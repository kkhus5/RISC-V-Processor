* File: AO211x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:02:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO211x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO211x2_ASAP7_75t_L.pex.sp.pex"
* File: AO211x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:02:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO211X2_ASAP7_75T_L%A1 2 5 8 11 13 23 25 26 32 VSS
c20 32 VSS 0.0154392f $X=0.0175 $Y=0.135
c21 26 VSS 6.352e-19 $X=0.0635 $Y=0.135
c22 25 VSS 9.99012e-19 $X=0.046 $Y=0.135
c23 23 VSS 5.74507e-19 $X=0.081 $Y=0.135
c24 11 VSS 0.00857795f $X=0.135 $Y=0.135
c25 8 VSS 0.0627962f $X=0.135 $Y=0.0675
c26 2 VSS 0.0686846f $X=0.081 $Y=0.135
r27 25 26 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r28 23 26 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r29 21 32 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r30 21 25 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.046 $Y2=0.135
r31 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r32 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r33 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r34 2 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r35 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
.ends

.subckt PM_AO211X2_ASAP7_75T_L%A2 2 7 10 13 21 29 VSS
c26 29 VSS 0.0040315f $X=0.137 $Y=0.1335
c27 21 VSS 7.18539e-19 $X=0.189 $Y=0.135
c28 10 VSS 0.0816994f $X=0.243 $Y=0.135
c29 2 VSS 0.0633997f $X=0.189 $Y=0.0675
r30 19 29 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.135 $Y2=0.135
r31 19 21 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.189 $Y2=0.135
r32 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r33 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r34 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r35 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r36 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO211X2_ASAP7_75T_L%B 2 7 10 13 25 VSS
c23 25 VSS 0.0114284f $X=0.298 $Y=0.1345
c24 10 VSS 0.0735411f $X=0.351 $Y=0.135
c25 2 VSS 0.0629692f $X=0.297 $Y=0.054
r26 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r27 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r28 5 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r29 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r30 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO211X2_ASAP7_75T_L%C 2 7 10 13 22 VSS
c13 22 VSS 0.00501966f $X=0.514 $Y=0.137
c14 10 VSS 0.0748382f $X=0.567 $Y=0.135
c15 2 VSS 0.0688401f $X=0.513 $Y=0.054
r16 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r17 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r18 5 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r19 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r20 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.054 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AO211X2_ASAP7_75T_L%7 2 7 10 13 15 17 22 25 27 30 32 33 36 37 39 40
+ 47 48 50 51 52 56 58 59 60 62 67 72 76 78 81 VSS
c56 85 VSS 7.08352e-19 $X=0.675 $Y=0.134
c57 81 VSS 0.00337493f $X=0.729 $Y=0.134
c58 78 VSS 0.0011573f $X=0.675 $Y=0.207
c59 77 VSS 0.00118958f $X=0.675 $Y=0.189
c60 76 VSS 0.00113947f $X=0.675 $Y=0.171
c61 75 VSS 7.78273e-19 $X=0.675 $Y=0.153
c62 74 VSS 0.00109324f $X=0.675 $Y=0.225
c63 72 VSS 0.00213713f $X=0.675 $Y=0.094
c64 71 VSS 0.00109324f $X=0.675 $Y=0.063
c65 70 VSS 0.00171628f $X=0.675 $Y=0.125
c66 68 VSS 0.00376564f $X=0.637 $Y=0.234
c67 67 VSS 0.00690843f $X=0.608 $Y=0.234
c68 62 VSS 0.00676815f $X=0.666 $Y=0.234
c69 61 VSS 0.00385934f $X=0.637 $Y=0.036
c70 60 VSS 0.00790562f $X=0.608 $Y=0.036
c71 59 VSS 0.00282595f $X=0.541 $Y=0.036
c72 58 VSS 0.00283359f $X=0.522 $Y=0.036
c73 56 VSS 0.0181937f $X=0.485 $Y=0.036
c74 52 VSS 5.50713e-19 $X=0.3175 $Y=0.036
c75 51 VSS 0.00739244f $X=0.311 $Y=0.036
c76 50 VSS 0.00537337f $X=0.252 $Y=0.036
c77 49 VSS 0.00245874f $X=0.215 $Y=0.036
c78 48 VSS 0.00487199f $X=0.203 $Y=0.036
c79 47 VSS 0.00290385f $X=0.144 $Y=0.036
c80 40 VSS 0.00544414f $X=0.108 $Y=0.036
c81 39 VSS 0.00198127f $X=0.108 $Y=0.036
c82 37 VSS 0.00625126f $X=0.666 $Y=0.036
c83 36 VSS 0.00358294f $X=0.54 $Y=0.2025
c84 32 VSS 6.74996e-19 $X=0.557 $Y=0.2025
c85 30 VSS 0.00534772f $X=0.488 $Y=0.054
c86 27 VSS 3.06948e-19 $X=0.503 $Y=0.054
c87 25 VSS 0.00581201f $X=0.322 $Y=0.054
c88 17 VSS 5.01261e-19 $X=0.125 $Y=0.0675
c89 13 VSS 0.00628305f $X=0.783 $Y=0.134
c90 10 VSS 0.0647467f $X=0.783 $Y=0.0675
c91 2 VSS 0.0652893f $X=0.729 $Y=0.0675
r92 79 85 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.134 $X2=0.675 $Y2=0.134
r93 79 81 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.134 $X2=0.729 $Y2=0.134
r94 77 78 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.189 $X2=0.675 $Y2=0.207
r95 76 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.171 $X2=0.675 $Y2=0.189
r96 75 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.153 $X2=0.675 $Y2=0.171
r97 74 78 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.225 $X2=0.675 $Y2=0.207
r98 73 85 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.143 $X2=0.675 $Y2=0.134
r99 73 75 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.143 $X2=0.675 $Y2=0.153
r100 71 72 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.063 $X2=0.675 $Y2=0.094
r101 70 85 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.125 $X2=0.675 $Y2=0.134
r102 70 72 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.125 $X2=0.675 $Y2=0.094
r103 69 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.045 $X2=0.675 $Y2=0.063
r104 67 68 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.608
+ $Y=0.234 $X2=0.637 $Y2=0.234
r105 64 67 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.608 $Y2=0.234
r106 62 74 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.234 $X2=0.675 $Y2=0.225
r107 62 68 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.234 $X2=0.637 $Y2=0.234
r108 60 61 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.608
+ $Y=0.036 $X2=0.637 $Y2=0.036
r109 59 60 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.541
+ $Y=0.036 $X2=0.608 $Y2=0.036
r110 58 59 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.541 $Y2=0.036
r111 56 57 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.485
+ $Y=0.036 $X2=0.4855 $Y2=0.036
r112 54 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.522 $Y2=0.036
r113 54 57 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.4855 $Y2=0.036
r114 51 52 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.036 $X2=0.3175 $Y2=0.036
r115 50 51 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.311 $Y2=0.036
r116 49 50 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.215
+ $Y=0.036 $X2=0.252 $Y2=0.036
r117 48 49 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.203
+ $Y=0.036 $X2=0.215 $Y2=0.036
r118 47 48 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.203 $Y2=0.036
r119 45 56 10.9321 $w=1.8e-08 $l=1.61e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.485 $Y2=0.036
r120 45 52 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.3175 $Y2=0.036
r121 39 47 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.144 $Y2=0.036
r122 39 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r123 37 69 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.036 $X2=0.675 $Y2=0.045
r124 37 61 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.637 $Y2=0.036
r125 36 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r126 33 36 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r127 32 36 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r128 30 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036
+ $X2=0.486 $Y2=0.036
r129 27 30 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.054 $X2=0.488 $Y2=0.054
r130 25 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r131 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.054 $X2=0.322 $Y2=0.054
r132 20 40 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.108 $Y=0.0675 $X2=0.108 $Y2=0.036
r133 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r134 13 15 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.134 $X2=0.783 $Y2=0.2025
r135 10 13 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.134
r136 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729 $Y=0.134
+ $X2=0.783 $Y2=0.134
r137 5 81 3.03549 $a=6.48e-16 $layer=V0LIG $count=2 $X=0.729 $Y=0.134 $X2=0.729
+ $Y2=0.134
r138 5 7 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.134 $X2=0.729 $Y2=0.2025
r139 2 5 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0675 $X2=0.729 $Y2=0.134
.ends

.subckt PM_AO211X2_ASAP7_75T_L%Y 1 2 6 7 10 14 16 23 28 29 30 VSS
c15 32 VSS 0.00270007f $X=0.837 $Y=0.184
c16 30 VSS 2.2091e-19 $X=0.837 $Y=0.13025
c17 29 VSS 0.00464972f $X=0.837 $Y=0.125
c18 28 VSS 5.1939e-19 $X=0.8375 $Y=0.1355
c19 26 VSS 0.00241318f $X=0.837 $Y=0.225
c20 24 VSS 0.00294383f $X=0.8125 $Y=0.234
c21 23 VSS 0.00532058f $X=0.797 $Y=0.234
c22 18 VSS 0.00579105f $X=0.828 $Y=0.234
c23 17 VSS 0.00294383f $X=0.8125 $Y=0.036
c24 16 VSS 0.00531887f $X=0.797 $Y=0.036
c25 14 VSS 0.00904224f $X=0.756 $Y=0.036
c26 11 VSS 0.00579105f $X=0.828 $Y=0.036
c27 10 VSS 0.00904121f $X=0.756 $Y=0.2025
c28 6 VSS 5.72268e-19 $X=0.773 $Y=0.2025
c29 1 VSS 5.72268e-19 $X=0.773 $Y=0.0675
r30 31 32 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.143 $X2=0.837 $Y2=0.184
r31 29 30 0.356481 $w=1.8e-08 $l=5.25e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.125 $X2=0.837 $Y2=0.13025
r32 28 31 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.1355 $X2=0.837 $Y2=0.143
r33 28 30 0.356481 $w=1.8e-08 $l=5.25e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.1355 $X2=0.837 $Y2=0.13025
r34 26 32 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.184
r35 25 29 5.4321 $w=1.8e-08 $l=8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.045 $X2=0.837 $Y2=0.125
r36 23 24 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.797
+ $Y=0.234 $X2=0.8125 $Y2=0.234
r37 20 23 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.797 $Y2=0.234
r38 18 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r39 18 24 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.8125 $Y2=0.234
r40 16 17 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.797
+ $Y=0.036 $X2=0.8125 $Y2=0.036
r41 13 16 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.797 $Y2=0.036
r42 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r43 11 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.036 $X2=0.837 $Y2=0.045
r44 11 17 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.8125 $Y2=0.036
r45 10 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234 $X2=0.756
+ $Y2=0.234
r46 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r47 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r48 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.756
+ $Y=0.0675 $X2=0.756 $Y2=0.036
r49 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
r50 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
.ends


* END of "./AO211x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO211x2_ASAP7_75t_L  VSS VDD A1 A2 B C Y
* 
* Y	Y
* C	C
* B	B
* A2	A2
* A1	A1
M0 noxref_11 N_A1_M0_g N_7_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M1 VSS N_A2_M1_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M2 N_7_M2_d N_B_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287 $Y=0.027
M3 VSS N_C_M3_g N_7_M3_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.503 $Y=0.027
M4 N_Y_M4_d N_7_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M5 N_Y_M5_d N_7_M5_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773 $Y=0.027
M6 VDD N_A1_M6_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 VDD N_A1_M7_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 VDD N_A2_M8_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 VDD N_A2_M9_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 noxref_9 N_B_M10_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 noxref_9 N_B_M11_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M12 N_7_M12_d N_C_M12_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M13 N_7_M13_d N_C_M13_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M14 N_Y_M14_d N_7_M14_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M15 N_Y_M15_d N_7_M15_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
*
* 
* .include "AO211x2_ASAP7_75t_L.pex.sp.AO211X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO211x2_ASAP7_75t_L.pex.sp.AO211X2_ASAP7_75T_L.pxi"
* File: AO211x2_ASAP7_75t_L.pex.sp.AO211X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:02:26 2017
* 
x_PM_AO211X2_ASAP7_75T_L%A1 N_A1_c_1_p N_A1_M6_g N_A1_M0_g N_A1_c_3_p N_A1_M7_g
+ N_A1_c_7_p N_A1_c_14_p N_A1_c_15_p A1 VSS PM_AO211X2_ASAP7_75T_L%A1
x_PM_AO211X2_ASAP7_75T_L%A2 N_A2_M1_g N_A2_M8_g N_A2_c_23_n N_A2_M9_g
+ N_A2_c_24_n A2 VSS PM_AO211X2_ASAP7_75T_L%A2
x_PM_AO211X2_ASAP7_75T_L%B N_B_M2_g N_B_M10_g N_B_c_49_n N_B_M11_g B VSS
+ PM_AO211X2_ASAP7_75T_L%B
x_PM_AO211X2_ASAP7_75T_L%C N_C_M3_g N_C_M12_g N_C_c_71_p N_C_M13_g C VSS
+ PM_AO211X2_ASAP7_75T_L%C
x_PM_AO211X2_ASAP7_75T_L%7 N_7_M4_g N_7_M14_g N_7_M5_g N_7_c_123_p N_7_M15_g
+ N_7_M0_s N_7_M2_d N_7_c_92_n N_7_M3_s N_7_c_98_n N_7_M13_d N_7_M12_d
+ N_7_c_100_n N_7_c_129_p N_7_c_83_n N_7_c_84_n N_7_c_86_n N_7_c_89_n N_7_c_93_n
+ N_7_c_94_n N_7_c_116_p N_7_c_97_n N_7_c_102_n N_7_c_104_n N_7_c_106_n
+ N_7_c_133_p N_7_c_107_n N_7_c_135_p N_7_c_115_p N_7_c_118_p N_7_c_130_p VSS
+ PM_AO211X2_ASAP7_75T_L%7
x_PM_AO211X2_ASAP7_75T_L%Y N_Y_M5_d N_Y_M4_d N_Y_M15_d N_Y_M14_d N_Y_c_141_n
+ N_Y_c_142_n N_Y_c_143_n N_Y_c_147_n Y N_Y_c_151_n N_Y_c_152_n VSS
+ PM_AO211X2_ASAP7_75T_L%Y
cc_1 N_A1_c_1_p N_A2_M1_g 2.69148e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_2 N_A1_M0_g N_A2_M1_g 0.00347357f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A1_c_3_p N_A2_c_23_n 0.0015471f $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_4 N_A1_c_3_p N_A2_c_24_n 5.75115e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_5 N_A1_M0_g A2 8.56946e-19 $X=0.135 $Y=0.0675 $X2=0.137 $Y2=0.1335
cc_6 N_A1_c_3_p A2 0.00274309f $X=0.135 $Y=0.135 $X2=0.137 $Y2=0.1335
cc_7 N_A1_c_7_p A2 9.16541e-19 $X=0.081 $Y=0.135 $X2=0.137 $Y2=0.1335
cc_8 A1 A2 0.00166694f $X=0.0175 $Y=0.135 $X2=0.137 $Y2=0.1335
cc_9 A1 N_7_c_83_n 8.45795e-19 $X=0.0175 $Y=0.135 $X2=0 $Y2=0
cc_10 N_A1_c_3_p N_7_c_84_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_11 A1 N_7_c_84_n 0.0011434f $X=0.0175 $Y=0.135 $X2=0 $Y2=0
cc_12 N_A1_M0_g N_7_c_86_n 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_13 VSS A1 0.00201602f $X=0.0175 $Y=0.135 $X2=0.189 $Y2=0.135
cc_14 VSS N_A1_c_14_p 2.97204e-19 $X=0.046 $Y=0.135 $X2=0.189 $Y2=0.135
cc_15 VSS N_A1_c_15_p 2.97204e-19 $X=0.0635 $Y=0.135 $X2=0.189 $Y2=0.135
cc_16 VSS A1 7.45437e-19 $X=0.0175 $Y=0.135 $X2=0.189 $Y2=0.135
cc_17 VSS N_A1_c_1_p 4.28653e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_18 VSS N_A1_c_3_p 3.24561e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_19 VSS N_A1_c_7_p 2.97204e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_20 VSS N_A1_M0_g 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_21 N_A2_M1_g N_B_M2_g 2.2125e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_22 N_A2_c_23_n N_B_M2_g 0.00333136f $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 N_A2_c_23_n N_B_c_49_n 0.00181947f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_24 N_A2_c_23_n B 0.00457636f $X=0.243 $Y=0.135 $X2=0.046 $Y2=0.135
cc_25 N_A2_c_24_n B 9.09825e-19 $X=0.189 $Y=0.135 $X2=0.046 $Y2=0.135
cc_26 A2 B 0.0018213f $X=0.137 $Y=0.1335 $X2=0.046 $Y2=0.135
cc_27 A2 N_7_c_84_n 0.00249808f $X=0.137 $Y=0.1335 $X2=0 $Y2=0
cc_28 A2 N_7_c_86_n 0.00374737f $X=0.137 $Y=0.1335 $X2=0 $Y2=0
cc_29 N_A2_M1_g N_7_c_89_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_A2_c_23_n N_7_c_89_n 3.09109e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 N_A2_c_24_n N_7_c_89_n 0.00121122f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_32 VSS A2 0.00156163f $X=0.137 $Y=0.1335 $X2=0.135 $Y2=0.135
cc_33 VSS A2 0.00375052f $X=0.137 $Y=0.1335 $X2=0.0175 $Y2=0.135
cc_34 VSS N_A2_c_24_n 0.00106008f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_35 VSS N_A2_M1_g 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_36 VSS N_A2_c_23_n 3.08494e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_37 VSS N_A2_c_23_n 2.34993e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_38 VSS N_A2_c_24_n 4.22525e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_39 N_B_c_49_n N_7_c_92_n 3.82299e-19 $X=0.351 $Y=0.135 $X2=0.046 $Y2=0.135
cc_40 B N_7_c_93_n 0.00350411f $X=0.298 $Y=0.1345 $X2=0 $Y2=0
cc_41 N_B_M2_g N_7_c_94_n 4.28653e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_42 N_B_c_49_n N_7_c_94_n 5.37757e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_43 B N_7_c_94_n 0.00103481f $X=0.298 $Y=0.1345 $X2=0 $Y2=0
cc_44 N_B_c_49_n N_7_c_97_n 4.62717e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_45 VSS B 0.00109884f $X=0.298 $Y=0.1345 $X2=0 $Y2=0
cc_46 VSS B 0.00375052f $X=0.298 $Y=0.1345 $X2=0 $Y2=0
cc_47 VSS B 5.23991e-19 $X=0.298 $Y=0.1345 $X2=0 $Y2=0
cc_48 VSS N_B_c_49_n 2.21754e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_49 VSS N_B_M2_g 4.28653e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_50 VSS B 5.23991e-19 $X=0.298 $Y=0.1345 $X2=0 $Y2=0
cc_51 VSS N_B_c_49_n 3.8028e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_52 VSS N_B_c_49_n 9.18375e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_53 VSS N_B_c_49_n 7.96506e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_54 VSS B 3.71763e-19 $X=0.298 $Y=0.1345 $X2=0 $Y2=0
cc_55 VSS N_B_c_49_n 3.97719e-19 $X=0.351 $Y=0.135 $X2=0.046 $Y2=0.135
cc_56 C N_7_c_98_n 0.00237967f $X=0.514 $Y=0.137 $X2=0 $Y2=0
cc_57 N_C_c_71_p N_7_M13_d 3.78279e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_58 N_C_c_71_p N_7_c_100_n 9.18375e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_59 C N_7_c_100_n 9.22768e-19 $X=0.514 $Y=0.137 $X2=0 $Y2=0
cc_60 N_C_M3_g N_7_c_102_n 2.34993e-19 $X=0.513 $Y=0.054 $X2=0 $Y2=0
cc_61 C N_7_c_102_n 0.00372137f $X=0.514 $Y=0.137 $X2=0 $Y2=0
cc_62 N_C_c_71_p N_7_c_104_n 7.31733e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_63 C N_7_c_104_n 2.5188e-19 $X=0.514 $Y=0.137 $X2=0 $Y2=0
cc_64 N_C_c_71_p N_7_c_106_n 4.62717e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_65 N_C_c_71_p N_7_c_107_n 2.64781e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_66 VSS N_C_M3_g 3.4229e-19 $X=0.513 $Y=0.054 $X2=0 $Y2=0
cc_67 VSS C 0.00373221f $X=0.514 $Y=0.137 $X2=0 $Y2=0
cc_68 VSS N_C_c_71_p 8.30831e-19 $X=0.567 $Y=0.135 $X2=0.297 $Y2=0.135
cc_69 VSS N_7_c_107_n 2.83135e-19 $X=0.608 $Y=0.234 $X2=0 $Y2=0
cc_70 VSS N_7_c_92_n 9.98826e-19 $X=0.322 $Y=0.054 $X2=0.081 $Y2=0.2025
cc_71 VSS N_7_c_98_n 8.59825e-19 $X=0.488 $Y=0.054 $X2=0 $Y2=0
cc_72 VSS N_7_c_100_n 0.00338163f $X=0.54 $Y=0.2025 $X2=0 $Y2=0
cc_73 VSS N_7_c_107_n 5.08059e-19 $X=0.608 $Y=0.234 $X2=0 $Y2=0
cc_74 VSS N_7_c_100_n 0.00369676f $X=0.54 $Y=0.2025 $X2=0 $Y2=0
cc_75 VSS N_7_c_107_n 0.00313156f $X=0.608 $Y=0.234 $X2=0 $Y2=0
cc_76 VSS N_7_c_115_p 4.23807e-19 $X=0.675 $Y=0.171 $X2=0 $Y2=0
cc_77 VSS N_7_c_116_p 7.89965e-19 $X=0.3175 $Y=0.036 $X2=0 $Y2=0
cc_78 VSS N_7_c_97_n 7.89965e-19 $X=0.485 $Y=0.036 $X2=0.046 $Y2=0.135
cc_79 VSS N_7_c_118_p 6.12996e-19 $X=0.675 $Y=0.207 $X2=0 $Y2=0
cc_80 VSS N_7_c_100_n 0.00126629f $X=0.54 $Y=0.2025 $X2=0.0175 $Y2=0.135
cc_81 VSS N_7_c_107_n 0.00678111f $X=0.608 $Y=0.234 $X2=0.0175 $Y2=0.135
cc_82 VSS N_7_c_100_n 0.00112576f $X=0.54 $Y=0.2025 $X2=0 $Y2=0
cc_83 VSS N_7_c_106_n 7.89965e-19 $X=0.608 $Y=0.036 $X2=0 $Y2=0
cc_84 N_7_c_123_p N_Y_M5_d 3.73743e-19 $X=0.783 $Y=0.134 $X2=0.081 $Y2=0.135
cc_85 N_7_c_123_p N_Y_M15_d 3.61125e-19 $X=0.783 $Y=0.134 $X2=0 $Y2=0
cc_86 N_7_c_123_p N_Y_c_141_n 4.78826e-19 $X=0.783 $Y=0.134 $X2=0.135 $Y2=0.135
cc_87 N_7_c_123_p N_Y_c_142_n 5.26265e-19 $X=0.783 $Y=0.134 $X2=0 $Y2=0
cc_88 N_7_M5_g N_Y_c_143_n 4.11429e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_89 N_7_c_123_p N_Y_c_143_n 4.0761e-19 $X=0.783 $Y=0.134 $X2=0 $Y2=0
cc_90 N_7_c_129_p N_Y_c_143_n 4.02904e-19 $X=0.666 $Y=0.036 $X2=0 $Y2=0
cc_91 N_7_c_130_p N_Y_c_143_n 7.6376e-19 $X=0.729 $Y=0.134 $X2=0 $Y2=0
cc_92 N_7_M5_g N_Y_c_147_n 4.32902e-19 $X=0.783 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_93 N_7_c_123_p N_Y_c_147_n 4.02718e-19 $X=0.783 $Y=0.134 $X2=0.081 $Y2=0.135
cc_94 N_7_c_133_p N_Y_c_147_n 3.9751e-19 $X=0.666 $Y=0.234 $X2=0.081 $Y2=0.135
cc_95 N_7_c_130_p N_Y_c_147_n 7.42958e-19 $X=0.729 $Y=0.134 $X2=0.081 $Y2=0.135
cc_96 N_7_c_135_p N_Y_c_151_n 3.20931e-19 $X=0.675 $Y=0.094 $X2=0 $Y2=0
cc_97 N_7_c_123_p N_Y_c_152_n 5.24018e-19 $X=0.783 $Y=0.134 $X2=0 $Y2=0
cc_98 N_7_c_130_p N_Y_c_152_n 0.00101708f $X=0.729 $Y=0.134 $X2=0 $Y2=0
cc_99 VSS N_7_c_89_n 4.14303e-19 $X=0.203 $Y=0.036 $X2=0.081 $Y2=0.135

* END of "./AO211x2_ASAP7_75t_L.pex.sp.AO211X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO21x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:02:49 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO21x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO21x1_ASAP7_75t_L.pex.sp.pex"
* File: AO21x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:02:49 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO21X1_ASAP7_75T_L%A1 2 5 7 17 VSS
c9 17 VSS 0.0149008f $X=0.0795 $Y=0.1355
c10 5 VSS 0.00273001f $X=0.081 $Y=0.135
c11 2 VSS 0.0661158f $X=0.081 $Y=0.0675
r12 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO21X1_ASAP7_75T_L%A2 2 5 7 10 VSS
c11 10 VSS 0.00170642f $X=0.1315 $Y=0.1355
c12 5 VSS 0.00129484f $X=0.135 $Y=0.135
c13 2 VSS 0.0614068f $X=0.135 $Y=0.0675
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO21X1_ASAP7_75T_L%B 2 5 7 10 VSS
c12 10 VSS 0.0016481f $X=0.1865 $Y=0.1355
c13 5 VSS 0.00110432f $X=0.189 $Y=0.135
c14 2 VSS 0.0607131f $X=0.189 $Y=0.0675
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO21X1_ASAP7_75T_L%6 2 5 7 9 10 14 15 18 21 27 29 31 33 34 37 40 44
+ VSS
c27 49 VSS 3.38114e-19 $X=0.243 $Y=0.1765
c28 47 VSS 3.56487e-19 $X=0.243 $Y=0.07
c29 46 VSS 2.62061e-20 $X=0.243 $Y=0.063
c30 44 VSS 0.0013899f $X=0.243 $Y=0.135
c31 40 VSS 0.00146362f $X=0.198 $Y=0.036
c32 39 VSS 0.00409617f $X=0.18 $Y=0.036
c33 37 VSS 0.00780544f $X=0.162 $Y=0.036
c34 34 VSS 0.00785727f $X=0.234 $Y=0.036
c35 33 VSS 4.97894e-20 $X=0.232 $Y=0.198
c36 32 VSS 0.00354056f $X=0.23 $Y=0.198
c37 31 VSS 5.31938e-19 $X=0.198 $Y=0.198
c38 30 VSS 2.03419e-19 $X=0.18 $Y=0.198
c39 29 VSS 2.44387e-19 $X=0.176 $Y=0.198
c40 28 VSS 1.23838e-19 $X=0.148 $Y=0.198
c41 27 VSS 8.46035e-21 $X=0.144 $Y=0.198
c42 26 VSS 5.69672e-19 $X=0.126 $Y=0.198
c43 21 VSS 1.3844e-19 $X=0.108 $Y=0.198
c44 19 VSS 8.26569e-20 $X=0.234 $Y=0.198
c45 18 VSS 0.00243919f $X=0.108 $Y=0.2025
c46 14 VSS 6.06806e-19 $X=0.125 $Y=0.2025
c47 9 VSS 5.72268e-19 $X=0.179 $Y=0.0675
c48 5 VSS 0.00173625f $X=0.243 $Y=0.135
c49 2 VSS 0.0654755f $X=0.243 $Y=0.0675
r50 48 49 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.164 $X2=0.243 $Y2=0.1765
r51 46 47 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.063 $X2=0.243 $Y2=0.07
r52 44 48 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.164
r53 44 47 4.41358 $w=1.8e-08 $l=6.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.07
r54 42 49 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.1765
r55 41 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.063
r56 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r57 36 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r58 36 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r59 34 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r60 34 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.198 $Y2=0.036
r61 32 33 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.198 $X2=0.232 $Y2=0.198
r62 31 32 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.198 $X2=0.23 $Y2=0.198
r63 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.198 $X2=0.198 $Y2=0.198
r64 29 30 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.198 $X2=0.18 $Y2=0.198
r65 28 29 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.198 $X2=0.176 $Y2=0.198
r66 27 28 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.198 $X2=0.148 $Y2=0.198
r67 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.198 $X2=0.144 $Y2=0.198
r68 21 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.198 $X2=0.126 $Y2=0.198
r69 19 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.198 $X2=0.243 $Y2=0.189
r70 19 33 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.232 $Y2=0.198
r71 18 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.198 $X2=0.108
+ $Y2=0.198
r72 15 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r73 14 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r74 13 37 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r75 10 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r76 9 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r77 5 44 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r78 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r79 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO21X1_ASAP7_75T_L%Y 1 4 6 9 17 21 23 VSS
c8 23 VSS 0.00999953f $X=0.286 $Y=0.202
c9 17 VSS 0.00839825f $X=0.286 $Y=0.054
c10 9 VSS 0.0126254f $X=0.268 $Y=0.2025
c11 4 VSS 0.0168216f $X=0.268 $Y=0.0675
r12 21 23 5.94136 $w=1.8e-08 $l=8.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.286
+ $Y=0.1145 $X2=0.286 $Y2=0.202
r13 17 21 4.10802 $w=1.8e-08 $l=6.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.286
+ $Y=0.054 $X2=0.286 $Y2=0.1145
r14 9 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.286 $Y=0.202 $X2=0.286
+ $Y2=0.202
r15 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.2025 $X2=0.268 $Y2=0.2025
r16 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.286 $Y=0.054 $X2=0.286
+ $Y2=0.054
r17 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.268 $Y2=0.0675
.ends


* END of "./AO21x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO21x1_ASAP7_75t_L  VSS VDD A1 A2 B Y
* 
* Y	Y
* B	B
* A2	A2
* A1	A1
M0 noxref_9 N_A1_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_A2_M1_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_B_M2_g N_6_M2_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_6_M3_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_6_M4_d N_A1_M4_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 noxref_7 N_A2_M5_g N_6_M5_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 VDD N_B_M6_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M7 N_Y_M7_d N_6_M7_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
*
* 
* .include "AO21x1_ASAP7_75t_L.pex.sp.AO21X1_ASAP7_75T_L.pxi"
* BEGIN of "./AO21x1_ASAP7_75t_L.pex.sp.AO21X1_ASAP7_75T_L.pxi"
* File: AO21x1_ASAP7_75t_L.pex.sp.AO21X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:02:49 2017
* 
x_PM_AO21X1_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M4_g A1 VSS
+ PM_AO21X1_ASAP7_75T_L%A1
x_PM_AO21X1_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_11_n N_A2_M5_g A2 VSS
+ PM_AO21X1_ASAP7_75T_L%A2
x_PM_AO21X1_ASAP7_75T_L%B N_B_M2_g N_B_c_23_n N_B_M6_g B VSS
+ PM_AO21X1_ASAP7_75T_L%B
x_PM_AO21X1_ASAP7_75T_L%6 N_6_M3_g N_6_c_39_n N_6_M7_g N_6_M2_s N_6_M1_d
+ N_6_M5_s N_6_M4_d N_6_c_46_p N_6_c_33_n N_6_c_35_n N_6_c_49_p N_6_c_40_n
+ N_6_c_59_p N_6_c_54_p N_6_c_37_n N_6_c_43_n N_6_c_45_n VSS
+ PM_AO21X1_ASAP7_75T_L%6
x_PM_AO21X1_ASAP7_75T_L%Y N_Y_M3_d N_Y_c_60_n N_Y_M7_d N_Y_c_62_n N_Y_c_63_n Y
+ N_Y_c_64_n VSS PM_AO21X1_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00361888f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_11_n 0.00120928f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A1 A2 0.00207308f $X=0.0795 $Y=0.1355 $X2=0.1315 $Y2=0.1355
cc_4 N_A1_M0_g N_B_M2_g 2.98169e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 A1 N_6_c_33_n 5.28865e-19 $X=0.0795 $Y=0.1355 $X2=0 $Y2=0
cc_6 VSS A1 0.00230205f $X=0.0795 $Y=0.1355 $X2=0.135 $Y2=0.135
cc_7 VSS A1 0.00134496f $X=0.0795 $Y=0.1355 $X2=0.135 $Y2=0.135
cc_8 VSS N_A1_M0_g 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_9 VSS A1 2.99763e-19 $X=0.0795 $Y=0.1355 $X2=0 $Y2=0
cc_10 N_A2_M1_g N_B_M2_g 0.00354623f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_11 N_A2_c_11_n N_B_c_23_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_12 A2 B 0.00406615f $X=0.1315 $Y=0.1355 $X2=0 $Y2=0
cc_13 N_A2_M1_g N_6_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_A2_M1_g N_6_c_35_n 2.76185e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 A2 N_6_c_35_n 0.0012322f $X=0.1315 $Y=0.1355 $X2=0 $Y2=0
cc_16 A2 N_6_c_37_n 0.0013399f $X=0.1315 $Y=0.1355 $X2=0 $Y2=0
cc_17 VSS N_A2_M1_g 2.08515e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_18 N_B_M2_g N_6_M3_g 0.00287079f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_19 N_B_c_23_n N_6_c_39_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_20 N_B_M2_g N_6_c_40_n 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_21 B N_6_c_40_n 0.0012322f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_22 B N_6_c_37_n 0.00114532f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_23 N_B_M2_g N_6_c_43_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 B N_6_c_43_n 0.00124805f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_25 B N_6_c_45_n 0.0037803f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_26 VSS N_6_c_46_p 0.00353012f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_27 VSS N_6_c_33_n 3.60466e-19 $X=0.108 $Y=0.198 $X2=0.081 $Y2=0.135
cc_28 VSS N_6_c_46_p 0.0035219f $X=0.108 $Y=0.2025 $X2=0 $Y2=0
cc_29 VSS N_6_c_49_p 0.00233206f $X=0.176 $Y=0.198 $X2=0 $Y2=0
cc_30 VSS N_6_c_37_n 0.00138157f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_31 VSS N_6_c_35_n 0.00347702f $X=0.144 $Y=0.198 $X2=0 $Y2=0
cc_32 VSS N_6_c_46_p 0.00248803f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_33 VSS N_6_c_33_n 0.00347702f $X=0.108 $Y=0.198 $X2=0.081 $Y2=0.135
cc_34 N_6_c_54_p N_Y_c_60_n 0.00182327f $X=0.234 $Y=0.036 $X2=0.081 $Y2=0.135
cc_35 N_6_c_37_n N_Y_c_60_n 3.37765e-19 $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_36 N_6_c_45_n N_Y_c_62_n 0.00104853f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_37 N_6_c_54_p N_Y_c_63_n 0.00957806f $X=0.234 $Y=0.036 $X2=0.0795 $Y2=0.1355
cc_38 N_6_M3_g N_Y_c_64_n 2.34993e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_6_c_59_p N_Y_c_64_n 0.00232476f $X=0.232 $Y=0.198 $X2=0 $Y2=0
cc_40 VSS N_Y_c_62_n 2.41798e-19 $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_41 VSS N_Y_c_64_n 4.32936e-19 $X=0.162 $Y=0.234 $X2=0 $Y2=0

* END of "./AO21x1_ASAP7_75t_L.pex.sp.AO21X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO21x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:03:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO21x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO21x2_ASAP7_75t_L.pex.sp.pex"
* File: AO21x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:03:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO21X2_ASAP7_75T_L%A1 2 5 7 17 VSS
c9 17 VSS 0.0149008f $X=0.0795 $Y=0.1355
c10 5 VSS 0.00273001f $X=0.081 $Y=0.135
c11 2 VSS 0.0661158f $X=0.081 $Y=0.0675
r12 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO21X2_ASAP7_75T_L%A2 2 5 7 10 VSS
c11 10 VSS 0.00170642f $X=0.1315 $Y=0.1355
c12 5 VSS 0.00129794f $X=0.135 $Y=0.135
c13 2 VSS 0.0614068f $X=0.135 $Y=0.0675
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO21X2_ASAP7_75T_L%B 2 5 7 10 VSS
c13 10 VSS 0.00173245f $X=0.1865 $Y=0.1355
c14 5 VSS 9.84213e-19 $X=0.189 $Y=0.135
c15 2 VSS 0.0593522f $X=0.189 $Y=0.0675
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO21X2_ASAP7_75T_L%6 2 7 10 13 15 17 18 22 23 26 29 35 37 39 41 42 45
+ 48 52 56 57 VSS
c37 59 VSS 3.38114e-19 $X=0.243 $Y=0.1765
c38 57 VSS 6.71733e-19 $X=0.243 $Y=0.111
c39 56 VSS 5.07501e-19 $X=0.243 $Y=0.087
c40 55 VSS 3.56487e-19 $X=0.243 $Y=0.07
c41 54 VSS 2.8341e-20 $X=0.243 $Y=0.063
c42 52 VSS 2.57607e-19 $X=0.243 $Y=0.135
c43 48 VSS 0.00146362f $X=0.198 $Y=0.036
c44 47 VSS 0.00409617f $X=0.18 $Y=0.036
c45 45 VSS 0.00780542f $X=0.162 $Y=0.036
c46 42 VSS 0.00785727f $X=0.234 $Y=0.036
c47 41 VSS 4.97894e-20 $X=0.232 $Y=0.198
c48 40 VSS 0.00354056f $X=0.23 $Y=0.198
c49 39 VSS 5.31938e-19 $X=0.198 $Y=0.198
c50 38 VSS 2.03419e-19 $X=0.18 $Y=0.198
c51 37 VSS 2.44387e-19 $X=0.176 $Y=0.198
c52 36 VSS 1.23838e-19 $X=0.148 $Y=0.198
c53 35 VSS 8.46035e-21 $X=0.144 $Y=0.198
c54 34 VSS 5.69672e-19 $X=0.126 $Y=0.198
c55 29 VSS 1.3844e-19 $X=0.108 $Y=0.198
c56 27 VSS 5.71502e-20 $X=0.234 $Y=0.198
c57 26 VSS 0.00243919f $X=0.108 $Y=0.2025
c58 22 VSS 6.06806e-19 $X=0.125 $Y=0.2025
c59 17 VSS 5.72268e-19 $X=0.179 $Y=0.0675
c60 13 VSS 0.00430272f $X=0.297 $Y=0.135
c61 10 VSS 0.0648587f $X=0.297 $Y=0.0675
c62 2 VSS 0.0608946f $X=0.243 $Y=0.0675
r63 58 59 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.164 $X2=0.243 $Y2=0.1765
r64 56 57 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.087 $X2=0.243 $Y2=0.111
r65 55 56 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.07 $X2=0.243 $Y2=0.087
r66 54 55 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.063 $X2=0.243 $Y2=0.07
r67 52 58 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.164
r68 52 57 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.111
r69 50 59 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.1765
r70 49 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.063
r71 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r72 44 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r73 44 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r74 42 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r75 42 48 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.198 $Y2=0.036
r76 40 41 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.198 $X2=0.232 $Y2=0.198
r77 39 40 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.198 $X2=0.23 $Y2=0.198
r78 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.198 $X2=0.198 $Y2=0.198
r79 37 38 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.198 $X2=0.18 $Y2=0.198
r80 36 37 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.198 $X2=0.176 $Y2=0.198
r81 35 36 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.198 $X2=0.148 $Y2=0.198
r82 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.198 $X2=0.144 $Y2=0.198
r83 29 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.198 $X2=0.126 $Y2=0.198
r84 27 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.198 $X2=0.243 $Y2=0.189
r85 27 41 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.232 $Y2=0.198
r86 26 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.198 $X2=0.108
+ $Y2=0.198
r87 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r88 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r89 21 45 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r90 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r91 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r92 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r93 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r94 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r95 5 52 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r96 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r97 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO21X2_ASAP7_75T_L%Y 1 2 5 6 7 10 11 13 20 25 29 VSS
c16 29 VSS 0.00271292f $X=0.285 $Y=0.054
c17 27 VSS 8.50351e-19 $X=0.324 $Y=0.216
c18 25 VSS 0.00909353f $X=0.3225 $Y=0.1145
c19 23 VSS 8.0311e-19 $X=0.324 $Y=0.225
c20 20 VSS 0.00365977f $X=0.315 $Y=0.078
c21 19 VSS 0.00189536f $X=0.2955 $Y=0.234
c22 18 VSS 0.00132025f $X=0.276 $Y=0.234
c23 13 VSS 0.00392797f $X=0.27 $Y=0.234
c24 11 VSS 0.00618369f $X=0.315 $Y=0.234
c25 10 VSS 0.010528f $X=0.27 $Y=0.2025
c26 6 VSS 5.38922e-19 $X=0.287 $Y=0.2025
c27 5 VSS 0.014693f $X=0.27 $Y=0.0675
c28 1 VSS 5.1537e-19 $X=0.287 $Y=0.0675
r29 29 32 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.285
+ $Y=0.054 $X2=0.285 $Y2=0.078
r30 26 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.207 $X2=0.324 $Y2=0.216
r31 25 26 6.28086 $w=1.8e-08 $l=9.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.1145 $X2=0.324 $Y2=0.207
r32 23 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.225 $X2=0.324 $Y2=0.216
r33 22 25 1.86728 $w=1.8e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.087 $X2=0.324 $Y2=0.1145
r34 21 32 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.294
+ $Y=0.078 $X2=0.285 $Y2=0.078
r35 20 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.315 $Y=0.078 $X2=0.324 $Y2=0.087
r36 20 21 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.315
+ $Y=0.078 $X2=0.294 $Y2=0.078
r37 18 19 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.276
+ $Y=0.234 $X2=0.2955 $Y2=0.234
r38 13 18 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.276 $Y2=0.234
r39 11 23 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.315 $Y=0.234 $X2=0.324 $Y2=0.225
r40 11 19 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.315
+ $Y=0.234 $X2=0.2955 $Y2=0.234
r41 10 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r42 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r43 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r44 5 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.285 $Y=0.054 $X2=0.285
+ $Y2=0.054
r45 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
r46 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends


* END of "./AO21x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO21x2_ASAP7_75t_L  VSS VDD A1 A2 B Y
* 
* Y	Y
* B	B
* A2	A2
* A1	A1
M0 noxref_9 N_A1_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_A2_M1_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_B_M2_g N_6_M2_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_6_M3_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_6_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_6_M5_d N_A1_M5_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M6 noxref_7 N_A2_M6_g N_6_M6_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 VDD N_B_M7_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M8 N_Y_M8_d N_6_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M9 N_Y_M9_d N_6_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
*
* 
* .include "AO21x2_ASAP7_75t_L.pex.sp.AO21X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO21x2_ASAP7_75t_L.pex.sp.AO21X2_ASAP7_75T_L.pxi"
* File: AO21x2_ASAP7_75t_L.pex.sp.AO21X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:03:11 2017
* 
x_PM_AO21X2_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M5_g A1 VSS
+ PM_AO21X2_ASAP7_75T_L%A1
x_PM_AO21X2_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_11_n N_A2_M6_g A2 VSS
+ PM_AO21X2_ASAP7_75T_L%A2
x_PM_AO21X2_ASAP7_75T_L%B N_B_M2_g N_B_c_23_n N_B_M7_g B VSS
+ PM_AO21X2_ASAP7_75T_L%B
x_PM_AO21X2_ASAP7_75T_L%6 N_6_M3_g N_6_M8_g N_6_M4_g N_6_c_41_n N_6_M9_g
+ N_6_M2_s N_6_M1_d N_6_M6_s N_6_M5_d N_6_c_48_p N_6_c_34_n N_6_c_36_n
+ N_6_c_51_p N_6_c_42_n N_6_c_66_p N_6_c_58_p N_6_c_38_n N_6_c_45_n N_6_c_62_p
+ N_6_c_47_n N_6_c_68_p VSS PM_AO21X2_ASAP7_75T_L%6
x_PM_AO21X2_ASAP7_75T_L%Y N_Y_M4_d N_Y_M3_d N_Y_c_71_n N_Y_M9_d N_Y_M8_d
+ N_Y_c_76_n N_Y_c_78_n N_Y_c_79_n N_Y_c_82_n Y N_Y_c_84_n VSS
+ PM_AO21X2_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00361888f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_11_n 0.00120928f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A1 A2 0.00207308f $X=0.0795 $Y=0.1355 $X2=0.1315 $Y2=0.1355
cc_4 N_A1_M0_g N_B_M2_g 2.98169e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 A1 N_6_c_34_n 5.28865e-19 $X=0.0795 $Y=0.1355 $X2=0 $Y2=0
cc_6 VSS A1 0.00230205f $X=0.0795 $Y=0.1355 $X2=0.135 $Y2=0.135
cc_7 VSS A1 0.00134496f $X=0.0795 $Y=0.1355 $X2=0.135 $Y2=0.135
cc_8 VSS N_A1_M0_g 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_9 VSS A1 2.99763e-19 $X=0.0795 $Y=0.1355 $X2=0 $Y2=0
cc_10 N_A2_M1_g N_B_M2_g 0.00354623f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_11 N_A2_c_11_n N_B_c_23_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_12 A2 B 0.00406615f $X=0.1315 $Y=0.1355 $X2=0 $Y2=0
cc_13 N_A2_M1_g N_6_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_A2_M1_g N_6_c_36_n 2.76185e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 A2 N_6_c_36_n 0.0012322f $X=0.1315 $Y=0.1355 $X2=0 $Y2=0
cc_16 A2 N_6_c_38_n 0.0013399f $X=0.1315 $Y=0.1355 $X2=0 $Y2=0
cc_17 VSS N_A2_M1_g 2.08515e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_18 N_B_M2_g N_6_M3_g 0.00287079f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_19 N_B_M2_g N_6_M4_g 2.34385e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_20 N_B_c_23_n N_6_c_41_n 9.59209e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_21 N_B_M2_g N_6_c_42_n 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_22 B N_6_c_42_n 0.0012322f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_23 B N_6_c_38_n 0.00114532f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_24 N_B_M2_g N_6_c_45_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_25 B N_6_c_45_n 0.00124805f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_26 B N_6_c_47_n 0.00377326f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_27 VSS N_6_c_48_p 0.00353012f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_28 VSS N_6_c_34_n 3.60466e-19 $X=0.108 $Y=0.198 $X2=0.081 $Y2=0.135
cc_29 VSS N_6_c_48_p 0.0035219f $X=0.108 $Y=0.2025 $X2=0 $Y2=0
cc_30 VSS N_6_c_51_p 0.00233206f $X=0.176 $Y=0.198 $X2=0 $Y2=0
cc_31 VSS N_6_c_38_n 0.00138157f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_32 VSS N_6_c_36_n 0.00347702f $X=0.144 $Y=0.198 $X2=0 $Y2=0
cc_33 VSS N_6_c_48_p 0.00248803f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_34 VSS N_6_c_34_n 0.00347702f $X=0.108 $Y=0.198 $X2=0.081 $Y2=0.135
cc_35 N_6_M4_g N_Y_c_71_n 0.00293521f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_36 N_6_c_41_n N_Y_c_71_n 0.00187466f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_37 N_6_c_58_p N_Y_c_71_n 0.00176852f $X=0.234 $Y=0.036 $X2=0.081 $Y2=0.135
cc_38 N_6_c_38_n N_Y_c_71_n 3.05411e-19 $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_39 N_6_c_41_n N_Y_M9_d 3.80663e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_40 N_6_c_41_n N_Y_c_76_n 8.00061e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_41 N_6_c_62_p N_Y_c_76_n 0.0015568f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_42 N_6_M4_g N_Y_c_78_n 2.57944e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_6_M3_g N_Y_c_79_n 2.34993e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_6_c_41_n N_Y_c_79_n 6.95747e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_45 N_6_c_66_p N_Y_c_79_n 0.00232476f $X=0.232 $Y=0.198 $X2=0 $Y2=0
cc_46 N_6_M4_g N_Y_c_82_n 3.12785e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_47 N_6_c_68_p Y 0.00214255f $X=0.243 $Y=0.111 $X2=0 $Y2=0
cc_48 N_6_c_41_n N_Y_c_84_n 5.04561e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_49 N_6_c_58_p N_Y_c_84_n 0.00318733f $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_50 VSS N_Y_c_79_n 4.45935e-19 $X=0.162 $Y=0.234 $X2=0 $Y2=0

* END of "./AO21x2_ASAP7_75t_L.pex.sp.AO21X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO221x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:03:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO221x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO221x1_ASAP7_75t_L.pex.sp.pex"
* File: AO221x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:03:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO221X1_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c11 10 VSS 6.95749e-19 $X=0.081 $Y=0.135
c12 5 VSS 0.00170784f $X=0.081 $Y=0.135
c13 2 VSS 0.0655264f $X=0.081 $Y=0.054
r14 10 14 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.148
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO221X1_ASAP7_75T_L%B2 2 5 7 10 VSS
c11 10 VSS 0.00105185f $X=0.133 $Y=0.109
c12 5 VSS 0.00114017f $X=0.135 $Y=0.135
c13 2 VSS 0.0608869f $X=0.135 $Y=0.054
r14 10 13 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.109 $X2=0.135 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO221X1_ASAP7_75T_L%C 2 5 7 10 VSS
c11 10 VSS 0.00138457f $X=0.188 $Y=0.123
c12 5 VSS 0.00120688f $X=0.189 $Y=0.135
c13 2 VSS 0.0599046f $X=0.189 $Y=0.054
r14 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.123 $X2=0.189 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO221X1_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c12 10 VSS 6.84433e-19 $X=0.243 $Y=0.135
c13 5 VSS 0.00114323f $X=0.243 $Y=0.135
c14 2 VSS 0.0596104f $X=0.243 $Y=0.054
r15 10 14 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.151
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO221X1_ASAP7_75T_L%A2 2 5 7 10 13 VSS
c9 13 VSS 5.28209e-19 $X=0.297 $Y=0.135
c10 10 VSS 7.94635e-19 $X=0.295 $Y=0.123
c11 5 VSS 0.00212633f $X=0.297 $Y=0.135
c12 2 VSS 0.0616967f $X=0.297 $Y=0.054
r13 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.123 $X2=0.297 $Y2=0.135
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO221X1_ASAP7_75T_L%8 2 5 7 9 12 14 15 18 19 20 23 27 28 37 39 42 44
+ 45 46 47 48 52 55 56 61 62 65 VSS
c37 65 VSS 0.00332792f $X=0.459 $Y=0.135
c38 63 VSS 0.00126105f $X=0.414 $Y=0.135
c39 62 VSS 0.00140379f $X=0.405 $Y=0.098
c40 61 VSS 0.00198282f $X=0.405 $Y=0.07
c41 60 VSS 9.72353e-19 $X=0.405 $Y=0.126
c42 57 VSS 1.45514e-19 $X=0.099 $Y=0.198
c43 56 VSS 8.46035e-21 $X=0.09 $Y=0.198
c44 55 VSS 4.76765e-19 $X=0.072 $Y=0.198
c45 54 VSS 1.91267e-19 $X=0.039 $Y=0.198
c46 52 VSS 5.70579e-19 $X=0.108 $Y=0.198
c47 50 VSS 0.00193008f $X=0.036 $Y=0.198
c48 49 VSS 0.00395192f $X=0.3675 $Y=0.036
c49 48 VSS 0.00611566f $X=0.339 $Y=0.036
c50 47 VSS 0.00146362f $X=0.306 $Y=0.036
c51 46 VSS 0.00368202f $X=0.288 $Y=0.036
c52 45 VSS 0.00146362f $X=0.252 $Y=0.036
c53 44 VSS 0.00331014f $X=0.234 $Y=0.036
c54 43 VSS 1.99947e-19 $X=0.2 $Y=0.036
c55 42 VSS 0.00142296f $X=0.198 $Y=0.036
c56 41 VSS 4.31197e-19 $X=0.18 $Y=0.036
c57 40 VSS 0.00564793f $X=0.176 $Y=0.036
c58 39 VSS 0.00146362f $X=0.144 $Y=0.036
c59 38 VSS 0.00345019f $X=0.126 $Y=0.036
c60 37 VSS 0.00146362f $X=0.09 $Y=0.036
c61 36 VSS 0.00353842f $X=0.072 $Y=0.036
c62 29 VSS 0.00340187f $X=0.036 $Y=0.036
c63 28 VSS 0.00653563f $X=0.396 $Y=0.036
c64 27 VSS 0.00423691f $X=0.027 $Y=0.164
c65 26 VSS 9.59589e-19 $X=0.027 $Y=0.07
c66 25 VSS 0.00112176f $X=0.027 $Y=0.189
c67 23 VSS 0.00233317f $X=0.108 $Y=0.2025
c68 19 VSS 5.91014e-19 $X=0.125 $Y=0.2025
c69 18 VSS 0.00607665f $X=0.216 $Y=0.054
c70 14 VSS 5.19811e-19 $X=0.233 $Y=0.054
c71 12 VSS 0.00319205f $X=0.056 $Y=0.054
c72 9 VSS 2.6657e-19 $X=0.071 $Y=0.054
c73 5 VSS 0.00384591f $X=0.459 $Y=0.135
c74 2 VSS 0.06855f $X=0.459 $Y=0.0675
r75 63 65 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.135 $X2=0.459 $Y2=0.135
r76 61 62 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.07 $X2=0.405 $Y2=0.098
r77 60 63 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.405 $Y=0.126 $X2=0.414 $Y2=0.135
r78 60 62 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.126 $X2=0.405 $Y2=0.098
r79 59 61 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.07
r80 56 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.198 $X2=0.099 $Y2=0.198
r81 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.198 $X2=0.09 $Y2=0.198
r82 54 55 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.039
+ $Y=0.198 $X2=0.072 $Y2=0.198
r83 52 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.198 $X2=0.099 $Y2=0.198
r84 50 54 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.198 $X2=0.039 $Y2=0.198
r85 48 49 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.339
+ $Y=0.036 $X2=0.3675 $Y2=0.036
r86 47 48 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.339 $Y2=0.036
r87 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r88 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r89 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r90 42 43 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.2 $Y2=0.036
r91 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r92 40 41 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.036 $X2=0.18 $Y2=0.036
r93 39 40 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.176 $Y2=0.036
r94 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r95 37 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.126 $Y2=0.036
r96 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r97 34 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.234 $Y2=0.036
r98 34 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.2 $Y2=0.036
r99 31 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.072 $Y2=0.036
r100 29 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.054 $Y2=0.036
r101 28 59 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r102 28 49 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.3675 $Y2=0.036
r103 26 27 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.164
r104 25 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.189 $X2=0.036 $Y2=0.198
r105 25 27 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.027 $Y2=0.164
r106 24 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r107 24 26 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r108 23 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.198
+ $X2=0.108 $Y2=0.198
r109 20 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r110 19 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r111 18 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r112 15 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.054 $X2=0.216 $Y2=0.054
r113 14 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.054 $X2=0.216 $Y2=0.054
r114 12 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r115 9 12 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r116 5 65 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r117 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r118 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AO221X1_ASAP7_75T_L%Y 1 6 13 21 22 23 VSS
c6 35 VSS 0.00260752f $X=0.504 $Y=0.234
c7 34 VSS 0.00278493f $X=0.513 $Y=0.234
c8 29 VSS 0.00183949f $X=0.486 $Y=0.234
c9 27 VSS 2.98008e-19 $X=0.513 $Y=0.216
c10 26 VSS 8.34402e-19 $X=0.513 $Y=0.207
c11 25 VSS 0.00106207f $X=0.513 $Y=0.189
c12 23 VSS 7.45333e-19 $X=0.513 $Y=0.144
c13 22 VSS 0.00346118f $X=0.513 $Y=0.126
c14 21 VSS 0.00126998f $X=0.509 $Y=0.1475
c15 19 VSS 7.30208e-19 $X=0.513 $Y=0.225
c16 14 VSS 0.00645609f $X=0.486 $Y=0.036
c17 13 VSS 0.00284415f $X=0.486 $Y=0.036
c18 11 VSS 0.00571562f $X=0.504 $Y=0.036
c19 9 VSS 0.00682422f $X=0.484 $Y=0.2025
c20 4 VSS 3.19577e-19 $X=0.484 $Y=0.0675
r21 35 36 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.5085 $Y2=0.234
r22 34 36 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.234 $X2=0.5085 $Y2=0.234
r23 29 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.504 $Y2=0.234
r24 26 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.207 $X2=0.513 $Y2=0.216
r25 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.513 $Y2=0.207
r26 24 25 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.164 $X2=0.513 $Y2=0.189
r27 22 23 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.126 $X2=0.513 $Y2=0.144
r28 21 24 1.12037 $w=1.8e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.1475 $X2=0.513 $Y2=0.164
r29 21 23 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.1475 $X2=0.513 $Y2=0.144
r30 19 34 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.234
r31 19 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.216
r32 18 22 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.126
r33 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036 $X2=0.486
+ $Y2=0.036
r34 11 18 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.036 $X2=0.513 $Y2=0.045
r35 11 13 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.486 $Y2=0.036
r36 9 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r37 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.2025 $X2=0.484 $Y2=0.2025
r38 4 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0675 $X2=0.486 $Y2=0.036
r39 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.0675 $X2=0.484 $Y2=0.0675
.ends


* END of "./AO221x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO221x1_ASAP7_75t_L  VSS VDD B1 B2 C A1 A2 Y
* 
* Y	Y
* A2	A2
* A1	A1
* C	C
* B2	B2
* B1	B1
M0 noxref_12 N_B1_M0_g N_8_M0_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 VSS N_B2_M1_g noxref_12 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 N_8_M2_d N_C_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 noxref_13 N_A1_M3_g N_8_M3_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 VSS N_A2_M4_g noxref_13 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.027
M5 N_Y_M5_d N_8_M5_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M6 N_8_M6_d N_B1_M6_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 noxref_9 N_B2_M7_g N_8_M7_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 noxref_10 N_C_M8_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 VDD N_A1_M9_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 noxref_10 N_A2_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_Y_M11_d N_8_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "AO221x1_ASAP7_75t_L.pex.sp.AO221X1_ASAP7_75T_L.pxi"
* BEGIN of "./AO221x1_ASAP7_75t_L.pex.sp.AO221X1_ASAP7_75T_L.pxi"
* File: AO221x1_ASAP7_75t_L.pex.sp.AO221X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:03:34 2017
* 
x_PM_AO221X1_ASAP7_75T_L%B1 N_B1_M0_g N_B1_c_2_p N_B1_M6_g N_B1_c_3_p B1 VSS
+ PM_AO221X1_ASAP7_75T_L%B1
x_PM_AO221X1_ASAP7_75T_L%B2 N_B2_M1_g N_B2_c_13_n N_B2_M7_g B2 VSS
+ PM_AO221X1_ASAP7_75T_L%B2
x_PM_AO221X1_ASAP7_75T_L%C N_C_M2_g N_C_c_25_n N_C_M8_g C VSS
+ PM_AO221X1_ASAP7_75T_L%C
x_PM_AO221X1_ASAP7_75T_L%A1 N_A1_M3_g N_A1_c_36_n N_A1_M9_g N_A1_c_37_n A1 VSS
+ PM_AO221X1_ASAP7_75T_L%A1
x_PM_AO221X1_ASAP7_75T_L%A2 N_A2_M4_g N_A2_c_48_n N_A2_M10_g A2 N_A2_c_54_p VSS
+ PM_AO221X1_ASAP7_75T_L%A2
x_PM_AO221X1_ASAP7_75T_L%8 N_8_M5_g N_8_c_90_p N_8_M11_g N_8_M0_s N_8_c_55_n
+ N_8_M3_s N_8_M2_d N_8_c_63_n N_8_M7_s N_8_M6_d N_8_c_74_p N_8_c_56_n
+ N_8_c_87_p N_8_c_57_n N_8_c_61_n N_8_c_64_n N_8_c_83_p N_8_c_67_n N_8_c_85_p
+ N_8_c_69_n N_8_c_82_p N_8_c_78_p N_8_c_72_p N_8_c_59_n N_8_c_89_p N_8_c_71_n
+ N_8_c_88_p VSS PM_AO221X1_ASAP7_75T_L%8
x_PM_AO221X1_ASAP7_75T_L%Y N_Y_M5_d N_Y_M11_d N_Y_c_92_n Y N_Y_c_95_n N_Y_c_96_n
+ VSS PM_AO221X1_ASAP7_75T_L%Y
cc_1 N_B1_M0_g N_B2_M1_g 0.00364065f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_B1_c_2_p N_B2_c_13_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_B1_c_3_p B2 0.00484691f $X=0.081 $Y=0.135 $X2=0.133 $Y2=0.109
cc_4 N_B1_M0_g N_C_M2_g 2.6588e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 N_B1_c_3_p N_8_c_55_n 3.87865e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_6 N_B1_c_3_p N_8_c_56_n 0.00441847f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_7 N_B1_M0_g N_8_c_57_n 2.64276e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_8 N_B1_c_3_p N_8_c_57_n 0.00124805f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_B1_M0_g N_8_c_59_n 2.68514e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_10 N_B1_c_3_p N_8_c_59_n 0.00121543f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 VSS N_B1_M0_g 2.38303e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_12 N_B2_M1_g N_C_M2_g 0.0032267f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_13 N_B2_c_13_n N_C_c_25_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 B2 C 0.00456406f $X=0.133 $Y=0.109 $X2=0.081 $Y2=0.135
cc_15 N_B2_M1_g N_A1_M3_g 2.60137e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_16 N_B2_M1_g N_8_c_61_n 2.64276e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_17 B2 N_8_c_61_n 0.00124805f $X=0.133 $Y=0.109 $X2=0 $Y2=0
cc_18 VSS N_B2_M1_g 3.57119e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_19 VSS B2 5.37372e-19 $X=0.133 $Y=0.109 $X2=0 $Y2=0
cc_20 N_C_M2_g N_A1_M3_g 0.00346636f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_21 N_C_c_25_n N_A1_c_36_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 C N_A1_c_37_n 0.00456406f $X=0.188 $Y=0.123 $X2=0.081 $Y2=0.135
cc_23 N_C_M2_g N_A2_M4_g 2.54394e-19 $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_24 C N_8_c_63_n 3.31541e-19 $X=0.188 $Y=0.123 $X2=0 $Y2=0
cc_25 N_C_M2_g N_8_c_64_n 2.56935e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_26 C N_8_c_64_n 0.00123064f $X=0.188 $Y=0.123 $X2=0 $Y2=0
cc_27 N_A1_M3_g N_A2_M4_g 0.00310323f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_28 N_A1_c_36_n N_A2_c_48_n 9.33263e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_29 N_A1_c_37_n A2 0.00484283f $X=0.243 $Y=0.135 $X2=0.133 $Y2=0.109
cc_30 N_A1_c_37_n N_8_c_63_n 3.87865e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 N_A1_M3_g N_8_c_67_n 2.64276e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_32 N_A1_c_37_n N_8_c_67_n 0.00124805f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_33 VSS N_A1_M3_g 3.62029e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_34 VSS N_A1_c_37_n 0.0012322f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_35 N_A2_M4_g N_8_c_69_n 2.64276e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_36 A2 N_8_c_69_n 0.00124805f $X=0.295 $Y=0.123 $X2=0 $Y2=0
cc_37 A2 N_8_c_71_n 0.00123483f $X=0.295 $Y=0.123 $X2=0 $Y2=0
cc_38 VSS N_A2_M4_g 3.62029e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_39 VSS N_A2_c_54_p 0.0012322f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_40 VSS N_8_c_72_p 2.47657e-19 $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.054
cc_41 VSS N_8_c_55_n 9.76646e-19 $X=0.056 $Y=0.054 $X2=0.081 $Y2=0.135
cc_42 VSS N_8_c_74_p 0.00371671f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_43 VSS N_8_c_56_n 3.97918e-19 $X=0.027 $Y=0.164 $X2=0.081 $Y2=0.135
cc_44 VSS N_8_c_72_p 0.00263302f $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.135
cc_45 VSS N_8_c_74_p 0.00333296f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_46 VSS N_8_c_78_p 4.57757e-19 $X=0.108 $Y=0.198 $X2=0.081 $Y2=0.135
cc_47 VSS N_8_c_74_p 0.00250965f $X=0.108 $Y=0.2025 $X2=0 $Y2=0
cc_48 VSS N_8_c_72_p 0.00752628f $X=0.072 $Y=0.198 $X2=0 $Y2=0
cc_49 VSS N_8_c_63_n 9.98826e-19 $X=0.216 $Y=0.054 $X2=0.081 $Y2=0.135
cc_50 VSS N_8_c_82_p 2.77965e-19 $X=0.339 $Y=0.036 $X2=0 $Y2=0
cc_51 VSS N_8_c_83_p 2.77965e-19 $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_52 VSS N_8_c_78_p 3.01089e-19 $X=0.108 $Y=0.198 $X2=0 $Y2=0
cc_53 VSS N_8_c_85_p 2.77965e-19 $X=0.288 $Y=0.036 $X2=0 $Y2=0
cc_54 N_8_M5_g N_Y_c_92_n 3.47719e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.148
cc_55 N_8_c_87_p N_Y_c_92_n 4.96595e-19 $X=0.396 $Y=0.036 $X2=0.081 $Y2=0.148
cc_56 N_8_c_88_p N_Y_c_92_n 2.74073e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.148
cc_57 N_8_c_89_p N_Y_c_95_n 7.5881e-19 $X=0.405 $Y=0.07 $X2=0 $Y2=0
cc_58 N_8_c_90_p N_Y_c_96_n 3.14625e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_59 N_8_c_88_p N_Y_c_96_n 0.00105849f $X=0.459 $Y=0.135 $X2=0 $Y2=0

* END of "./AO221x1_ASAP7_75t_L.pex.sp.AO221X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO221x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:03:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO221x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO221x2_ASAP7_75t_L.pex.sp.pex"
* File: AO221x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:03:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO221X2_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c11 10 VSS 6.95749e-19 $X=0.081 $Y=0.135
c12 5 VSS 0.00170784f $X=0.081 $Y=0.135
c13 2 VSS 0.0655264f $X=0.081 $Y=0.054
r14 10 14 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.148
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO221X2_ASAP7_75T_L%B2 2 5 7 10 VSS
c11 10 VSS 0.00105185f $X=0.133 $Y=0.109
c12 5 VSS 0.00114017f $X=0.135 $Y=0.135
c13 2 VSS 0.0608869f $X=0.135 $Y=0.054
r14 10 13 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.109 $X2=0.135 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO221X2_ASAP7_75T_L%C 2 5 7 10 VSS
c11 10 VSS 0.00138457f $X=0.188 $Y=0.123
c12 5 VSS 0.00120688f $X=0.189 $Y=0.135
c13 2 VSS 0.0599046f $X=0.189 $Y=0.054
r14 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.123 $X2=0.189 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO221X2_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c12 10 VSS 6.84433e-19 $X=0.243 $Y=0.135
c13 5 VSS 0.00114323f $X=0.243 $Y=0.135
c14 2 VSS 0.0596104f $X=0.243 $Y=0.054
r15 10 14 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.151
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO221X2_ASAP7_75T_L%A2 2 5 7 10 13 VSS
c9 13 VSS 5.09476e-19 $X=0.297 $Y=0.135
c10 10 VSS 7.94635e-19 $X=0.295 $Y=0.123
c11 5 VSS 0.00212633f $X=0.297 $Y=0.135
c12 2 VSS 0.0616967f $X=0.297 $Y=0.054
r13 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.123 $X2=0.297 $Y2=0.135
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO221X2_ASAP7_75T_L%8 2 7 10 13 15 17 20 22 23 26 27 28 31 35 36 45
+ 47 50 52 53 54 55 56 60 63 64 69 70 73 VSS
c45 73 VSS 0.00307769f $X=0.459 $Y=0.135
c46 71 VSS 0.00126105f $X=0.414 $Y=0.135
c47 70 VSS 0.00149017f $X=0.405 $Y=0.098
c48 69 VSS 0.00211517f $X=0.405 $Y=0.07
c49 68 VSS 0.00108523f $X=0.405 $Y=0.126
c50 65 VSS 1.45514e-19 $X=0.099 $Y=0.198
c51 64 VSS 8.46035e-21 $X=0.09 $Y=0.198
c52 63 VSS 4.76765e-19 $X=0.072 $Y=0.198
c53 62 VSS 1.91267e-19 $X=0.039 $Y=0.198
c54 60 VSS 5.70579e-19 $X=0.108 $Y=0.198
c55 58 VSS 0.00193008f $X=0.036 $Y=0.198
c56 57 VSS 0.00395192f $X=0.3675 $Y=0.036
c57 56 VSS 0.00611566f $X=0.339 $Y=0.036
c58 55 VSS 0.00146362f $X=0.306 $Y=0.036
c59 54 VSS 0.00368202f $X=0.288 $Y=0.036
c60 53 VSS 0.00146362f $X=0.252 $Y=0.036
c61 52 VSS 0.00331014f $X=0.234 $Y=0.036
c62 51 VSS 1.99947e-19 $X=0.2 $Y=0.036
c63 50 VSS 0.00142296f $X=0.198 $Y=0.036
c64 49 VSS 4.31197e-19 $X=0.18 $Y=0.036
c65 48 VSS 0.00564793f $X=0.176 $Y=0.036
c66 47 VSS 0.00146362f $X=0.144 $Y=0.036
c67 46 VSS 0.00345019f $X=0.126 $Y=0.036
c68 45 VSS 0.00146362f $X=0.09 $Y=0.036
c69 44 VSS 0.00353842f $X=0.072 $Y=0.036
c70 37 VSS 0.00340187f $X=0.036 $Y=0.036
c71 36 VSS 0.00653563f $X=0.396 $Y=0.036
c72 35 VSS 0.00423691f $X=0.027 $Y=0.164
c73 34 VSS 9.59589e-19 $X=0.027 $Y=0.07
c74 33 VSS 0.00112176f $X=0.027 $Y=0.189
c75 31 VSS 0.00233317f $X=0.108 $Y=0.2025
c76 27 VSS 5.91014e-19 $X=0.125 $Y=0.2025
c77 26 VSS 0.00607665f $X=0.216 $Y=0.054
c78 22 VSS 5.19811e-19 $X=0.233 $Y=0.054
c79 20 VSS 0.00319205f $X=0.056 $Y=0.054
c80 17 VSS 2.6657e-19 $X=0.071 $Y=0.054
c81 13 VSS 0.00558302f $X=0.513 $Y=0.135
c82 10 VSS 0.0641916f $X=0.513 $Y=0.0675
c83 2 VSS 0.0645799f $X=0.459 $Y=0.0675
r84 71 73 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.135 $X2=0.459 $Y2=0.135
r85 69 70 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.07 $X2=0.405 $Y2=0.098
r86 68 71 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.405 $Y=0.126 $X2=0.414 $Y2=0.135
r87 68 70 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.126 $X2=0.405 $Y2=0.098
r88 67 69 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.07
r89 64 65 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.198 $X2=0.099 $Y2=0.198
r90 63 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.198 $X2=0.09 $Y2=0.198
r91 62 63 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.039
+ $Y=0.198 $X2=0.072 $Y2=0.198
r92 60 65 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.198 $X2=0.099 $Y2=0.198
r93 58 62 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.198 $X2=0.039 $Y2=0.198
r94 56 57 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.339
+ $Y=0.036 $X2=0.3675 $Y2=0.036
r95 55 56 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.339 $Y2=0.036
r96 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r97 53 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r98 52 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r99 50 51 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.2 $Y2=0.036
r100 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r101 48 49 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.036 $X2=0.18 $Y2=0.036
r102 47 48 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.176 $Y2=0.036
r103 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r104 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.126 $Y2=0.036
r105 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r106 42 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.234 $Y2=0.036
r107 42 51 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.2 $Y2=0.036
r108 39 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.072 $Y2=0.036
r109 37 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.054 $Y2=0.036
r110 36 67 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r111 36 57 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.3675 $Y2=0.036
r112 34 35 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.164
r113 33 58 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.189 $X2=0.036 $Y2=0.198
r114 33 35 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.027 $Y2=0.164
r115 32 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r116 32 34 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r117 31 60 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.198
+ $X2=0.108 $Y2=0.198
r118 28 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r119 27 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r120 26 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r121 23 26 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.054 $X2=0.216 $Y2=0.054
r122 22 26 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.054 $X2=0.216 $Y2=0.054
r123 20 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r124 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r125 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r126 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r127 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r128 5 73 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r129 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r130 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AO221X2_ASAP7_75T_L%Y 1 2 6 7 10 11 13 14 18 20 28 29 30 VSS
c14 34 VSS 8.50351e-19 $X=0.54 $Y=0.216
c15 33 VSS 0.00163777f $X=0.54 $Y=0.207
c16 32 VSS 0.00191308f $X=0.54 $Y=0.189
c17 30 VSS 5.47546e-19 $X=0.54 $Y=0.144
c18 29 VSS 0.00691258f $X=0.54 $Y=0.126
c19 28 VSS 0.00149354f $X=0.537 $Y=0.1475
c20 26 VSS 8.0311e-19 $X=0.54 $Y=0.225
c21 20 VSS 0.00178743f $X=0.486 $Y=0.234
c22 18 VSS 0.00906391f $X=0.531 $Y=0.234
c23 14 VSS 0.00902228f $X=0.486 $Y=0.036
c24 13 VSS 0.00273288f $X=0.486 $Y=0.036
c25 11 VSS 0.00893562f $X=0.531 $Y=0.036
c26 10 VSS 0.00904513f $X=0.486 $Y=0.2025
c27 6 VSS 5.58795e-19 $X=0.503 $Y=0.2025
c28 1 VSS 5.25448e-19 $X=0.503 $Y=0.0675
r29 33 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.207 $X2=0.54 $Y2=0.216
r30 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.189 $X2=0.54 $Y2=0.207
r31 31 32 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.164 $X2=0.54 $Y2=0.189
r32 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.126 $X2=0.54 $Y2=0.144
r33 28 31 1.12037 $w=1.8e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.1475 $X2=0.54 $Y2=0.164
r34 28 30 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.1475 $X2=0.54 $Y2=0.144
r35 26 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.225 $X2=0.54 $Y2=0.216
r36 25 29 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.045 $X2=0.54 $Y2=0.126
r37 18 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.531 $Y=0.234 $X2=0.54 $Y2=0.225
r38 18 20 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.531
+ $Y=0.234 $X2=0.486 $Y2=0.234
r39 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036 $X2=0.486
+ $Y2=0.036
r40 11 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.531 $Y=0.036 $X2=0.54 $Y2=0.045
r41 11 13 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.531
+ $Y=0.036 $X2=0.486 $Y2=0.036
r42 10 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r43 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.486 $Y2=0.2025
r44 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.2025 $X2=0.486 $Y2=0.2025
r45 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0675 $X2=0.486 $Y2=0.036
r46 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.0675 $X2=0.486 $Y2=0.0675
r47 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0675 $X2=0.486 $Y2=0.0675
.ends


* END of "./AO221x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO221x2_ASAP7_75t_L  VSS VDD B1 B2 C A1 A2 Y
* 
* Y	Y
* A2	A2
* A1	A1
* C	C
* B2	B2
* B1	B1
M0 noxref_12 N_B1_M0_g N_8_M0_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 VSS N_B2_M1_g noxref_12 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 N_8_M2_d N_C_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 noxref_13 N_A1_M3_g N_8_M3_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 VSS N_A2_M4_g noxref_13 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.027
M5 N_Y_M5_d N_8_M5_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M6 N_Y_M6_d N_8_M6_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M7 N_8_M7_d N_B1_M7_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M8 noxref_9 N_B2_M8_g N_8_M8_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M9 noxref_10 N_C_M9_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M10 VDD N_A1_M10_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M11 noxref_10 N_A2_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M12 N_Y_M12_d N_8_M12_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M13 N_Y_M13_d N_8_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
*
* 
* .include "AO221x2_ASAP7_75t_L.pex.sp.AO221X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO221x2_ASAP7_75t_L.pex.sp.AO221X2_ASAP7_75T_L.pxi"
* File: AO221x2_ASAP7_75t_L.pex.sp.AO221X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:03:56 2017
* 
x_PM_AO221X2_ASAP7_75T_L%B1 N_B1_M0_g N_B1_c_2_p N_B1_M7_g N_B1_c_3_p B1 VSS
+ PM_AO221X2_ASAP7_75T_L%B1
x_PM_AO221X2_ASAP7_75T_L%B2 N_B2_M1_g N_B2_c_13_n N_B2_M8_g B2 VSS
+ PM_AO221X2_ASAP7_75T_L%B2
x_PM_AO221X2_ASAP7_75T_L%C N_C_M2_g N_C_c_25_n N_C_M9_g C VSS
+ PM_AO221X2_ASAP7_75T_L%C
x_PM_AO221X2_ASAP7_75T_L%A1 N_A1_M3_g N_A1_c_36_n N_A1_M10_g N_A1_c_37_n A1 VSS
+ PM_AO221X2_ASAP7_75T_L%A1
x_PM_AO221X2_ASAP7_75T_L%A2 N_A2_M4_g N_A2_c_48_n N_A2_M11_g A2 N_A2_c_54_p VSS
+ PM_AO221X2_ASAP7_75T_L%A2
x_PM_AO221X2_ASAP7_75T_L%8 N_8_M5_g N_8_M12_g N_8_M6_g N_8_c_86_p N_8_M13_g
+ N_8_M0_s N_8_c_55_n N_8_M3_s N_8_M2_d N_8_c_63_n N_8_M8_s N_8_M7_d N_8_c_74_p
+ N_8_c_56_n N_8_c_92_p N_8_c_57_n N_8_c_61_n N_8_c_64_n N_8_c_83_p N_8_c_67_n
+ N_8_c_85_p N_8_c_69_n N_8_c_82_p N_8_c_78_p N_8_c_72_p N_8_c_59_n N_8_c_98_p
+ N_8_c_71_n N_8_c_93_p VSS PM_AO221X2_ASAP7_75T_L%8
x_PM_AO221X2_ASAP7_75T_L%Y N_Y_M6_d N_Y_M5_d N_Y_M13_d N_Y_M12_d N_Y_c_102_n
+ N_Y_c_103_n N_Y_c_104_n N_Y_c_108_n N_Y_c_109_n N_Y_c_110_n Y N_Y_c_111_n
+ N_Y_c_113_n VSS PM_AO221X2_ASAP7_75T_L%Y
cc_1 N_B1_M0_g N_B2_M1_g 0.00364065f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_B1_c_2_p N_B2_c_13_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_B1_c_3_p B2 0.00484691f $X=0.081 $Y=0.135 $X2=0.133 $Y2=0.109
cc_4 N_B1_M0_g N_C_M2_g 2.6588e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 N_B1_c_3_p N_8_c_55_n 3.87865e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_6 N_B1_c_3_p N_8_c_56_n 0.00441847f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_7 N_B1_M0_g N_8_c_57_n 2.64276e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_8 N_B1_c_3_p N_8_c_57_n 0.00124805f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_B1_M0_g N_8_c_59_n 2.68514e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_10 N_B1_c_3_p N_8_c_59_n 0.00121543f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 VSS N_B1_M0_g 2.38303e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_12 N_B2_M1_g N_C_M2_g 0.0032267f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_13 N_B2_c_13_n N_C_c_25_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 B2 C 0.00456406f $X=0.133 $Y=0.109 $X2=0.081 $Y2=0.135
cc_15 N_B2_M1_g N_A1_M3_g 2.60137e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_16 N_B2_M1_g N_8_c_61_n 2.64276e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_17 B2 N_8_c_61_n 0.00124805f $X=0.133 $Y=0.109 $X2=0 $Y2=0
cc_18 VSS N_B2_M1_g 3.57119e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_19 VSS B2 5.37372e-19 $X=0.133 $Y=0.109 $X2=0 $Y2=0
cc_20 N_C_M2_g N_A1_M3_g 0.00346636f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_21 N_C_c_25_n N_A1_c_36_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 C N_A1_c_37_n 0.00456406f $X=0.188 $Y=0.123 $X2=0.081 $Y2=0.135
cc_23 N_C_M2_g N_A2_M4_g 2.54394e-19 $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_24 C N_8_c_63_n 3.31541e-19 $X=0.188 $Y=0.123 $X2=0 $Y2=0
cc_25 N_C_M2_g N_8_c_64_n 2.56935e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_26 C N_8_c_64_n 0.00123064f $X=0.188 $Y=0.123 $X2=0 $Y2=0
cc_27 N_A1_M3_g N_A2_M4_g 0.00310323f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_28 N_A1_c_36_n N_A2_c_48_n 9.33263e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_29 N_A1_c_37_n A2 0.00484283f $X=0.243 $Y=0.135 $X2=0.133 $Y2=0.109
cc_30 N_A1_c_37_n N_8_c_63_n 3.87865e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 N_A1_M3_g N_8_c_67_n 2.64276e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_32 N_A1_c_37_n N_8_c_67_n 0.00124805f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_33 VSS N_A1_M3_g 3.62029e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_34 VSS N_A1_c_37_n 0.0012322f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_35 N_A2_M4_g N_8_c_69_n 2.64276e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_36 A2 N_8_c_69_n 0.00124805f $X=0.295 $Y=0.123 $X2=0 $Y2=0
cc_37 A2 N_8_c_71_n 0.00123483f $X=0.295 $Y=0.123 $X2=0 $Y2=0
cc_38 VSS N_A2_M4_g 3.62029e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_39 VSS N_A2_c_54_p 0.0012322f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_40 VSS N_8_c_72_p 2.47657e-19 $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.054
cc_41 VSS N_8_c_55_n 9.76646e-19 $X=0.056 $Y=0.054 $X2=0.081 $Y2=0.135
cc_42 VSS N_8_c_74_p 0.00371671f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_43 VSS N_8_c_56_n 3.97918e-19 $X=0.027 $Y=0.164 $X2=0.081 $Y2=0.135
cc_44 VSS N_8_c_72_p 0.00263302f $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.135
cc_45 VSS N_8_c_74_p 0.00333296f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_46 VSS N_8_c_78_p 4.57757e-19 $X=0.108 $Y=0.198 $X2=0.081 $Y2=0.135
cc_47 VSS N_8_c_74_p 0.00250965f $X=0.108 $Y=0.2025 $X2=0 $Y2=0
cc_48 VSS N_8_c_72_p 0.00752628f $X=0.072 $Y=0.198 $X2=0 $Y2=0
cc_49 VSS N_8_c_63_n 9.98826e-19 $X=0.216 $Y=0.054 $X2=0.081 $Y2=0.135
cc_50 VSS N_8_c_82_p 2.77965e-19 $X=0.339 $Y=0.036 $X2=0 $Y2=0
cc_51 VSS N_8_c_83_p 2.77965e-19 $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_52 VSS N_8_c_78_p 3.01089e-19 $X=0.108 $Y=0.198 $X2=0 $Y2=0
cc_53 VSS N_8_c_85_p 2.77965e-19 $X=0.288 $Y=0.036 $X2=0 $Y2=0
cc_54 N_8_c_86_p N_Y_M6_d 3.8044e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.054
cc_55 N_8_c_86_p N_Y_M13_d 3.8044e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_56 N_8_c_86_p N_Y_c_102_n 8.00061e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.135
cc_57 N_8_M6_g N_Y_c_103_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_58 N_8_M5_g N_Y_c_104_n 3.49779e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.148
cc_59 N_8_c_86_p N_Y_c_104_n 5.88586e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.148
cc_60 N_8_c_92_p N_Y_c_104_n 5.0963e-19 $X=0.396 $Y=0.036 $X2=0.081 $Y2=0.148
cc_61 N_8_c_93_p N_Y_c_104_n 2.47393e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.148
cc_62 N_8_c_86_p N_Y_c_108_n 8.00061e-19 $X=0.513 $Y=0.135 $X2=0.076 $Y2=0.148
cc_63 N_8_M6_g N_Y_c_109_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_8_c_86_p N_Y_c_110_n 5.35675e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_65 N_8_c_86_p N_Y_c_111_n 3.51153e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_66 N_8_c_98_p N_Y_c_111_n 4.82822e-19 $X=0.405 $Y=0.07 $X2=0 $Y2=0
cc_67 N_8_c_93_p N_Y_c_113_n 4.99147e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0

* END of "./AO221x2_ASAP7_75t_L.pex.sp.AO221X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO222x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:04:19 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO222x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO222x2_ASAP7_75t_L.pex.sp.pex"
* File: AO222x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:04:19 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO222X2_ASAP7_75T_L%A1 2 5 8 11 13 25 VSS
c14 29 VSS 0.00199488f $X=0.081 $Y=0.135
c15 25 VSS 0.0243989f $X=0.061 $Y=0.1335
c16 11 VSS 0.00514703f $X=0.135 $Y=0.135
c17 8 VSS 0.0623423f $X=0.135 $Y=0.0675
c18 2 VSS 0.067361f $X=0.081 $Y=0.135
r19 25 29 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.061
+ $Y=0.135 $X2=0.081 $Y2=0.135
r20 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r21 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r22 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r23 2 29 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r24 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
.ends

.subckt PM_AO222X2_ASAP7_75T_L%A2 2 7 10 13 22 VSS
c16 22 VSS 0.0071796f $X=0.242 $Y=0.1365
c17 10 VSS 0.0735665f $X=0.243 $Y=0.135
c18 2 VSS 0.0630916f $X=0.189 $Y=0.0675
r19 10 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r20 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r21 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO222X2_ASAP7_75T_L%B2 2 5 8 11 13 23 25 VSS
c22 25 VSS 0.00136606f $X=0.405 $Y=0.135
c23 23 VSS 0.00745695f $X=0.385 $Y=0.1335
c24 11 VSS 0.00767224f $X=0.459 $Y=0.135
c25 8 VSS 0.0648902f $X=0.459 $Y=0.0675
c26 2 VSS 0.0682653f $X=0.405 $Y=0.135
r27 23 25 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.385
+ $Y=0.135 $X2=0.405 $Y2=0.135
r28 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r29 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r30 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r31 2 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r32 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
.ends

.subckt PM_AO222X2_ASAP7_75T_L%B1 2 7 10 13 22 VSS
c21 22 VSS 0.00344167f $X=0.512 $Y=0.1415
c22 10 VSS 0.0731244f $X=0.567 $Y=0.135
c23 2 VSS 0.0637664f $X=0.513 $Y=0.0675
r24 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r25 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r26 5 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r27 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r28 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AO222X2_ASAP7_75T_L%C1 2 5 8 11 13 22 VSS
c18 22 VSS 0.00410504f $X=0.729 $Y=0.1405
c19 11 VSS 0.00438535f $X=0.783 $Y=0.135
c20 8 VSS 0.0641408f $X=0.783 $Y=0.0675
c21 2 VSS 0.0685112f $X=0.729 $Y=0.135
r22 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.135 $X2=0.783 $Y2=0.2025
r23 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0675 $X2=0.783 $Y2=0.135
r24 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.135 $X2=0.783 $Y2=0.135
r25 2 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.729 $Y=0.135 $X2=0.729
+ $Y2=0.135
r26 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.135 $X2=0.729 $Y2=0.2025
.ends

.subckt PM_AO222X2_ASAP7_75T_L%C2 2 7 10 13 21 VSS
c23 21 VSS 0.00528042f $X=0.904 $Y=0.1335
c24 10 VSS 0.0755161f $X=0.891 $Y=0.135
c25 2 VSS 0.0648902f $X=0.837 $Y=0.0675
r26 17 21 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.135 $X2=0.904 $Y2=0.135
r27 10 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.135 $X2=0.891
+ $Y2=0.135
r28 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.135 $X2=0.891 $Y2=0.2025
r29 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.837
+ $Y=0.135 $X2=0.891 $Y2=0.135
r30 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.2025
r31 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.0675 $X2=0.837 $Y2=0.135
.ends

.subckt PM_AO222X2_ASAP7_75T_L%9 2 7 10 13 15 17 22 27 32 33 36 37 38 41 42 44
+ 45 51 52 53 54 55 56 57 58 59 62 63 64 65 66 67 69 77 78 80 82 85 87 91 94 VSS
c84 94 VSS 4.03344e-19 $X=0.999 $Y=0.135
c85 91 VSS 0.00316031f $X=1.052 $Y=0.135
c86 88 VSS 5.62236e-19 $X=0.999 $Y=0.216
c87 87 VSS 0.00112681f $X=0.999 $Y=0.207
c88 86 VSS 0.00120599f $X=0.999 $Y=0.189
c89 85 VSS 0.00159654f $X=0.999 $Y=0.171
c90 84 VSS 5.31001e-19 $X=0.999 $Y=0.225
c91 82 VSS 0.00186623f $X=0.999 $Y=0.0945
c92 81 VSS 0.00109324f $X=0.999 $Y=0.063
c93 80 VSS 0.00134208f $X=0.999 $Y=0.126
c94 78 VSS 0.00228373f $X=0.954 $Y=0.234
c95 77 VSS 0.0155159f $X=0.932 $Y=0.234
c96 69 VSS 0.00757627f $X=0.99 $Y=0.234
c97 68 VSS 0.00208651f $X=0.972 $Y=0.036
c98 67 VSS 0.00329905f $X=0.954 $Y=0.036
c99 66 VSS 0.00332626f $X=0.917 $Y=0.036
c100 65 VSS 0.0158447f $X=0.877 $Y=0.036
c101 64 VSS 0.00311606f $X=0.738 $Y=0.036
c102 63 VSS 0.0184488f $X=0.701 $Y=0.036
c103 62 VSS 0.00450651f $X=0.756 $Y=0.036
c104 59 VSS 7.78824e-19 $X=0.531 $Y=0.036
c105 58 VSS 0.00308768f $X=0.522 $Y=0.036
c106 57 VSS 0.0095766f $X=0.485 $Y=0.036
c107 56 VSS 0.00491144f $X=0.419 $Y=0.036
c108 55 VSS 0.00348601f $X=0.36 $Y=0.036
c109 54 VSS 0.00834035f $X=0.323 $Y=0.036
c110 53 VSS 0.00495294f $X=0.252 $Y=0.036
c111 52 VSS 0.0119456f $X=0.215 $Y=0.036
c112 51 VSS 0.00439671f $X=0.54 $Y=0.036
c113 45 VSS 0.00454982f $X=0.108 $Y=0.036
c114 44 VSS 0.00114698f $X=0.108 $Y=0.036
c115 42 VSS 0.00496487f $X=0.99 $Y=0.036
c116 41 VSS 0.00495547f $X=0.864 $Y=0.2025
c117 37 VSS 5.86873e-19 $X=0.881 $Y=0.2025
c118 36 VSS 0.00297664f $X=0.756 $Y=0.2025
c119 32 VSS 6.4808e-19 $X=0.773 $Y=0.2025
c120 27 VSS 4.59792e-19 $X=0.773 $Y=0.0675
c121 25 VSS 4.59792e-19 $X=0.538 $Y=0.0675
c122 17 VSS 4.59792e-19 $X=0.125 $Y=0.0675
c123 13 VSS 0.0059175f $X=1.107 $Y=0.135
c124 10 VSS 0.0647446f $X=1.107 $Y=0.0675
c125 2 VSS 0.0652872f $X=1.053 $Y=0.0675
r126 89 94 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.008
+ $Y=0.135 $X2=0.999 $Y2=0.135
r127 89 91 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.008
+ $Y=0.135 $X2=1.052 $Y2=0.135
r128 87 88 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.207 $X2=0.999 $Y2=0.216
r129 86 87 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.189 $X2=0.999 $Y2=0.207
r130 85 86 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.171 $X2=0.999 $Y2=0.189
r131 84 88 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.225 $X2=0.999 $Y2=0.216
r132 83 94 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.144 $X2=0.999 $Y2=0.135
r133 83 85 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.144 $X2=0.999 $Y2=0.171
r134 81 82 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.063 $X2=0.999 $Y2=0.0945
r135 80 94 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.126 $X2=0.999 $Y2=0.135
r136 80 82 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.126 $X2=0.999 $Y2=0.0945
r137 79 81 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.045 $X2=0.999 $Y2=0.063
r138 77 78 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.932
+ $Y=0.234 $X2=0.954 $Y2=0.234
r139 75 77 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.932 $Y2=0.234
r140 71 75 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.864 $Y2=0.234
r141 69 84 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.99 $Y=0.234 $X2=0.999 $Y2=0.225
r142 69 78 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.99
+ $Y=0.234 $X2=0.954 $Y2=0.234
r143 67 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.036 $X2=0.972 $Y2=0.036
r144 66 67 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.917
+ $Y=0.036 $X2=0.954 $Y2=0.036
r145 65 66 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.877
+ $Y=0.036 $X2=0.917 $Y2=0.036
r146 63 64 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.701
+ $Y=0.036 $X2=0.738 $Y2=0.036
r147 61 65 8.21605 $w=1.8e-08 $l=1.21e-07 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.877 $Y2=0.036
r148 61 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.738 $Y2=0.036
r149 61 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036
+ $X2=0.756 $Y2=0.036
r150 58 59 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.531 $Y2=0.036
r151 57 58 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.485
+ $Y=0.036 $X2=0.522 $Y2=0.036
r152 56 57 4.48148 $w=1.8e-08 $l=6.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.419
+ $Y=0.036 $X2=0.485 $Y2=0.036
r153 55 56 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.419 $Y2=0.036
r154 54 55 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.323
+ $Y=0.036 $X2=0.36 $Y2=0.036
r155 53 54 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.323 $Y2=0.036
r156 52 53 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.215
+ $Y=0.036 $X2=0.252 $Y2=0.036
r157 50 63 10.9321 $w=1.8e-08 $l=1.61e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.701 $Y2=0.036
r158 50 59 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.531 $Y2=0.036
r159 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r160 44 52 7.26543 $w=1.8e-08 $l=1.07e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.215 $Y2=0.036
r161 44 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r162 42 79 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.99 $Y=0.036 $X2=0.999 $Y2=0.045
r163 42 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.99
+ $Y=0.036 $X2=0.972 $Y2=0.036
r164 41 75 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234
+ $X2=0.864 $Y2=0.234
r165 38 41 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2025 $X2=0.864 $Y2=0.2025
r166 37 41 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2025 $X2=0.864 $Y2=0.2025
r167 36 71 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234
+ $X2=0.756 $Y2=0.234
r168 33 36 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r169 32 36 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r170 30 62 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.756 $Y=0.0675 $X2=0.756 $Y2=0.036
r171 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.758 $Y2=0.0675
r172 25 51 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r173 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.538 $Y2=0.0675
r174 20 45 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.108 $Y=0.0675 $X2=0.108 $Y2=0.036
r175 17 20 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.11 $Y2=0.0675
r176 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.135 $X2=1.107 $Y2=0.2025
r177 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.0675 $X2=1.107 $Y2=0.135
r178 5 13 50 $w=2.2e-08 $l=5.5e-08 $layer=LIG $thickness=5e-08 $X=1.052 $Y=0.135
+ $X2=1.107 $Y2=0.135
r179 5 91 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.052 $Y=0.135 $X2=1.052
+ $Y2=0.135
r180 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.135 $X2=1.053 $Y2=0.2025
r181 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.0675 $X2=1.053 $Y2=0.135
.ends

.subckt PM_AO222X2_ASAP7_75T_L%Y 1 2 6 7 10 11 14 16 24 25 26 VSS
c13 28 VSS 0.0026303f $X=1.161 $Y=0.1845
c14 26 VSS 3.47847e-19 $X=1.161 $Y=0.13375
c15 25 VSS 0.0046845f $X=1.161 $Y=0.126
c16 24 VSS 4.26393e-19 $X=1.161 $Y=0.1415
c17 22 VSS 0.00236896f $X=1.161 $Y=0.225
c18 16 VSS 0.0145473f $X=1.152 $Y=0.234
c19 14 VSS 0.00931001f $X=1.08 $Y=0.036
c20 11 VSS 0.0145473f $X=1.152 $Y=0.036
c21 10 VSS 0.00914519f $X=1.08 $Y=0.2025
c22 6 VSS 5.72268e-19 $X=1.097 $Y=0.2025
c23 1 VSS 5.72268e-19 $X=1.097 $Y=0.0675
r24 27 28 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.144 $X2=1.161 $Y2=0.1845
r25 25 26 0.526235 $w=1.8e-08 $l=7.75e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.126 $X2=1.161 $Y2=0.13375
r26 24 27 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.1415 $X2=1.161 $Y2=0.144
r27 24 26 0.526235 $w=1.8e-08 $l=7.75e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.1415 $X2=1.161 $Y2=0.13375
r28 22 28 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.225 $X2=1.161 $Y2=0.1845
r29 21 25 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.045 $X2=1.161 $Y2=0.126
r30 16 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.152 $Y=0.234 $X2=1.161 $Y2=0.225
r31 16 18 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.152
+ $Y=0.234 $X2=1.08 $Y2=0.234
r32 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.036 $X2=1.08
+ $Y2=0.036
r33 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.152 $Y=0.036 $X2=1.161 $Y2=0.045
r34 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.152
+ $Y=0.036 $X2=1.08 $Y2=0.036
r35 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234 $X2=1.08
+ $Y2=0.234
r36 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2025 $X2=1.08 $Y2=0.2025
r37 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.097 $Y=0.2025 $X2=1.08 $Y2=0.2025
r38 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.08
+ $Y=0.0675 $X2=1.08 $Y2=0.036
r39 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.063
+ $Y=0.0675 $X2=1.08 $Y2=0.0675
r40 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.097
+ $Y=0.0675 $X2=1.08 $Y2=0.0675
.ends


* END of "./AO222x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO222x2_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 C1 C2 Y
* 
* Y	Y
* C2	C2
* C1	C1
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 noxref_13 N_A1_M0_g N_9_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M1 VSS N_A2_M1_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M2 noxref_14 N_B2_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M3 N_9_M3_d N_B1_M3_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M4 noxref_15 N_C1_M4_g N_9_M4_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.027
M5 VSS N_C2_M5_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.027
M6 N_Y_M6_d N_9_M6_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=1.043 $Y=0.027
M7 N_Y_M7_d N_9_M7_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=1.097 $Y=0.027
M8 noxref_10 N_A1_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M9 noxref_10 N_A1_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M10 noxref_10 N_A2_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M11 noxref_10 N_A2_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M12 noxref_11 N_B2_M12_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M13 noxref_11 N_B2_M13_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M14 noxref_11 N_B1_M14_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
M15 noxref_11 N_B1_M15_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M16 N_9_M16_d N_C1_M16_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.719 $Y=0.162
M17 N_9_M17_d N_C1_M17_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.773 $Y=0.162
M18 N_9_M18_d N_C2_M18_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.827 $Y=0.162
M19 N_9_M19_d N_C2_M19_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.881 $Y=0.162
M20 N_Y_M20_d N_9_M20_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.162
M21 N_Y_M21_d N_9_M21_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.162
*
* 
* .include "AO222x2_ASAP7_75t_L.pex.sp.AO222X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO222x2_ASAP7_75t_L.pex.sp.AO222X2_ASAP7_75T_L.pxi"
* File: AO222x2_ASAP7_75t_L.pex.sp.AO222X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:04:19 2017
* 
x_PM_AO222X2_ASAP7_75T_L%A1 N_A1_c_1_p N_A1_M8_g N_A1_M0_g N_A1_c_4_p N_A1_M9_g
+ A1 VSS PM_AO222X2_ASAP7_75T_L%A1
x_PM_AO222X2_ASAP7_75T_L%A2 N_A2_M1_g N_A2_M10_g N_A2_c_17_n N_A2_M11_g A2 VSS
+ PM_AO222X2_ASAP7_75T_L%A2
x_PM_AO222X2_ASAP7_75T_L%B2 N_B2_c_32_p N_B2_M12_g N_B2_M2_g N_B2_c_35_p
+ N_B2_M13_g B2 N_B2_c_40_p VSS PM_AO222X2_ASAP7_75T_L%B2
x_PM_AO222X2_ASAP7_75T_L%B1 N_B1_M3_g N_B1_M14_g N_B1_c_55_n N_B1_M15_g B1 VSS
+ PM_AO222X2_ASAP7_75T_L%B1
x_PM_AO222X2_ASAP7_75T_L%C1 N_C1_c_74_p N_C1_M16_g N_C1_M4_g N_C1_c_77_p
+ N_C1_M17_g C1 VSS PM_AO222X2_ASAP7_75T_L%C1
x_PM_AO222X2_ASAP7_75T_L%C2 N_C2_M5_g N_C2_M18_g N_C2_c_94_n N_C2_M19_g C2 VSS
+ PM_AO222X2_ASAP7_75T_L%C2
x_PM_AO222X2_ASAP7_75T_L%9 N_9_M6_g N_9_M20_g N_9_M7_g N_9_c_184_p N_9_M21_g
+ N_9_M0_s N_9_M3_d N_9_M4_s N_9_M17_d N_9_M16_d N_9_c_136_n N_9_M19_d N_9_M18_d
+ N_9_c_145_n N_9_c_189_p N_9_c_115_n N_9_c_117_n N_9_c_129_n N_9_c_119_n
+ N_9_c_122_n N_9_c_161_p N_9_c_124_n N_9_c_125_n N_9_c_128_n N_9_c_131_n
+ N_9_c_133_n N_9_c_137_n N_9_c_134_n N_9_c_139_n N_9_c_141_n N_9_c_148_n
+ N_9_c_150_n N_9_c_193_p N_9_c_143_n N_9_c_154_n N_9_c_155_n N_9_c_156_n
+ N_9_c_173_p N_9_c_180_p N_9_c_196_p N_9_c_157_n VSS PM_AO222X2_ASAP7_75T_L%9
x_PM_AO222X2_ASAP7_75T_L%Y N_Y_M7_d N_Y_M6_d N_Y_M21_d N_Y_M20_d N_Y_c_201_n
+ N_Y_c_202_n N_Y_c_205_n N_Y_c_206_n Y N_Y_c_209_n N_Y_c_211_n VSS
+ PM_AO222X2_ASAP7_75T_L%Y
cc_1 N_A1_c_1_p N_A2_M1_g 2.69148e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_2 N_A1_M0_g N_A2_M1_g 0.00323392f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A1_M0_g N_A2_c_17_n 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_4 N_A1_c_4_p N_A2_c_17_n 0.00163635f $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_5 N_A1_c_4_p N_9_c_115_n 5.21154e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_6 A1 N_9_c_115_n 8.46903e-19 $X=0.061 $Y=0.1335 $X2=0 $Y2=0
cc_7 N_A1_c_4_p N_9_c_117_n 8.0006e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_8 A1 N_9_c_117_n 0.00166117f $X=0.061 $Y=0.1335 $X2=0 $Y2=0
cc_9 N_A1_M0_g N_9_c_119_n 4.58656e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_10 VSS N_A1_c_4_p 3.80485e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_11 VSS N_A1_c_4_p 8.0006e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_12 VSS N_A1_c_4_p 5.20568e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_13 VSS A1 5.33049e-19 $X=0.061 $Y=0.1335 $X2=0 $Y2=0
cc_14 VSS N_A1_M0_g 4.58656e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 A2 B2 0.00272345f $X=0.242 $Y=0.1365 $X2=0 $Y2=0
cc_16 N_A2_M1_g N_9_c_119_n 4.58656e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_17 N_A2_c_17_n N_9_c_119_n 4.88232e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_18 N_A2_c_17_n N_9_c_122_n 2.38303e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_19 A2 N_9_c_122_n 0.00374964f $X=0.242 $Y=0.1365 $X2=0 $Y2=0
cc_20 VSS N_A2_c_17_n 3.80455e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_21 VSS N_A2_c_17_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_22 VSS A2 0.00161606f $X=0.242 $Y=0.1365 $X2=0.135 $Y2=0.135
cc_23 VSS N_A2_M1_g 4.58656e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 VSS N_A2_c_17_n 3.83955e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_25 VSS N_A2_c_17_n 2.34993e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_26 VSS A2 0.00372802f $X=0.242 $Y=0.1365 $X2=0.135 $Y2=0.135
cc_27 N_B2_c_32_p N_B1_M3_g 2.74891e-19 $X=0.405 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_28 N_B2_M2_g N_B1_M3_g 0.00372052f $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_29 N_B2_M2_g N_B1_c_55_n 3.09654e-19 $X=0.459 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_30 N_B2_c_35_p N_B1_c_55_n 0.00135537f $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.135
cc_31 B2 B1 3.69601e-19 $X=0.385 $Y=0.1335 $X2=0.242 $Y2=0.1365
cc_32 B2 N_9_c_124_n 0.00375203f $X=0.385 $Y=0.1335 $X2=0 $Y2=0
cc_33 N_B2_c_32_p N_9_c_125_n 4.28653e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_34 N_B2_c_35_p N_9_c_125_n 7.71172e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_35 N_B2_c_40_p N_9_c_125_n 0.00123965f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_36 N_B2_M2_g N_9_c_128_n 4.62717e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_37 VSS B2 0.00148665f $X=0.385 $Y=0.1335 $X2=0 $Y2=0
cc_38 VSS B2 0.00373029f $X=0.385 $Y=0.1335 $X2=0 $Y2=0
cc_39 VSS N_B2_c_40_p 5.36267e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_40 VSS N_B2_c_32_p 4.28653e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_41 VSS N_B2_c_40_p 5.36267e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_42 VSS N_B2_M2_g 2.21754e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_43 VSS N_B2_c_35_p 3.8028e-19 $X=0.459 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_44 VSS N_B2_c_35_p 8.0006e-19 $X=0.459 $Y=0.135 $X2=0.189 $Y2=0.135
cc_45 VSS N_B2_c_35_p 7.7076e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_46 VSS B2 3.72854e-19 $X=0.385 $Y=0.1335 $X2=0 $Y2=0
cc_47 VSS N_B2_M2_g 3.97719e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_48 N_B1_c_55_n N_9_c_129_n 8.0006e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_49 B1 N_9_c_129_n 0.00181344f $X=0.512 $Y=0.1415 $X2=0 $Y2=0
cc_50 N_B1_M3_g N_9_c_131_n 2.34993e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_51 B1 N_9_c_131_n 0.00397452f $X=0.512 $Y=0.1415 $X2=0 $Y2=0
cc_52 N_B1_c_55_n N_9_c_133_n 5.07795e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_53 N_B1_c_55_n N_9_c_134_n 4.62717e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_54 VSS B1 0.0313331f $X=0.512 $Y=0.1415 $X2=0 $Y2=0
cc_55 VSS N_B1_M3_g 2.38303e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_56 VSS N_B1_c_55_n 2.64781e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_57 VSS N_B1_c_55_n 3.80246e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_58 VSS N_B1_c_55_n 8.0006e-19 $X=0.567 $Y=0.135 $X2=0.459 $Y2=0.135
cc_59 VSS B1 3.21813e-19 $X=0.512 $Y=0.1415 $X2=0.459 $Y2=0.135
cc_60 VSS N_B1_M3_g 2.56447e-19 $X=0.513 $Y=0.0675 $X2=0.459 $Y2=0.135
cc_61 VSS B1 0.00376032f $X=0.512 $Y=0.1415 $X2=0.459 $Y2=0.135
cc_62 VSS N_B1_c_55_n 0.0012804f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_63 VSS B1 3.15243e-19 $X=0.512 $Y=0.1415 $X2=0.405 $Y2=0.135
cc_64 N_C1_c_74_p N_C2_M5_g 3.09654e-19 $X=0.729 $Y=0.135 $X2=0.513 $Y2=0.0675
cc_65 N_C1_M4_g N_C2_M5_g 0.00372052f $X=0.783 $Y=0.0675 $X2=0.513 $Y2=0.0675
cc_66 N_C1_M4_g N_C2_c_94_n 2.74891e-19 $X=0.783 $Y=0.0675 $X2=0.567 $Y2=0.135
cc_67 N_C1_c_77_p N_C2_c_94_n 0.00163635f $X=0.783 $Y=0.135 $X2=0.567 $Y2=0.135
cc_68 N_C1_c_77_p N_9_M17_d 3.80246e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_69 N_C1_c_77_p N_9_c_136_n 8.0006e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_70 N_C1_c_77_p N_9_c_137_n 8.0006e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_71 C1 N_9_c_137_n 0.00217241f $X=0.729 $Y=0.1405 $X2=0 $Y2=0
cc_72 N_C1_c_74_p N_9_c_139_n 2.38303e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_73 C1 N_9_c_139_n 0.00372924f $X=0.729 $Y=0.1405 $X2=0 $Y2=0
cc_74 N_C1_M4_g N_9_c_141_n 4.62717e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_75 N_C1_c_77_p N_9_c_141_n 5.14245e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_76 N_C1_M4_g N_9_c_143_n 2.64781e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_77 VSS C1 0.0314327f $X=0.729 $Y=0.1405 $X2=0 $Y2=0
cc_78 VSS N_C1_c_74_p 3.37536e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_79 VSS C1 0.00373921f $X=0.729 $Y=0.1405 $X2=0 $Y2=0
cc_80 VSS N_C1_c_77_p 8.7969e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_81 VSS N_C1_M4_g 3.97719e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_82 N_C2_c_94_n N_9_M19_d 3.80413e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_83 N_C2_c_94_n N_9_c_145_n 8.0006e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_84 N_C2_M5_g N_9_c_141_n 4.62717e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_85 N_C2_c_94_n N_9_c_141_n 7.70721e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_86 N_C2_c_94_n N_9_c_148_n 4.28653e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_87 C2 N_9_c_148_n 4.56869e-19 $X=0.904 $Y=0.1335 $X2=0 $Y2=0
cc_88 C2 N_9_c_150_n 0.00415841f $X=0.904 $Y=0.1335 $X2=0 $Y2=0
cc_89 N_C2_M5_g N_9_c_143_n 2.64781e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_90 N_C2_c_94_n N_9_c_143_n 2.64781e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_91 C2 N_9_c_143_n 3.33942e-19 $X=0.904 $Y=0.1335 $X2=0 $Y2=0
cc_92 C2 N_9_c_154_n 3.33942e-19 $X=0.904 $Y=0.1335 $X2=0 $Y2=0
cc_93 C2 N_9_c_155_n 0.00144692f $X=0.904 $Y=0.1335 $X2=0 $Y2=0
cc_94 C2 N_9_c_156_n 0.00144692f $X=0.904 $Y=0.1335 $X2=0 $Y2=0
cc_95 C2 N_9_c_157_n 0.00144692f $X=0.904 $Y=0.1335 $X2=0 $Y2=0
cc_96 VSS C2 0.00101254f $X=0.904 $Y=0.1335 $X2=0 $Y2=0
cc_97 VSS N_C2_M5_g 3.97719e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_98 VSS N_C2_c_94_n 8.66837e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_99 VSS N_C2_c_94_n 2.62734e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_100 VSS C2 0.00101254f $X=0.904 $Y=0.1335 $X2=0 $Y2=0
cc_101 VSS N_9_c_117_n 0.00104998f $X=0.108 $Y=0.036 $X2=0.081 $Y2=0.2025
cc_102 VSS N_9_c_115_n 4.62858e-19 $X=0.108 $Y=0.036 $X2=0 $Y2=0
cc_103 VSS N_9_c_119_n 2.31429e-19 $X=0.215 $Y=0.036 $X2=0 $Y2=0
cc_104 VSS N_9_c_161_p 2.31429e-19 $X=0.323 $Y=0.036 $X2=0 $Y2=0
cc_105 VSS N_9_c_125_n 2.31429e-19 $X=0.419 $Y=0.036 $X2=0 $Y2=0
cc_106 VSS N_9_c_128_n 2.31429e-19 $X=0.485 $Y=0.036 $X2=0 $Y2=0
cc_107 VSS N_9_c_143_n 2.93863e-19 $X=0.932 $Y=0.234 $X2=0 $Y2=0
cc_108 VSS N_9_c_129_n 0.00137166f $X=0.54 $Y=0.036 $X2=0.135 $Y2=0.135
cc_109 VSS N_9_c_136_n 0.00332785f $X=0.756 $Y=0.2025 $X2=0 $Y2=0
cc_110 VSS N_9_c_143_n 5.10653e-19 $X=0.932 $Y=0.234 $X2=0 $Y2=0
cc_111 VSS N_9_c_136_n 0.00361305f $X=0.756 $Y=0.2025 $X2=0 $Y2=0
cc_112 VSS N_9_c_145_n 0.00350515f $X=0.864 $Y=0.2025 $X2=0 $Y2=0
cc_113 VSS N_9_c_143_n 0.00250965f $X=0.932 $Y=0.234 $X2=0 $Y2=0
cc_114 VSS N_9_c_145_n 0.00350506f $X=0.864 $Y=0.2025 $X2=0.061 $Y2=0.135
cc_115 VSS N_9_c_143_n 0.00312698f $X=0.932 $Y=0.234 $X2=0.061 $Y2=0.135
cc_116 VSS N_9_c_173_p 4.08738e-19 $X=0.999 $Y=0.171 $X2=0.061 $Y2=0.135
cc_117 VSS N_9_c_125_n 5.33787e-19 $X=0.419 $Y=0.036 $X2=0 $Y2=0
cc_118 VSS N_9_c_128_n 5.33787e-19 $X=0.485 $Y=0.036 $X2=0 $Y2=0
cc_119 VSS N_9_c_133_n 5.33787e-19 $X=0.531 $Y=0.036 $X2=0 $Y2=0
cc_120 VSS N_9_c_134_n 5.33787e-19 $X=0.701 $Y=0.036 $X2=0.135 $Y2=0.135
cc_121 VSS N_9_c_141_n 5.33787e-19 $X=0.877 $Y=0.036 $X2=0 $Y2=0
cc_122 VSS N_9_c_148_n 5.33787e-19 $X=0.917 $Y=0.036 $X2=0 $Y2=0
cc_123 VSS N_9_c_180_p 6.06775e-19 $X=0.999 $Y=0.207 $X2=0 $Y2=0
cc_124 VSS N_9_c_136_n 0.00233206f $X=0.756 $Y=0.2025 $X2=0 $Y2=0
cc_125 VSS N_9_c_145_n 0.00233206f $X=0.864 $Y=0.2025 $X2=0 $Y2=0
cc_126 VSS N_9_c_143_n 0.0155792f $X=0.932 $Y=0.234 $X2=0 $Y2=0
cc_127 N_9_c_184_p N_Y_M7_d 3.80529e-19 $X=1.107 $Y=0.135 $X2=0.081 $Y2=0.135
cc_128 N_9_c_184_p N_Y_M21_d 3.80529e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_129 N_9_c_184_p N_Y_c_201_n 8.00061e-19 $X=1.107 $Y=0.135 $X2=0.135 $Y2=0.135
cc_130 N_9_M7_g N_Y_c_202_n 4.59284e-19 $X=1.107 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_131 N_9_c_184_p N_Y_c_202_n 5.51214e-19 $X=1.107 $Y=0.135 $X2=0.135 $Y2=0.135
cc_132 N_9_c_189_p N_Y_c_202_n 4.03778e-19 $X=0.99 $Y=0.036 $X2=0.135 $Y2=0.135
cc_133 N_9_c_184_p N_Y_c_205_n 8.00061e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_134 N_9_M7_g N_Y_c_206_n 4.59284e-19 $X=1.107 $Y=0.0675 $X2=0 $Y2=0
cc_135 N_9_c_184_p N_Y_c_206_n 5.51214e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_136 N_9_c_193_p N_Y_c_206_n 4.00248e-19 $X=0.99 $Y=0.234 $X2=0 $Y2=0
cc_137 N_9_c_184_p N_Y_c_209_n 4.96657e-19 $X=1.107 $Y=0.135 $X2=0.061
+ $Y2=0.1335
cc_138 N_9_c_156_n N_Y_c_209_n 3.19589e-19 $X=0.999 $Y=0.0945 $X2=0.061
+ $Y2=0.1335
cc_139 N_9_c_196_p N_Y_c_211_n 2.25338e-19 $X=1.052 $Y=0.135 $X2=0 $Y2=0
cc_140 VSS N_9_c_119_n 4.62297e-19 $X=0.215 $Y=0.036 $X2=0.081 $Y2=0.135
cc_141 VSS N_9_c_141_n 4.54171e-19 $X=0.877 $Y=0.036 $X2=0.081 $Y2=0.135

* END of "./AO222x2_ASAP7_75t_L.pex.sp.AO222X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO22x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:04:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO22x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO22x1_ASAP7_75t_L.pex.sp.pex"
* File: AO22x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:04:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO22X1_ASAP7_75T_L%A1 2 5 7 16 19 21 22 26 VSS
c14 26 VSS 0.0124301f $X=0.018 $Y=0.135
c15 22 VSS 7.38238e-19 $X=0.0635 $Y=0.135
c16 21 VSS 8.96246e-19 $X=0.046 $Y=0.135
c17 19 VSS 9.39933e-19 $X=0.081 $Y=0.135
c18 16 VSS 0.00531417f $X=0.018 $Y=0.151
c19 5 VSS 0.00274291f $X=0.081 $Y=0.135
c20 2 VSS 0.0645488f $X=0.081 $Y=0.054
r21 21 22 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r22 19 22 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r23 17 26 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r24 17 21 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.046 $Y2=0.135
r25 13 26 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r26 13 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.151
r27 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r28 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r29 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO22X1_ASAP7_75T_L%A2 2 5 7 12 17 19 VSS
c17 19 VSS 1.81759e-19 $X=0.135 $Y=0.164
c18 17 VSS 0.00314757f $X=0.134 $Y=0.186
c19 12 VSS 0.00147988f $X=0.135 $Y=0.135
c20 5 VSS 0.00116811f $X=0.135 $Y=0.135
c21 2 VSS 0.0602966f $X=0.135 $Y=0.054
r22 18 19 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.164
r23 17 19 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.186 $X2=0.135 $Y2=0.164
r24 12 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r25 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r26 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r27 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO22X1_ASAP7_75T_L%B2 2 5 7 10 VSS
c12 10 VSS 6.22747e-19 $X=0.188 $Y=0.115
c13 5 VSS 0.00110682f $X=0.189 $Y=0.135
c14 2 VSS 0.0604449f $X=0.189 $Y=0.054
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO22X1_ASAP7_75T_L%B1 2 5 7 11 13 VSS
c12 13 VSS 5.17197e-19 $X=0.243 $Y=0.135
c13 11 VSS 0.00374061f $X=0.243 $Y=0.081
c14 5 VSS 0.00210567f $X=0.243 $Y=0.135
c15 2 VSS 0.0631344f $X=0.243 $Y=0.054
r16 11 13 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r19 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO22X1_ASAP7_75T_L%7 2 5 7 9 10 13 14 15 18 19 21 27 30 37 38 39 42
+ 43 44 47 51 VSS
c29 55 VSS 4.18034e-19 $X=0.351 $Y=0.135
c30 51 VSS 0.00340617f $X=0.405 $Y=0.135
c31 48 VSS 5.18771e-19 $X=0.351 $Y=0.1765
c32 47 VSS 6.20958e-19 $X=0.351 $Y=0.164
c33 46 VSS 3.04011e-19 $X=0.351 $Y=0.189
c34 44 VSS 9.74222e-19 $X=0.351 $Y=0.081
c35 43 VSS 9.5529e-19 $X=0.351 $Y=0.063
c36 42 VSS 0.00159541f $X=0.351 $Y=0.126
c37 40 VSS 2.02755e-19 $X=0.287 $Y=0.198
c38 39 VSS 4.31692e-19 $X=0.284 $Y=0.198
c39 38 VSS 8.46035e-21 $X=0.252 $Y=0.198
c40 37 VSS 5.02599e-19 $X=0.234 $Y=0.198
c41 32 VSS 0.00627269f $X=0.342 $Y=0.198
c42 31 VSS 0.0035163f $X=0.3145 $Y=0.036
c43 30 VSS 0.00748237f $X=0.287 $Y=0.036
c44 29 VSS 0.00311169f $X=0.234 $Y=0.036
c45 28 VSS 4.32241e-19 $X=0.202 $Y=0.036
c46 27 VSS 0.00146362f $X=0.198 $Y=0.036
c47 26 VSS 0.00269651f $X=0.18 $Y=0.036
c48 21 VSS 0.00479518f $X=0.162 $Y=0.036
c49 19 VSS 0.00652675f $X=0.342 $Y=0.036
c50 18 VSS 0.00219578f $X=0.216 $Y=0.216
c51 14 VSS 5.7036e-19 $X=0.233 $Y=0.216
c52 13 VSS 0.00428109f $X=0.162 $Y=0.054
c53 9 VSS 5.3314e-19 $X=0.179 $Y=0.054
c54 5 VSS 0.00384735f $X=0.405 $Y=0.135
c55 2 VSS 0.067966f $X=0.405 $Y=0.0675
r56 49 55 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.135 $X2=0.351 $Y2=0.135
r57 49 51 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.135 $X2=0.405 $Y2=0.135
r58 47 48 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.164 $X2=0.351 $Y2=0.1765
r59 46 48 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.1765
r60 45 55 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.144 $X2=0.351 $Y2=0.135
r61 45 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.144 $X2=0.351 $Y2=0.164
r62 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.063 $X2=0.351 $Y2=0.081
r63 42 55 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.135
r64 42 44 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.081
r65 41 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.063
r66 39 40 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.198 $X2=0.287 $Y2=0.198
r67 38 39 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.284 $Y2=0.198
r68 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.252 $Y2=0.198
r69 34 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.234 $Y2=0.198
r70 32 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.198 $X2=0.351 $Y2=0.189
r71 32 40 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.287 $Y2=0.198
r72 30 31 1.86728 $w=1.8e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.287
+ $Y=0.036 $X2=0.3145 $Y2=0.036
r73 29 30 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.287 $Y2=0.036
r74 28 29 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.036 $X2=0.234 $Y2=0.036
r75 27 28 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.202 $Y2=0.036
r76 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r77 21 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r78 19 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.036 $X2=0.351 $Y2=0.045
r79 19 31 1.86728 $w=1.8e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.3145 $Y2=0.036
r80 18 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r81 15 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.216 $X2=0.216 $Y2=0.216
r82 14 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.216 $X2=0.216 $Y2=0.216
r83 13 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r84 10 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.162 $Y2=0.054
r85 9 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.054 $X2=0.162 $Y2=0.054
r86 5 51 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r87 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r88 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO22X1_ASAP7_75T_L%Y 1 6 14 15 16 18 20 30 VSS
c6 36 VSS 0.00267977f $X=0.45 $Y=0.234
c7 35 VSS 0.00278493f $X=0.459 $Y=0.234
c8 30 VSS 0.00161219f $X=0.432 $Y=0.234
c9 26 VSS 0.00267977f $X=0.45 $Y=0.036
c10 25 VSS 0.00278493f $X=0.459 $Y=0.036
c11 21 VSS 0.00641078f $X=0.432 $Y=0.036
c12 20 VSS 0.00141731f $X=0.432 $Y=0.036
c13 18 VSS 0.00286206f $X=0.459 $Y=0.207
c14 16 VSS 2.52491e-19 $X=0.459 $Y=0.132
c15 15 VSS 0.00391028f $X=0.459 $Y=0.126
c16 14 VSS 4.87872e-19 $X=0.459 $Y=0.138
c17 12 VSS 0.00102822f $X=0.459 $Y=0.225
c18 9 VSS 0.00675415f $X=0.43 $Y=0.2025
c19 4 VSS 3.41873e-19 $X=0.43 $Y=0.0675
r20 36 37 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.4545 $Y2=0.234
r21 35 37 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.234 $X2=0.4545 $Y2=0.234
r22 30 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.45 $Y2=0.234
r23 26 27 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r24 25 27 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r25 20 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r26 20 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r27 17 18 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.144 $X2=0.459 $Y2=0.207
r28 15 16 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.126 $X2=0.459 $Y2=0.132
r29 14 17 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.138 $X2=0.459 $Y2=0.144
r30 14 16 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.138 $X2=0.459 $Y2=0.132
r31 12 35 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.234
r32 12 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.207
r33 11 25 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r34 11 15 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.126
r35 9 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r36 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2025 $X2=0.43 $Y2=0.2025
r37 4 21 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r38 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.43 $Y2=0.0675
.ends


* END of "./AO22x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO22x1_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 Y
* 
* Y	Y
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 noxref_10 N_A1_M0_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_7_M1_d N_A2_M1_g noxref_10 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 noxref_11 N_B2_M2_g N_7_M2_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.027
M3 VSS N_B1_M3_g noxref_11 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_7_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M5 VDD N_A1_M5_g noxref_8 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M6 noxref_8 N_A2_M6_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M7 N_7_M7_d N_B2_M7_g noxref_8 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M8 noxref_8 N_B1_M8_g N_7_M8_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M9 N_Y_M9_d N_7_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.162
*
* 
* .include "AO22x1_ASAP7_75t_L.pex.sp.AO22X1_ASAP7_75T_L.pxi"
* BEGIN of "./AO22x1_ASAP7_75t_L.pex.sp.AO22X1_ASAP7_75T_L.pxi"
* File: AO22x1_ASAP7_75t_L.pex.sp.AO22X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:04:41 2017
* 
x_PM_AO22X1_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M5_g A1 N_A1_c_3_p
+ N_A1_c_11_p N_A1_c_12_p N_A1_c_4_p VSS PM_AO22X1_ASAP7_75T_L%A1
x_PM_AO22X1_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_16_n N_A2_M6_g N_A2_c_17_n A2
+ N_A2_c_20_n VSS PM_AO22X1_ASAP7_75T_L%A2
x_PM_AO22X1_ASAP7_75T_L%B2 N_B2_M2_g N_B2_c_34_n N_B2_M7_g B2 VSS
+ PM_AO22X1_ASAP7_75T_L%B2
x_PM_AO22X1_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_46_n N_B1_M8_g B1 N_B1_c_51_p VSS
+ PM_AO22X1_ASAP7_75T_L%B1
x_PM_AO22X1_ASAP7_75T_L%7 N_7_M4_g N_7_c_80_p N_7_M9_g N_7_M2_s N_7_M1_d
+ N_7_c_57_n N_7_M8_s N_7_M7_d N_7_c_72_p N_7_c_83_p N_7_c_56_n N_7_c_62_n
+ N_7_c_64_n N_7_c_60_n N_7_c_66_n N_7_c_68_n N_7_c_69_n N_7_c_79_p N_7_c_70_n
+ N_7_c_82_p N_7_c_81_p VSS PM_AO22X1_ASAP7_75T_L%7
x_PM_AO22X1_ASAP7_75T_L%Y N_Y_M4_d N_Y_M9_d Y N_Y_c_85_n N_Y_c_86_n N_Y_c_88_n
+ N_Y_c_89_n N_Y_c_90_n VSS PM_AO22X1_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00315405f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A1_c_2_p N_A2_c_16_n 0.00120928f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p N_A2_c_17_n 8.78098e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A1_c_4_p N_A2_c_17_n 0.00104667f $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.135
cc_5 A1 A2 3.12618e-19 $X=0.018 $Y=0.151 $X2=0.134 $Y2=0.186
cc_6 A1 N_A2_c_20_n 8.11421e-19 $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.164
cc_7 N_A1_M0_g N_B2_M2_g 2.60137e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_8 N_A1_c_4_p N_7_c_56_n 4.58091e-19 $X=0.018 $Y=0.135 $X2=0 $Y2=0
cc_9 VSS A1 0.00131018f $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.135
cc_10 VSS A1 7.45437e-19 $X=0.018 $Y=0.151 $X2=0.134 $Y2=0.186
cc_11 VSS N_A1_c_11_p 3.14847e-19 $X=0.046 $Y=0.135 $X2=0.134 $Y2=0.186
cc_12 VSS N_A1_c_12_p 3.14847e-19 $X=0.0635 $Y=0.135 $X2=0.134 $Y2=0.186
cc_13 VSS N_A1_M0_g 4.28653e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_14 VSS N_A1_c_3_p 3.14847e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_15 N_A2_M1_g N_B2_M2_g 0.00353901f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_16 N_A2_c_16_n N_B2_c_34_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_17 N_A2_c_17_n B2 0.00436278f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_18 N_A2_M1_g N_B1_M3_g 2.949e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_19 N_A2_c_17_n N_7_c_57_n 6.66766e-19 $X=0.135 $Y=0.135 $X2=0.018 $Y2=0.144
cc_20 N_A2_M1_g N_7_c_56_n 2.34993e-19 $X=0.135 $Y=0.054 $X2=0.046 $Y2=0.135
cc_21 N_A2_c_17_n N_7_c_56_n 0.00399258f $X=0.135 $Y=0.135 $X2=0.046 $Y2=0.135
cc_22 A2 N_7_c_60_n 4.29446e-19 $X=0.134 $Y=0.186 $X2=0 $Y2=0
cc_23 VSS A2 6.13941e-19 $X=0.134 $Y=0.186 $X2=0 $Y2=0
cc_24 VSS N_A2_M1_g 2.34993e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_25 VSS A2 0.00375082f $X=0.134 $Y=0.186 $X2=0 $Y2=0
cc_26 N_B2_M2_g N_B1_M3_g 0.00358983f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_27 N_B2_c_34_n N_B1_c_46_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_28 B2 B1 0.00480954f $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_29 B2 N_7_c_57_n 3.87865e-19 $X=0.188 $Y=0.115 $X2=0.018 $Y2=0.144
cc_30 N_B2_M2_g N_7_c_62_n 2.64276e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_31 B2 N_7_c_62_n 0.00124805f $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_32 VSS N_B2_M2_g 3.57119e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_33 VSS B2 5.37372e-19 $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_34 N_B1_M3_g N_7_c_64_n 2.34993e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_35 B1 N_7_c_64_n 0.00497576f $X=0.243 $Y=0.081 $X2=0 $Y2=0
cc_36 N_B1_M3_g N_7_c_66_n 2.76185e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_37 N_B1_c_51_p N_7_c_66_n 0.00123353f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_38 B1 N_7_c_68_n 3.92634e-19 $X=0.243 $Y=0.081 $X2=0 $Y2=0
cc_39 N_B1_c_51_p N_7_c_69_n 0.00143736f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_40 B1 N_7_c_70_n 5.57293e-19 $X=0.243 $Y=0.081 $X2=0 $Y2=0
cc_41 VSS N_B1_M3_g 2.08515e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_42 VSS N_7_c_57_n 6.80422e-19 $X=0.162 $Y=0.054 $X2=0 $Y2=0
cc_43 VSS N_7_c_72_p 0.00288888f $X=0.216 $Y=0.216 $X2=0 $Y2=0
cc_44 VSS N_7_c_60_n 3.94585e-19 $X=0.234 $Y=0.198 $X2=0 $Y2=0
cc_45 VSS N_7_c_72_p 0.00302498f $X=0.216 $Y=0.216 $X2=0 $Y2=0
cc_46 VSS N_7_c_68_n 0.00397265f $X=0.284 $Y=0.198 $X2=0 $Y2=0
cc_47 VSS N_7_c_66_n 0.00352873f $X=0.252 $Y=0.198 $X2=0 $Y2=0
cc_48 VSS N_7_c_72_p 0.00250965f $X=0.216 $Y=0.216 $X2=0 $Y2=0
cc_49 VSS N_7_c_60_n 0.00352873f $X=0.234 $Y=0.198 $X2=0 $Y2=0
cc_50 N_7_c_79_p N_Y_c_85_n 7.67125e-19 $X=0.351 $Y=0.063 $X2=0.018 $Y2=0.151
cc_51 N_7_c_80_p N_Y_c_86_n 3.14724e-19 $X=0.405 $Y=0.135 $X2=0.018 $Y2=0.151
cc_52 N_7_c_81_p N_Y_c_86_n 0.00101388f $X=0.405 $Y=0.135 $X2=0.018 $Y2=0.151
cc_53 N_7_c_82_p N_Y_c_88_n 6.45145e-19 $X=0.351 $Y=0.164 $X2=0.081 $Y2=0.135
cc_54 N_7_c_83_p N_Y_c_89_n 3.79692e-19 $X=0.342 $Y=0.036 $X2=0.081 $Y2=0.135
cc_55 VSS N_7_c_56_n 2.90855e-19 $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.054
cc_56 VSS N_Y_c_90_n 2.40402e-19 $X=0.27 $Y=0.234 $X2=0 $Y2=0

* END of "./AO22x1_ASAP7_75t_L.pex.sp.AO22X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO22x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:05:04 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO22x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO22x2_ASAP7_75t_L.pex.sp.pex"
* File: AO22x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:05:04 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO22X2_ASAP7_75T_L%A1 2 5 7 16 19 21 22 26 VSS
c14 26 VSS 0.0122468f $X=0.018 $Y=0.135
c15 22 VSS 6.65175e-19 $X=0.0635 $Y=0.135
c16 21 VSS 0.00101906f $X=0.046 $Y=0.135
c17 19 VSS 0.00105225f $X=0.081 $Y=0.135
c18 16 VSS 0.00492582f $X=0.018 $Y=0.151
c19 5 VSS 0.00274291f $X=0.081 $Y=0.135
c20 2 VSS 0.0645488f $X=0.081 $Y=0.0675
r21 21 22 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r22 19 22 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r23 17 26 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r24 17 21 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.046 $Y2=0.135
r25 13 26 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r26 13 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.151
r27 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r28 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r29 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO22X2_ASAP7_75T_L%A2 2 5 7 12 17 19 VSS
c17 19 VSS 2.43609e-19 $X=0.135 $Y=0.164
c18 17 VSS 0.0027918f $X=0.134 $Y=0.186
c19 12 VSS 0.00183316f $X=0.135 $Y=0.135
c20 5 VSS 0.00116811f $X=0.135 $Y=0.135
c21 2 VSS 0.0602966f $X=0.135 $Y=0.0675
r22 18 19 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.164
r23 17 19 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.186 $X2=0.135 $Y2=0.164
r24 12 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r25 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO22X2_ASAP7_75T_L%B2 2 5 7 10 VSS
c12 10 VSS 5.22847e-19 $X=0.188 $Y=0.115
c13 5 VSS 0.00110682f $X=0.189 $Y=0.135
c14 2 VSS 0.0604449f $X=0.189 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO22X2_ASAP7_75T_L%B1 2 5 7 11 13 VSS
c12 13 VSS 0.00162001f $X=0.243 $Y=0.135
c13 11 VSS 0.00258486f $X=0.243 $Y=0.081
c14 5 VSS 0.00210567f $X=0.243 $Y=0.135
c15 2 VSS 0.0631344f $X=0.243 $Y=0.0675
r16 11 13 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO22X2_ASAP7_75T_L%7 2 7 10 13 15 17 18 22 23 26 27 29 30 35 37 38 45
+ 46 47 50 52 55 59 VSS
c38 63 VSS 4.18034e-19 $X=0.351 $Y=0.135
c39 59 VSS 0.00322784f $X=0.405 $Y=0.135
c40 56 VSS 7.76721e-19 $X=0.351 $Y=0.1765
c41 55 VSS 9.50916e-19 $X=0.351 $Y=0.164
c42 54 VSS 7.17985e-19 $X=0.351 $Y=0.189
c43 52 VSS 0.00113859f $X=0.351 $Y=0.081
c44 51 VSS 0.00109324f $X=0.351 $Y=0.063
c45 50 VSS 0.00278428f $X=0.351 $Y=0.126
c46 48 VSS 2.02755e-19 $X=0.287 $Y=0.198
c47 47 VSS 4.4302e-19 $X=0.284 $Y=0.198
c48 46 VSS 8.46035e-21 $X=0.252 $Y=0.198
c49 45 VSS 4.59335e-19 $X=0.234 $Y=0.198
c50 40 VSS 0.00636518f $X=0.342 $Y=0.198
c51 39 VSS 0.0035163f $X=0.3145 $Y=0.036
c52 38 VSS 0.00753002f $X=0.287 $Y=0.036
c53 37 VSS 0.00291823f $X=0.234 $Y=0.036
c54 36 VSS 4.1976e-19 $X=0.202 $Y=0.036
c55 35 VSS 0.00146362f $X=0.198 $Y=0.036
c56 34 VSS 0.00264888f $X=0.18 $Y=0.036
c57 30 VSS 0.00503645f $X=0.162 $Y=0.036
c58 29 VSS 0.00474537f $X=0.162 $Y=0.036
c59 27 VSS 0.00652675f $X=0.342 $Y=0.036
c60 26 VSS 0.00243084f $X=0.216 $Y=0.2025
c61 22 VSS 5.75997e-19 $X=0.233 $Y=0.2025
c62 17 VSS 5.38922e-19 $X=0.179 $Y=0.0675
c63 13 VSS 0.00546085f $X=0.459 $Y=0.135
c64 10 VSS 0.0634956f $X=0.459 $Y=0.0675
c65 2 VSS 0.0640381f $X=0.405 $Y=0.0675
r66 57 63 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.135 $X2=0.351 $Y2=0.135
r67 57 59 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.135 $X2=0.405 $Y2=0.135
r68 55 56 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.164 $X2=0.351 $Y2=0.1765
r69 54 56 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.1765
r70 53 63 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.144 $X2=0.351 $Y2=0.135
r71 53 55 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.144 $X2=0.351 $Y2=0.164
r72 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.063 $X2=0.351 $Y2=0.081
r73 50 63 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.135
r74 50 52 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.081
r75 49 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.063
r76 47 48 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.198 $X2=0.287 $Y2=0.198
r77 46 47 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.284 $Y2=0.198
r78 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.252 $Y2=0.198
r79 42 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.234 $Y2=0.198
r80 40 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.198 $X2=0.351 $Y2=0.189
r81 40 48 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.287 $Y2=0.198
r82 38 39 1.86728 $w=1.8e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.287
+ $Y=0.036 $X2=0.3145 $Y2=0.036
r83 37 38 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.287 $Y2=0.036
r84 36 37 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.036 $X2=0.234 $Y2=0.036
r85 35 36 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.202 $Y2=0.036
r86 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r87 29 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r88 29 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r89 27 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.036 $X2=0.351 $Y2=0.045
r90 27 39 1.86728 $w=1.8e-08 $l=2.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.3145 $Y2=0.036
r91 26 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r92 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r93 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r94 21 30 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r95 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r96 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r97 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r98 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r99 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r100 5 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r101 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r102 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO22X2_ASAP7_75T_L%Y 1 2 6 7 10 11 13 14 18 20 28 29 30 32 VSS
c14 32 VSS 0.00379776f $X=0.513 $Y=0.207
c15 30 VSS 2.69413e-19 $X=0.513 $Y=0.132
c16 29 VSS 0.00468461f $X=0.513 $Y=0.126
c17 28 VSS 5.05149e-19 $X=0.513 $Y=0.138
c18 26 VSS 8.85605e-19 $X=0.513 $Y=0.225
c19 20 VSS 0.00158432f $X=0.432 $Y=0.234
c20 18 VSS 0.0130697f $X=0.504 $Y=0.234
c21 14 VSS 0.00904188f $X=0.432 $Y=0.036
c22 13 VSS 0.00138529f $X=0.432 $Y=0.036
c23 11 VSS 0.0130697f $X=0.504 $Y=0.036
c24 10 VSS 0.00904877f $X=0.432 $Y=0.2025
c25 6 VSS 5.58795e-19 $X=0.449 $Y=0.2025
c26 1 VSS 5.58795e-19 $X=0.449 $Y=0.0675
r27 31 32 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.144 $X2=0.513 $Y2=0.207
r28 29 30 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.126 $X2=0.513 $Y2=0.132
r29 28 31 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.138 $X2=0.513 $Y2=0.144
r30 28 30 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.138 $X2=0.513 $Y2=0.132
r31 26 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.207
r32 25 29 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.126
r33 18 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.234 $X2=0.513 $Y2=0.225
r34 18 20 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.432 $Y2=0.234
r35 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r36 11 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.036 $X2=0.513 $Y2=0.045
r37 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.432 $Y2=0.036
r38 10 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r39 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r40 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r41 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r42 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.432 $Y2=0.0675
r43 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.449
+ $Y=0.0675 $X2=0.432 $Y2=0.0675
.ends


* END of "./AO22x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO22x2_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 Y
* 
* Y	Y
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 noxref_10 N_A1_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_7_M1_d N_A2_M1_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_11 N_B2_M2_g N_7_M2_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_B1_M3_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_7_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M5 N_Y_M5_d N_7_M5_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M6 VDD N_A1_M6_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 noxref_8 N_A2_M7_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 N_7_M8_d N_B2_M8_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 noxref_8 N_B1_M9_g N_7_M9_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 N_Y_M10_d N_7_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M11 N_Y_M11_d N_7_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "AO22x2_ASAP7_75t_L.pex.sp.AO22X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO22x2_ASAP7_75t_L.pex.sp.AO22X2_ASAP7_75T_L.pxi"
* File: AO22x2_ASAP7_75t_L.pex.sp.AO22X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:05:04 2017
* 
x_PM_AO22X2_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M6_g A1 N_A1_c_3_p
+ N_A1_c_11_p N_A1_c_12_p N_A1_c_4_p VSS PM_AO22X2_ASAP7_75T_L%A1
x_PM_AO22X2_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_16_n N_A2_M7_g N_A2_c_17_n A2
+ N_A2_c_20_n VSS PM_AO22X2_ASAP7_75T_L%A2
x_PM_AO22X2_ASAP7_75T_L%B2 N_B2_M2_g N_B2_c_34_n N_B2_M8_g B2 VSS
+ PM_AO22X2_ASAP7_75T_L%B2
x_PM_AO22X2_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_46_n N_B1_M9_g B1 N_B1_c_51_p VSS
+ PM_AO22X2_ASAP7_75T_L%B1
x_PM_AO22X2_ASAP7_75T_L%7 N_7_M4_g N_7_M10_g N_7_M5_g N_7_c_79_p N_7_M11_g
+ N_7_M2_s N_7_M1_d N_7_M9_s N_7_M8_d N_7_c_71_p N_7_c_84_p N_7_c_56_n
+ N_7_c_59_n N_7_c_62_n N_7_c_93_p N_7_c_64_n N_7_c_60_n N_7_c_66_n N_7_c_68_n
+ N_7_c_69_n N_7_c_70_n N_7_c_91_p N_7_c_90_p VSS PM_AO22X2_ASAP7_75T_L%7
x_PM_AO22X2_ASAP7_75T_L%Y N_Y_M5_d N_Y_M4_d N_Y_M11_d N_Y_M10_d N_Y_c_96_n
+ N_Y_c_97_n N_Y_c_98_n N_Y_c_100_n N_Y_c_101_n N_Y_c_102_n Y N_Y_c_103_n
+ N_Y_c_105_n N_Y_c_106_n VSS PM_AO22X2_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00315405f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_16_n 0.00120928f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p N_A2_c_17_n 8.78098e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A1_c_4_p N_A2_c_17_n 7.94587e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.135
cc_5 A1 A2 3.12618e-19 $X=0.018 $Y=0.151 $X2=0.134 $Y2=0.186
cc_6 A1 N_A2_c_20_n 4.69126e-19 $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.164
cc_7 N_A1_M0_g N_B2_M2_g 2.60137e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_8 N_A1_c_4_p N_7_c_56_n 4.58091e-19 $X=0.018 $Y=0.135 $X2=0 $Y2=0
cc_9 VSS A1 0.00201602f $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.135
cc_10 VSS A1 7.45434e-19 $X=0.018 $Y=0.151 $X2=0.134 $Y2=0.186
cc_11 VSS N_A1_c_11_p 3.04973e-19 $X=0.046 $Y=0.135 $X2=0.134 $Y2=0.186
cc_12 VSS N_A1_c_12_p 3.04973e-19 $X=0.0635 $Y=0.135 $X2=0.134 $Y2=0.186
cc_13 VSS N_A1_M0_g 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_14 VSS N_A1_c_3_p 3.04973e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_15 N_A2_M1_g N_B2_M2_g 0.00353901f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_A2_c_16_n N_B2_c_34_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_17 N_A2_c_17_n B2 0.00382022f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_18 N_A2_M1_g N_B1_M3_g 2.949e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_19 N_A2_M1_g N_7_c_56_n 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_20 N_A2_c_17_n N_7_c_56_n 0.00399257f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_21 N_A2_c_17_n N_7_c_59_n 0.00160911f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_22 A2 N_7_c_60_n 4.29446e-19 $X=0.134 $Y=0.186 $X2=0 $Y2=0
cc_23 VSS N_A2_c_20_n 0.00123948f $X=0.135 $Y=0.164 $X2=0 $Y2=0
cc_24 VSS N_A2_M1_g 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_25 VSS A2 0.00375082f $X=0.134 $Y=0.186 $X2=0 $Y2=0
cc_26 N_B2_M2_g N_B1_M3_g 0.00358983f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_27 N_B2_c_34_n N_B1_c_46_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_28 B2 B1 0.00468225f $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_29 B2 N_7_c_59_n 0.0013399f $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_30 N_B2_M2_g N_7_c_62_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_31 B2 N_7_c_62_n 0.00124805f $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_32 VSS N_B2_M2_g 3.57119e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_33 VSS B2 5.37372e-19 $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_34 N_B1_M3_g N_7_c_64_n 2.34993e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_35 B1 N_7_c_64_n 0.00497575f $X=0.243 $Y=0.081 $X2=0 $Y2=0
cc_36 N_B1_M3_g N_7_c_66_n 2.76185e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_B1_c_51_p N_7_c_66_n 0.00123353f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_38 B1 N_7_c_68_n 3.60257e-19 $X=0.243 $Y=0.081 $X2=0 $Y2=0
cc_39 N_B1_c_51_p N_7_c_69_n 0.00117553f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_40 B1 N_7_c_70_n 5.57293e-19 $X=0.243 $Y=0.081 $X2=0 $Y2=0
cc_41 VSS N_B1_M3_g 2.08515e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_42 VSS N_7_c_71_p 0.00369767f $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_43 VSS N_7_c_59_n 0.00107252f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_44 VSS N_7_c_60_n 3.94585e-19 $X=0.234 $Y=0.198 $X2=0 $Y2=0
cc_45 VSS N_7_c_71_p 0.00360077f $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_46 VSS N_7_c_68_n 0.00288786f $X=0.284 $Y=0.198 $X2=0 $Y2=0
cc_47 VSS N_7_c_66_n 0.00352872f $X=0.252 $Y=0.198 $X2=0 $Y2=0
cc_48 VSS N_7_c_71_p 0.00250965f $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_49 VSS N_7_c_60_n 0.00352872f $X=0.234 $Y=0.198 $X2=0 $Y2=0
cc_50 N_7_c_79_p N_Y_M5_d 3.80485e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_51 N_7_c_79_p N_Y_M11_d 3.80485e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_52 N_7_c_79_p N_Y_c_96_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_53 N_7_M5_g N_Y_c_97_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_54 N_7_c_79_p N_Y_c_98_n 5.20568e-19 $X=0.459 $Y=0.135 $X2=0.018 $Y2=0.144
cc_55 N_7_c_84_p N_Y_c_98_n 4.00023e-19 $X=0.342 $Y=0.036 $X2=0.018 $Y2=0.144
cc_56 N_7_c_79_p N_Y_c_100_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_57 N_7_M5_g N_Y_c_101_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_58 N_7_c_79_p N_Y_c_102_n 5.20568e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.135
cc_59 N_7_c_79_p N_Y_c_103_n 4.85747e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_60 N_7_c_70_n N_Y_c_103_n 3.19725e-19 $X=0.351 $Y=0.081 $X2=0 $Y2=0
cc_61 N_7_c_90_p N_Y_c_105_n 2.31129e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_62 N_7_c_91_p N_Y_c_106_n 3.22582e-19 $X=0.351 $Y=0.164 $X2=0 $Y2=0
cc_63 VSS N_7_c_56_n 2.82273e-19 $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_64 VSS N_7_c_93_p 3.19955e-19 $X=0.234 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_65 VSS N_Y_c_102_n 2.68802e-19 $X=0.27 $Y=0.234 $X2=0.081 $Y2=0.135

* END of "./AO22x2_ASAP7_75t_L.pex.sp.AO22X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO31x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:05:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO31x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO31x2_ASAP7_75t_L.pex.sp.pex"
* File: AO31x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:05:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO31X2_ASAP7_75T_L%A3 2 7 10 13 15 25 VSS
c18 25 VSS 0.0201929f $X=0.08 $Y=0.136
c19 13 VSS 0.00774036f $X=0.135 $Y=0.135
c20 10 VSS 0.0630502f $X=0.135 $Y=0.0675
c21 2 VSS 0.0670913f $X=0.081 $Y=0.0675
r22 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r23 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r24 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r25 5 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO31X2_ASAP7_75T_L%B 2 7 10 13 21 VSS
c30 21 VSS 0.00683156f $X=0.189 $Y=0.134
c31 10 VSS 0.0724175f $X=0.243 $Y=0.135
c32 2 VSS 0.0625257f $X=0.189 $Y=0.054
r33 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r34 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r35 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r36 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r37 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO31X2_ASAP7_75T_L%A2 2 7 10 13 15 34 VSS
c33 34 VSS 0.00550204f $X=0.403 $Y=0.137
c34 13 VSS 0.00374929f $X=0.459 $Y=0.135
c35 10 VSS 0.0631881f $X=0.459 $Y=0.0675
c36 2 VSS 0.0663501f $X=0.405 $Y=0.0675
r37 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r38 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r39 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r40 5 34 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r41 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r42 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO31X2_ASAP7_75T_L%A1 2 7 10 13 15 32 VSS
c29 32 VSS 0.00265998f $X=0.569 $Y=0.137
c30 13 VSS 0.00407881f $X=0.567 $Y=0.135
c31 10 VSS 0.0659479f $X=0.567 $Y=0.0675
c32 2 VSS 0.0628224f $X=0.513 $Y=0.0675
r33 13 32 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r34 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r35 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r36 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r37 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r38 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AO31X2_ASAP7_75T_L%7 2 7 10 13 15 17 20 22 23 27 28 31 34 35 36 40 41
+ 42 43 44 45 46 48 49 50 53 55 59 60 62 63 64 65 66 75 81 90 95 99 VSS
c76 99 VSS 4.33032e-19 $X=0.675 $Y=0.135
c77 96 VSS 2.67452e-19 $X=0.234 $Y=0.072
c78 95 VSS 3.64491e-19 $X=0.243 $Y=0.072
c79 90 VSS 5.88777e-19 $X=0.216 $Y=0.072
c80 87 VSS 1.77025e-19 $X=0.234 $Y=0.198
c81 81 VSS 3.58568e-19 $X=0.216 $Y=0.198
c82 75 VSS 0.00340212f $X=0.729 $Y=0.135
c83 72 VSS 0.00108998f $X=0.675 $Y=0.207
c84 71 VSS 0.00165812f $X=0.675 $Y=0.189
c85 70 VSS 0.00147802f $X=0.675 $Y=0.171
c86 69 VSS 3.13694e-19 $X=0.675 $Y=0.149
c87 68 VSS 0.00108989f $X=0.675 $Y=0.225
c88 66 VSS 7.23521e-19 $X=0.675 $Y=0.1125
c89 65 VSS 0.00101735f $X=0.675 $Y=0.099
c90 64 VSS 0.0011573f $X=0.675 $Y=0.081
c91 63 VSS 0.00104754f $X=0.675 $Y=0.063
c92 62 VSS 5.67204e-19 $X=0.675 $Y=0.126
c93 60 VSS 0.00330674f $X=0.63 $Y=0.234
c94 59 VSS 0.0075595f $X=0.666 $Y=0.234
c95 58 VSS 9.25907e-19 $X=0.621 $Y=0.225
c96 56 VSS 0.00286272f $X=0.63 $Y=0.036
c97 55 VSS 0.00687824f $X=0.608 $Y=0.036
c98 53 VSS 0.00282724f $X=0.54 $Y=0.036
c99 50 VSS 0.00757274f $X=0.666 $Y=0.036
c100 49 VSS 0.00363572f $X=0.608 $Y=0.198
c101 48 VSS 5.17397e-19 $X=0.576 $Y=0.198
c102 47 VSS 1.38834e-19 $X=0.558 $Y=0.198
c103 46 VSS 1.63363e-19 $X=0.554 $Y=0.198
c104 45 VSS 0.00129855f $X=0.522 $Y=0.198
c105 44 VSS 0.00152244f $X=0.485 $Y=0.198
c106 43 VSS 8.46035e-21 $X=0.414 $Y=0.198
c107 42 VSS 0.00390607f $X=0.396 $Y=0.198
c108 41 VSS 6.15423e-19 $X=0.325 $Y=0.198
c109 40 VSS 4.75287e-19 $X=0.288 $Y=0.198
c110 39 VSS 1.43629e-19 $X=0.252 $Y=0.198
c111 38 VSS 7.77903e-19 $X=0.612 $Y=0.198
c112 37 VSS 2.24414e-20 $X=0.243 $Y=0.18
c113 36 VSS 3.03855e-19 $X=0.243 $Y=0.171
c114 34 VSS 3.66662e-19 $X=0.243 $Y=0.126
c115 33 VSS 5.82045e-20 $X=0.243 $Y=0.189
c116 31 VSS 0.00295586f $X=0.216 $Y=0.2025
c117 27 VSS 5.87574e-19 $X=0.233 $Y=0.2025
c118 22 VSS 7.12523e-19 $X=0.557 $Y=0.0675
c119 20 VSS 0.00580086f $X=0.214 $Y=0.054
c120 13 VSS 0.00681065f $X=0.783 $Y=0.135
c121 10 VSS 0.0647446f $X=0.783 $Y=0.0675
c122 2 VSS 0.0652872f $X=0.729 $Y=0.0675
r123 96 97 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.2385 $Y2=0.072
r124 95 97 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.072 $X2=0.2385 $Y2=0.072
r125 90 96 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.072 $X2=0.234 $Y2=0.072
r126 87 88 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.2385 $Y2=0.198
r127 86 88 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.198 $X2=0.2385 $Y2=0.198
r128 81 87 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.234 $Y2=0.198
r129 73 99 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.135 $X2=0.675 $Y2=0.135
r130 73 75 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.135 $X2=0.729 $Y2=0.135
r131 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.189 $X2=0.675 $Y2=0.207
r132 70 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.171 $X2=0.675 $Y2=0.189
r133 69 70 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.149 $X2=0.675 $Y2=0.171
r134 68 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.225 $X2=0.675 $Y2=0.207
r135 67 99 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.144 $X2=0.675 $Y2=0.135
r136 67 69 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.144 $X2=0.675 $Y2=0.149
r137 65 66 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.099 $X2=0.675 $Y2=0.1125
r138 64 65 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.081 $X2=0.675 $Y2=0.099
r139 63 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.063 $X2=0.675 $Y2=0.081
r140 62 99 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.126 $X2=0.675 $Y2=0.135
r141 62 66 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.126 $X2=0.675 $Y2=0.1125
r142 61 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.045 $X2=0.675 $Y2=0.063
r143 59 68 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.234 $X2=0.675 $Y2=0.225
r144 59 60 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.234 $X2=0.63 $Y2=0.234
r145 58 60 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.621 $Y=0.225 $X2=0.63 $Y2=0.234
r146 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.207 $X2=0.621 $Y2=0.225
r147 55 56 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.608
+ $Y=0.036 $X2=0.63 $Y2=0.036
r148 52 55 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.608 $Y2=0.036
r149 52 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r150 50 61 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.036 $X2=0.675 $Y2=0.045
r151 50 56 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.63 $Y2=0.036
r152 48 49 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.198 $X2=0.608 $Y2=0.198
r153 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.198 $X2=0.576 $Y2=0.198
r154 46 47 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.554
+ $Y=0.198 $X2=0.558 $Y2=0.198
r155 45 46 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.198 $X2=0.554 $Y2=0.198
r156 44 45 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.485
+ $Y=0.198 $X2=0.522 $Y2=0.198
r157 43 44 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.485 $Y2=0.198
r158 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.414 $Y2=0.198
r159 41 42 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.325
+ $Y=0.198 $X2=0.396 $Y2=0.198
r160 40 41 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.325 $Y2=0.198
r161 39 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.243 $Y2=0.198
r162 39 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.288 $Y2=0.198
r163 38 57 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.198 $X2=0.621 $Y2=0.207
r164 38 49 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.198 $X2=0.608 $Y2=0.198
r165 36 37 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.171 $X2=0.243 $Y2=0.18
r166 35 36 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.144 $X2=0.243 $Y2=0.171
r167 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.144
r168 33 86 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.198
r169 33 37 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.18
r170 32 95 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.072
r171 32 34 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.126
r172 31 81 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198
+ $X2=0.216 $Y2=0.198
r173 28 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r174 27 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r175 26 53 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r176 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r177 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r178 20 90 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072
+ $X2=0.216 $Y2=0.072
r179 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.054 $X2=0.214 $Y2=0.054
r180 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.135 $X2=0.783 $Y2=0.2025
r181 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.135
r182 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.135 $X2=0.783 $Y2=0.135
r183 5 75 3.03549 $a=6.48e-16 $layer=V0LIG $count=2 $X=0.729 $Y=0.135 $X2=0.729
+ $Y2=0.135
r184 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.135 $X2=0.729 $Y2=0.2025
r185 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0675 $X2=0.729 $Y2=0.135
.ends

.subckt PM_AO31X2_ASAP7_75T_L%Y 1 2 6 7 16 23 28 29 30 VSS
c11 32 VSS 0.00271925f $X=0.837 $Y=0.1845
c12 30 VSS 1.052e-19 $X=0.837 $Y=0.1285
c13 29 VSS 0.00476898f $X=0.837 $Y=0.126
c14 28 VSS 6.35132e-19 $X=0.839 $Y=0.131
c15 26 VSS 0.0023684f $X=0.837 $Y=0.225
c16 24 VSS 0.00294383f $X=0.8125 $Y=0.036
c17 23 VSS 0.00552654f $X=0.797 $Y=0.036
c18 21 VSS 0.00904121f $X=0.756 $Y=0.036
c19 18 VSS 0.00579105f $X=0.828 $Y=0.036
c20 17 VSS 0.00294383f $X=0.8125 $Y=0.234
c21 16 VSS 0.00557175f $X=0.797 $Y=0.234
c22 11 VSS 0.00579156f $X=0.828 $Y=0.234
c23 10 VSS 0.00904119f $X=0.756 $Y=0.2025
c24 6 VSS 5.61153e-19 $X=0.773 $Y=0.2025
c25 1 VSS 5.72268e-19 $X=0.773 $Y=0.0675
r26 31 32 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.144 $X2=0.837 $Y2=0.1845
r27 29 30 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.126 $X2=0.837 $Y2=0.1285
r28 28 31 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.131 $X2=0.837 $Y2=0.144
r29 28 30 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.131 $X2=0.837 $Y2=0.1285
r30 26 32 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.1845
r31 25 29 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.045 $X2=0.837 $Y2=0.126
r32 23 24 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.797
+ $Y=0.036 $X2=0.8125 $Y2=0.036
r33 20 23 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.797 $Y2=0.036
r34 20 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r35 18 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.036 $X2=0.837 $Y2=0.045
r36 18 24 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.8125 $Y2=0.036
r37 16 17 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.797
+ $Y=0.234 $X2=0.8125 $Y2=0.234
r38 13 16 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.797 $Y2=0.234
r39 11 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r40 11 17 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.8125 $Y2=0.234
r41 10 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234 $X2=0.756
+ $Y2=0.234
r42 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r43 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r44 5 21 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.756
+ $Y=0.0675 $X2=0.756 $Y2=0.036
r45 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
r46 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
.ends


* END of "./AO31x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO31x2_ASAP7_75t_L  VSS VDD A3 B A2 A1 Y
* 
* Y	Y
* A1	A1
* A2	A2
* B	B
* A3	A3
M0 noxref_9 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_9 N_A3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_7_M2_d N_B_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 noxref_9 N_A2_M3_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 noxref_9 N_A2_M4_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M5 N_7_M5_d N_A1_M5_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_A1_M6_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M7 N_Y_M7_d N_7_M7_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M8 N_Y_M8_d N_7_M8_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773 $Y=0.027
M9 VDD N_A3_M9_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M10 VDD N_A3_M10_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M11 N_7_M11_d N_B_M11_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M12 N_7_M12_d N_B_M12_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M13 noxref_8 N_A2_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M14 noxref_8 N_A2_M14_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M15 noxref_8 N_A1_M15_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M16 noxref_8 N_A1_M16_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M17 N_Y_M17_d N_7_M17_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M18 N_Y_M18_d N_7_M18_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
*
* 
* .include "AO31x2_ASAP7_75t_L.pex.sp.AO31X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO31x2_ASAP7_75t_L.pex.sp.AO31X2_ASAP7_75T_L.pxi"
* File: AO31x2_ASAP7_75t_L.pex.sp.AO31X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:05:26 2017
* 
x_PM_AO31X2_ASAP7_75T_L%A3 N_A3_M0_g N_A3_M9_g N_A3_M1_g N_A3_c_4_p N_A3_M10_g
+ A3 VSS PM_AO31X2_ASAP7_75T_L%A3
x_PM_AO31X2_ASAP7_75T_L%B N_B_M2_g N_B_M11_g N_B_c_21_n N_B_M12_g B VSS
+ PM_AO31X2_ASAP7_75T_L%B
x_PM_AO31X2_ASAP7_75T_L%A2 N_A2_M3_g N_A2_M13_g N_A2_M4_g N_A2_c_52_p N_A2_M14_g
+ A2 VSS PM_AO31X2_ASAP7_75T_L%A2
x_PM_AO31X2_ASAP7_75T_L%A1 N_A1_M5_g N_A1_M15_g N_A1_M6_g N_A1_c_85_n N_A1_M16_g
+ A1 VSS PM_AO31X2_ASAP7_75T_L%A1
x_PM_AO31X2_ASAP7_75T_L%7 N_7_M7_g N_7_M17_g N_7_M8_g N_7_c_176_p N_7_M18_g
+ N_7_M2_d N_7_c_111_n N_7_M6_d N_7_M5_d N_7_M12_d N_7_M11_d N_7_c_113_n
+ N_7_c_114_n N_7_c_116_n N_7_c_118_n N_7_c_151_p N_7_c_127_n N_7_c_128_n
+ N_7_c_129_n N_7_c_131_n N_7_c_135_n N_7_c_137_n N_7_c_139_n N_7_c_175_p
+ N_7_c_182_p N_7_c_141_n N_7_c_143_n N_7_c_179_p N_7_c_158_p N_7_c_144_n
+ N_7_c_168_p N_7_c_172_p N_7_c_169_p N_7_c_145_n N_7_c_180_p N_7_c_120_n
+ N_7_c_122_n N_7_c_133_n N_7_c_146_n VSS PM_AO31X2_ASAP7_75T_L%7
x_PM_AO31X2_ASAP7_75T_L%Y N_Y_M8_d N_Y_M7_d N_Y_M18_d N_Y_M17_d N_Y_c_189_n
+ N_Y_c_192_n Y N_Y_c_195_n N_Y_c_196_n VSS PM_AO31X2_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_B_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.054
cc_2 N_A3_M1_g N_B_M2_g 0.00323392f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.054
cc_3 N_A3_M1_g N_B_c_21_n 2.69148e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_4 N_A3_c_4_p N_B_c_21_n 0.00149358f $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_5 N_A3_M1_g B 5.93459e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.134
cc_6 N_A3_c_4_p B 0.0032047f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.134
cc_7 A3 B 0.002207f $X=0.08 $Y=0.136 $X2=0.189 $Y2=0.134
cc_8 VSS A3 2.23359e-19 $X=0.08 $Y=0.136 $X2=0.189 $Y2=0.054
cc_9 VSS A3 0.00225004f $X=0.08 $Y=0.136 $X2=0.189 $Y2=0.135
cc_10 VSS A3 0.00179824f $X=0.08 $Y=0.136 $X2=0 $Y2=0
cc_11 VSS N_A3_M0_g 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_12 VSS N_A3_c_4_p 3.08494e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_13 VSS A3 2.73034e-19 $X=0.08 $Y=0.136 $X2=0 $Y2=0
cc_14 VSS N_A3_M1_g 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 VSS N_A3_c_4_p 3.80277e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.054
cc_16 VSS A3 5.97636e-19 $X=0.08 $Y=0.136 $X2=0.243 $Y2=0.2025
cc_17 VSS N_A3_c_4_p 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.2025
cc_18 VSS N_A3_M1_g 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 N_B_c_21_n N_7_c_111_n 3.82299e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_20 N_B_c_21_n N_7_M12_d 3.80413e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_21 N_B_c_21_n N_7_c_113_n 9.18375e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_22 N_B_c_21_n N_7_c_114_n 7.54008e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_23 B N_7_c_114_n 6.4382e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_24 N_B_c_21_n N_7_c_116_n 0.00127415f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_25 B N_7_c_116_n 8.41056e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_26 N_B_c_21_n N_7_c_118_n 4.86057e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_27 B N_7_c_118_n 5.36365e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_28 N_B_c_21_n N_7_c_120_n 4.65864e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_29 B N_7_c_120_n 3.81366e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_30 N_B_c_21_n N_7_c_122_n 4.18066e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 B N_7_c_122_n 3.7129e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_32 VSS B 0.0015422f $X=0.189 $Y=0.134 $X2=0.135 $Y2=0.0675
cc_33 VSS B 0.00375052f $X=0.189 $Y=0.134 $X2=0.081 $Y2=0.135
cc_34 VSS B 9.80823e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_35 VSS N_B_M2_g 4.23295e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_36 VSS N_B_c_21_n 2.28374e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_37 VSS B 0.002132f $X=0.189 $Y=0.134 $X2=0.135 $Y2=0.135
cc_38 VSS B 0.00374737f $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_39 VSS N_B_M2_g 4.28653e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_40 VSS B 0.00100241f $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_41 VSS N_B_c_21_n 2.34993e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_42 N_A2_M3_g N_A1_M5_g 2.74891e-19 $X=0.405 $Y=0.0675 $X2=0.189 $Y2=0.054
cc_43 N_A2_M4_g N_A1_M5_g 0.00335739f $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.054
cc_44 N_A2_M4_g N_A1_M6_g 2.74891e-19 $X=0.459 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_45 N_A2_c_52_p N_A1_c_85_n 0.00134829f $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.2025
cc_46 A2 A1 9.98825e-19 $X=0.403 $Y=0.137 $X2=0.189 $Y2=0.135
cc_47 A2 N_7_c_114_n 0.00122088f $X=0.403 $Y=0.137 $X2=0.243 $Y2=0.135
cc_48 A2 N_7_c_116_n 0.00122088f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_49 A2 N_7_c_118_n 0.00122088f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_50 A2 N_7_c_127_n 0.00473421f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_51 A2 N_7_c_128_n 9.41469e-19 $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_52 N_A2_M3_g N_7_c_129_n 3.08685e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_53 A2 N_7_c_129_n 7.78596e-19 $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_54 N_A2_M4_g N_7_c_131_n 3.99641e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_55 N_A2_c_52_p N_7_c_131_n 7.95511e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_56 A2 N_7_c_133_n 0.00122088f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_57 VSS A2 3.23443e-19 $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_58 VSS N_A2_c_52_p 3.80246e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_59 VSS N_A2_c_52_p 8.00061e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_60 VSS N_A2_M3_g 2.38303e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_61 VSS N_A2_M4_g 2.64781e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_62 VSS N_A2_c_52_p 3.80246e-19 $X=0.459 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_63 VSS N_A2_M3_g 2.38303e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_64 VSS A2 9.86796e-19 $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_65 VSS N_A2_c_52_p 8.00061e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_66 VSS A2 3.28046e-19 $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_67 VSS A2 0.0012344f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_68 VSS A2 9.86796e-19 $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_69 VSS A2 2.07179e-19 $X=0.403 $Y=0.137 $X2=0.189 $Y2=0.054
cc_70 VSS A2 0.00218013f $X=0.403 $Y=0.137 $X2=0.189 $Y2=0.135
cc_71 VSS N_A2_M3_g 2.52885e-19 $X=0.405 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_72 VSS A2 0.00473602f $X=0.403 $Y=0.137 $X2=0.189 $Y2=0.135
cc_73 VSS N_A2_c_52_p 7.92563e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_74 VSS N_A2_M4_g 4.95023e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_75 N_A1_c_85_n N_7_M6_d 3.76312e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_76 N_A1_M5_g N_7_c_135_n 2.56447e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_77 A1 N_7_c_135_n 0.00374659f $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_78 N_A1_c_85_n N_7_c_137_n 4.6296e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_79 A1 N_7_c_137_n 6.90614e-19 $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_80 N_A1_M6_g N_7_c_139_n 3.8357e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_81 A1 N_7_c_139_n 7.68517e-19 $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_82 N_A1_c_85_n N_7_c_141_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_83 A1 N_7_c_141_n 0.00135416f $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_84 N_A1_M6_g N_7_c_143_n 2.38303e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_85 A1 N_7_c_144_n 2.70873e-19 $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_86 A1 N_7_c_145_n 2.70873e-19 $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_87 A1 N_7_c_146_n 2.70873e-19 $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_88 VSS N_A1_c_85_n 3.80246e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_89 VSS N_A1_c_85_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_90 VSS A1 3.21662e-19 $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_91 VSS N_A1_M5_g 2.38303e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_92 VSS A1 3.24853e-19 $X=0.569 $Y=0.137 $X2=0.459 $Y2=0.0675
cc_93 VSS A1 3.21676e-19 $X=0.569 $Y=0.137 $X2=0.459 $Y2=0.2025
cc_94 VSS A1 4.01534e-19 $X=0.569 $Y=0.137 $X2=0.405 $Y2=0.135
cc_95 VSS N_A1_M5_g 3.4229e-19 $X=0.513 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_96 VSS A1 0.00335398f $X=0.569 $Y=0.137 $X2=0.405 $Y2=0.135
cc_97 VSS N_A1_M6_g 2.52885e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_98 VSS A1 0.00335398f $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_99 VSS N_7_c_113_n 0.00392515f $X=0.216 $Y=0.2025 $X2=0.135 $Y2=0.0675
cc_100 VSS N_7_c_120_n 4.02834e-19 $X=0.216 $Y=0.198 $X2=0.135 $Y2=0.0675
cc_101 VSS N_7_c_113_n 0.00356257f $X=0.216 $Y=0.2025 $X2=0.135 $Y2=0.2025
cc_102 VSS N_7_c_118_n 5.87812e-19 $X=0.243 $Y=0.171 $X2=0.135 $Y2=0.2025
cc_103 VSS N_7_c_151_p 0.00294986f $X=0.288 $Y=0.198 $X2=0.135 $Y2=0.2025
cc_104 VSS N_7_c_131_n 0.00226064f $X=0.485 $Y=0.198 $X2=0 $Y2=0
cc_105 VSS N_7_c_137_n 0.00217957f $X=0.554 $Y=0.198 $X2=0.08 $Y2=0.136
cc_106 VSS N_7_c_141_n 0.00131461f $X=0.54 $Y=0.036 $X2=0.08 $Y2=0.136
cc_107 VSS N_7_c_113_n 0.00249183f $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_108 VSS N_7_c_120_n 0.0145f $X=0.216 $Y=0.198 $X2=0 $Y2=0
cc_109 VSS N_7_c_127_n 0.0145f $X=0.325 $Y=0.198 $X2=0 $Y2=0
cc_110 VSS N_7_c_158_p 3.94426e-19 $X=0.63 $Y=0.234 $X2=0 $Y2=0
cc_111 VSS N_7_c_143_n 3.14186e-19 $X=0.608 $Y=0.036 $X2=0 $Y2=0
cc_112 VSS N_7_c_111_n 0.0032087f $X=0.214 $Y=0.054 $X2=0 $Y2=0
cc_113 VSS N_7_c_122_n 0.00480914f $X=0.216 $Y=0.072 $X2=0 $Y2=0
cc_114 VSS N_7_c_151_p 2.36616e-19 $X=0.288 $Y=0.198 $X2=0 $Y2=0
cc_115 VSS N_7_c_128_n 2.36616e-19 $X=0.396 $Y=0.198 $X2=0.08 $Y2=0.136
cc_116 VSS N_7_c_141_n 0.00332785f $X=0.54 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_117 VSS N_7_c_143_n 4.46182e-19 $X=0.608 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_118 VSS N_7_c_141_n 0.0037002f $X=0.54 $Y=0.036 $X2=0.135 $Y2=0.2025
cc_119 VSS N_7_c_143_n 0.00313249f $X=0.608 $Y=0.036 $X2=0.135 $Y2=0.2025
cc_120 VSS N_7_c_168_p 2.68628e-19 $X=0.675 $Y=0.063 $X2=0.135 $Y2=0.2025
cc_121 VSS N_7_c_169_p 4.06163e-19 $X=0.675 $Y=0.099 $X2=0.135 $Y2=0.2025
cc_122 VSS N_7_c_128_n 3.03534e-19 $X=0.396 $Y=0.198 $X2=0 $Y2=0
cc_123 VSS N_7_c_131_n 3.03534e-19 $X=0.485 $Y=0.198 $X2=0 $Y2=0
cc_124 VSS N_7_c_172_p 6.1248e-19 $X=0.675 $Y=0.081 $X2=0.081 $Y2=0.135
cc_125 VSS N_7_c_141_n 0.00238933f $X=0.54 $Y=0.036 $X2=0 $Y2=0
cc_126 VSS N_7_c_143_n 0.00678112f $X=0.608 $Y=0.036 $X2=0 $Y2=0
cc_127 VSS N_7_c_175_p 3.03534e-19 $X=0.608 $Y=0.198 $X2=0 $Y2=0
cc_128 N_7_c_176_p N_Y_M8_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_129 N_7_c_176_p N_Y_M18_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_130 N_7_M8_g N_Y_c_189_n 4.28653e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_131 N_7_c_179_p N_Y_c_189_n 3.90216e-19 $X=0.666 $Y=0.234 $X2=0 $Y2=0
cc_132 N_7_c_180_p N_Y_c_189_n 7.7415e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_133 N_7_M8_g N_Y_c_192_n 4.28653e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_134 N_7_c_182_p N_Y_c_192_n 3.9751e-19 $X=0.666 $Y=0.036 $X2=0 $Y2=0
cc_135 N_7_c_180_p N_Y_c_192_n 7.56738e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_136 N_7_c_172_p N_Y_c_195_n 3.17816e-19 $X=0.675 $Y=0.081 $X2=0.081 $Y2=0.135
cc_137 N_7_c_176_p N_Y_c_196_n 5.11279e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_138 N_7_c_180_p N_Y_c_196_n 0.00102f $X=0.729 $Y=0.135 $X2=0 $Y2=0

* END of "./AO31x2_ASAP7_75t_L.pex.sp.AO31X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO322x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:05:49 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO322x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO322x2_ASAP7_75t_L.pex.sp.pex"
* File: AO322x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:05:49 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO322X2_ASAP7_75T_L%A1 2 5 7 17 21 VSS
c11 21 VSS 0.00164036f $X=0.081 $Y=0.135
c12 17 VSS 0.0180882f $X=0.0505 $Y=0.1385
c13 5 VSS 0.00274291f $X=0.081 $Y=0.135
c14 2 VSS 0.0621257f $X=0.081 $Y=0.0675
r15 17 21 2.07099 $w=1.8e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.0505
+ $Y=0.135 $X2=0.081 $Y2=0.135
r16 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO322X2_ASAP7_75T_L%A2 2 5 7 12 17 24 29 VSS
c17 29 VSS 6.00769e-19 $X=0.1355 $Y=0.1905
c18 24 VSS 5.87439e-19 $X=0.135 $Y=0.198
c19 19 VSS 4.34718e-19 $X=0.135 $Y=0.18
c20 18 VSS 3.43106e-19 $X=0.135 $Y=0.171
c21 17 VSS 2.2242e-19 $X=0.135 $Y=0.164
c22 12 VSS 0.00104151f $X=0.135 $Y=0.135
c23 10 VSS 4.20973e-19 $X=0.135 $Y=0.189
c24 5 VSS 0.00116811f $X=0.135 $Y=0.135
c25 2 VSS 0.0576817f $X=0.135 $Y=0.0675
r26 24 29 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.198 $X2=0.1355 $Y2=0.198
r27 18 19 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.171 $X2=0.135 $Y2=0.18
r28 17 18 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.164 $X2=0.135 $Y2=0.171
r29 16 17 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.164
r30 12 16 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r31 10 24 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.135 $Y2=0.198
r32 10 19 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.135 $Y2=0.18
r33 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r34 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r35 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO322X2_ASAP7_75T_L%A3 2 5 7 10 VSS
c11 10 VSS 7.12602e-19 $X=0.1885 $Y=0.0905
c12 5 VSS 0.00108938f $X=0.189 $Y=0.135
c13 2 VSS 0.0577177f $X=0.189 $Y=0.0675
r14 10 13 3.02161 $w=1.8e-08 $l=4.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.0905 $X2=0.189 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO322X2_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c11 10 VSS 0.00107235f $X=0.243 $Y=0.135
c12 5 VSS 0.00114557f $X=0.243 $Y=0.135
c13 2 VSS 0.058856f $X=0.243 $Y=0.054
r14 10 14 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.1505
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO322X2_ASAP7_75T_L%B1 2 5 7 12 14 VSS
c15 14 VSS 5.36833e-19 $X=0.297 $Y=0.135
c16 12 VSS 0.00119714f $X=0.2995 $Y=0.0865
c17 5 VSS 0.00206319f $X=0.297 $Y=0.135
c18 2 VSS 0.0634905f $X=0.297 $Y=0.054
r19 12 14 3.29321 $w=1.8e-08 $l=4.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.0865 $X2=0.297 $Y2=0.135
r20 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r21 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r22 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO322X2_ASAP7_75T_L%C1 2 5 7 10 VSS
c8 10 VSS 0.00124462f $X=0.4585 $Y=0.0825
c9 5 VSS 0.00184379f $X=0.459 $Y=0.135
c10 2 VSS 0.063921f $X=0.459 $Y=0.054
r11 10 13 3.56481 $w=1.8e-08 $l=5.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.0825 $X2=0.459 $Y2=0.135
r12 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r14 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.054 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AO322X2_ASAP7_75T_L%C2 2 5 7 11 16 VSS
c8 11 VSS 0.00497173f $X=0.513 $Y=0.135
c9 5 VSS 0.00189109f $X=0.513 $Y=0.135
c10 2 VSS 0.063464f $X=0.513 $Y=0.054
r11 11 16 1.12037 $w=1.8e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.1515
r12 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r14 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.054 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AO322X2_ASAP7_75T_L%10 2 7 10 13 15 17 22 25 27 30 32 35 37 40 42 44
+ 45 52 54 55 56 57 58 59 60 61 66 67 68 69 71 80 81 83 88 90 92 95 99 VSS
c56 102 VSS 9.9667e-19 $X=0.423 $Y=0.036
c57 101 VSS 0.00203534f $X=0.414 $Y=0.036
c58 99 VSS 0.00313874f $X=0.432 $Y=0.036
c59 95 VSS 5.05467e-19 $X=0.6545 $Y=0.135
c60 94 VSS 0.00491915f $X=0.634 $Y=0.135
c61 92 VSS 6.14176e-19 $X=0.675 $Y=0.135
c62 90 VSS 0.00110556f $X=0.576 $Y=0.135
c63 89 VSS 9.26504e-20 $X=0.567 $Y=0.1765
c64 88 VSS 5.85687e-19 $X=0.567 $Y=0.164
c65 87 VSS 8.89444e-20 $X=0.567 $Y=0.189
c66 85 VSS 3.94527e-19 $X=0.5495 $Y=0.198
c67 84 VSS 0.00111453f $X=0.541 $Y=0.198
c68 83 VSS 5.31938e-19 $X=0.522 $Y=0.198
c69 82 VSS 2.34042e-19 $X=0.504 $Y=0.198
c70 81 VSS 5.47206e-19 $X=0.5 $Y=0.198
c71 80 VSS 8.46035e-21 $X=0.468 $Y=0.198
c72 79 VSS 1.22834e-19 $X=0.45 $Y=0.198
c73 78 VSS 4.17733e-19 $X=0.446 $Y=0.198
c74 71 VSS 4.5273e-19 $X=0.414 $Y=0.198
c75 70 VSS 0.00174591f $X=0.558 $Y=0.198
c76 69 VSS 3.86556e-20 $X=0.405 $Y=0.171
c77 68 VSS 2.07969e-19 $X=0.405 $Y=0.164
c78 67 VSS 0.00193608f $X=0.405 $Y=0.153
c79 66 VSS 2.79537e-19 $X=0.405 $Y=0.081
c80 65 VSS 3.16111e-19 $X=0.405 $Y=0.07
c81 64 VSS 3.82671e-20 $X=0.405 $Y=0.063
c82 63 VSS 6.69116e-20 $X=0.405 $Y=0.189
c83 61 VSS 0.00134427f $X=0.338 $Y=0.036
c84 60 VSS 0.00287092f $X=0.325 $Y=0.036
c85 59 VSS 0.00364813f $X=0.288 $Y=0.036
c86 58 VSS 0.00142296f $X=0.252 $Y=0.036
c87 57 VSS 0.00663192f $X=0.234 $Y=0.036
c88 56 VSS 0.00142296f $X=0.198 $Y=0.036
c89 55 VSS 0.00375557f $X=0.18 $Y=0.036
c90 54 VSS 0.00308768f $X=0.144 $Y=0.036
c91 53 VSS 0.00144693f $X=0.107 $Y=0.036
c92 52 VSS 0.00368527f $X=0.095 $Y=0.036
c93 45 VSS 0.00343598f $X=0.054 $Y=0.036
c94 44 VSS 0.00191587f $X=0.054 $Y=0.036
c95 42 VSS 0.00709587f $X=0.396 $Y=0.036
c96 40 VSS 0.00215284f $X=0.538 $Y=0.2025
c97 35 VSS 0.0023045f $X=0.434 $Y=0.2025
c98 32 VSS 2.69461e-19 $X=0.449 $Y=0.2025
c99 30 VSS 0.00336564f $X=0.434 $Y=0.054
c100 27 VSS 2.98509e-19 $X=0.449 $Y=0.054
c101 25 VSS 0.00350329f $X=0.322 $Y=0.054
c102 17 VSS 3.33606e-19 $X=0.071 $Y=0.0675
c103 13 VSS 0.00935851f $X=0.729 $Y=0.135
c104 10 VSS 0.0661363f $X=0.729 $Y=0.0675
c105 2 VSS 0.0654521f $X=0.675 $Y=0.0675
r106 101 102 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.423 $Y2=0.036
r107 99 102 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.423 $Y2=0.036
r108 97 101 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.036 $X2=0.414 $Y2=0.036
r109 94 95 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.634
+ $Y=0.135 $X2=0.6545 $Y2=0.135
r110 92 95 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.135 $X2=0.6545 $Y2=0.135
r111 90 94 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.135 $X2=0.634 $Y2=0.135
r112 88 89 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.164 $X2=0.567 $Y2=0.1765
r113 87 89 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.567 $Y2=0.1765
r114 86 90 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.567 $Y=0.144 $X2=0.576 $Y2=0.135
r115 86 88 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.144 $X2=0.567 $Y2=0.164
r116 84 85 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.541
+ $Y=0.198 $X2=0.5495 $Y2=0.198
r117 82 83 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.198 $X2=0.522 $Y2=0.198
r118 81 82 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.5
+ $Y=0.198 $X2=0.504 $Y2=0.198
r119 80 81 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.198 $X2=0.5 $Y2=0.198
r120 79 80 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.198 $X2=0.468 $Y2=0.198
r121 78 79 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.446
+ $Y=0.198 $X2=0.45 $Y2=0.198
r122 76 84 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.198 $X2=0.541 $Y2=0.198
r123 76 83 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.198 $X2=0.522 $Y2=0.198
r124 73 78 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.433
+ $Y=0.198 $X2=0.446 $Y2=0.198
r125 71 73 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.433 $Y2=0.198
r126 70 87 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.198 $X2=0.567 $Y2=0.189
r127 70 85 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.198 $X2=0.5495 $Y2=0.198
r128 68 69 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.164 $X2=0.405 $Y2=0.171
r129 67 68 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.405 $Y2=0.164
r130 66 67 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.081 $X2=0.405 $Y2=0.153
r131 65 66 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.07 $X2=0.405 $Y2=0.081
r132 64 65 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.063 $X2=0.405 $Y2=0.07
r133 63 71 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.405 $Y=0.189 $X2=0.414 $Y2=0.198
r134 63 69 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.171
r135 62 97 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.036
r136 62 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.063
r137 60 61 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.325
+ $Y=0.036 $X2=0.338 $Y2=0.036
r138 58 59 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r139 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r140 56 57 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.234 $Y2=0.036
r141 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r142 54 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.18 $Y2=0.036
r143 53 54 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.036 $X2=0.144 $Y2=0.036
r144 52 53 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.036 $X2=0.107 $Y2=0.036
r145 50 60 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.325 $Y2=0.036
r146 50 59 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.288 $Y2=0.036
r147 44 52 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.095 $Y2=0.036
r148 44 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r149 42 97 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.405 $Y2=0.036
r150 42 61 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.338 $Y2=0.036
r151 40 76 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.198 $X2=0.54
+ $Y2=0.198
r152 37 40 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.538 $Y2=0.2025
r153 35 73 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.433 $Y=0.198
+ $X2=0.433 $Y2=0.198
r154 32 35 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.434 $Y2=0.2025
r155 30 99 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r156 27 30 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.054 $X2=0.434 $Y2=0.054
r157 25 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r158 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.054 $X2=0.322 $Y2=0.054
r159 20 45 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.054 $Y=0.0675 $X2=0.054 $Y2=0.036
r160 17 20 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r161 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.135 $X2=0.729 $Y2=0.2025
r162 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.135
r163 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.729 $Y2=0.135
r164 5 92 3.03549 $a=6.48e-16 $layer=V0LIG $count=2 $X=0.675 $Y=0.135 $X2=0.675
+ $Y2=0.135
r165 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.2025
r166 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0675 $X2=0.675 $Y2=0.135
.ends

.subckt PM_AO322X2_ASAP7_75T_L%Y 1 6 11 14 16 24 29 39 44 48 49 VSS
c16 50 VSS 4.55454e-19 $X=0.783 $Y=0.216
c17 49 VSS 0.00307026f $X=0.783 $Y=0.207
c18 48 VSS 7.46953e-19 $X=0.783 $Y=0.144
c19 46 VSS 6.70981e-19 $X=0.783 $Y=0.081
c20 45 VSS 8.85605e-19 $X=0.783 $Y=0.063
c21 44 VSS 0.00249415f $X=0.7835 $Y=0.1145
c22 42 VSS 4.30151e-19 $X=0.783 $Y=0.225
c23 40 VSS 6.22498e-19 $X=0.7495 $Y=0.234
c24 39 VSS 0.0124703f $X=0.743 $Y=0.234
c25 31 VSS 0.00581326f $X=0.774 $Y=0.234
c26 30 VSS 6.22498e-19 $X=0.7495 $Y=0.036
c27 29 VSS 0.0126189f $X=0.743 $Y=0.036
c28 28 VSS 0.00635284f $X=0.756 $Y=0.036
c29 24 VSS 0.00678229f $X=0.648 $Y=0.036
c30 21 VSS 0.00581326f $X=0.774 $Y=0.036
c31 19 VSS 0.0066597f $X=0.754 $Y=0.2025
c32 14 VSS 0.00569926f $X=0.65 $Y=0.2025
c33 11 VSS 3.33606e-19 $X=0.665 $Y=0.2025
c34 9 VSS 3.06859e-19 $X=0.754 $Y=0.0675
c35 1 VSS 3.33606e-19 $X=0.665 $Y=0.0675
r36 49 50 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.207 $X2=0.783 $Y2=0.216
r37 48 49 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.144 $X2=0.783 $Y2=0.207
r38 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.126 $X2=0.783 $Y2=0.144
r39 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.063 $X2=0.783 $Y2=0.081
r40 44 47 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.1145 $X2=0.783 $Y2=0.126
r41 44 46 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.1145 $X2=0.783 $Y2=0.081
r42 42 50 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.225 $X2=0.783 $Y2=0.216
r43 41 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.063
r44 39 40 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.743
+ $Y=0.234 $X2=0.7495 $Y2=0.234
r45 37 40 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.7495 $Y2=0.234
r46 33 39 6.45062 $w=1.8e-08 $l=9.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.743 $Y2=0.234
r47 31 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.774 $Y=0.234 $X2=0.783 $Y2=0.225
r48 31 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.234 $X2=0.756 $Y2=0.234
r49 29 30 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.743
+ $Y=0.036 $X2=0.7495 $Y2=0.036
r50 27 30 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.7495 $Y2=0.036
r51 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r52 23 29 6.45062 $w=1.8e-08 $l=9.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.743 $Y2=0.036
r53 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036 $X2=0.648
+ $Y2=0.036
r54 21 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.774 $Y=0.036 $X2=0.783 $Y2=0.045
r55 21 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.036 $X2=0.756 $Y2=0.036
r56 19 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234 $X2=0.756
+ $Y2=0.234
r57 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.754 $Y2=0.2025
r58 14 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234 $X2=0.648
+ $Y2=0.234
r59 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.65 $Y2=0.2025
r60 9 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.756
+ $Y=0.0675 $X2=0.756 $Y2=0.036
r61 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.0675 $X2=0.754 $Y2=0.0675
r62 4 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.648
+ $Y=0.0675 $X2=0.648 $Y2=0.036
r63 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.665
+ $Y=0.0675 $X2=0.65 $Y2=0.0675
.ends


* END of "./AO322x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO322x2_ASAP7_75t_L  VSS VDD A1 A2 A3 B2 B1 C1 C2 Y
* 
* Y	Y
* C2	C2
* C1	C1
* B1	B1
* B2	B2
* A3	A3
* A2	A2
* A1	A1
M0 noxref_14 N_A1_M0_g N_10_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_15 N_A2_M1_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_A3_M2_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_16 N_B2_M3_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 N_10_M4_d N_B1_M4_g noxref_16 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.027
M5 noxref_17 N_C1_M5_g N_10_M5_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.449
+ $Y=0.027
M6 VSS N_C2_M6_g noxref_17 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.503
+ $Y=0.027
M7 VSS N_10_M7_g N_Y_M7_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M8 VSS N_10_M8_g N_Y_M8_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M9 noxref_11 N_A1_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M10 VDD N_A2_M10_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M11 noxref_11 N_A3_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M12 noxref_12 N_B2_M12_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M13 noxref_11 N_B1_M13_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M14 noxref_12 N_C1_M14_g N_10_M14_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M15 N_10_M15_d N_C2_M15_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
M16 VDD N_10_M16_g N_Y_M16_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
M17 VDD N_10_M17_g N_Y_M17_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
*
* 
* .include "AO322x2_ASAP7_75t_L.pex.sp.AO322X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO322x2_ASAP7_75t_L.pex.sp.AO322X2_ASAP7_75T_L.pxi"
* File: AO322x2_ASAP7_75t_L.pex.sp.AO322X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:05:49 2017
* 
x_PM_AO322X2_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M9_g A1 N_A1_c_4_p VSS
+ PM_AO322X2_ASAP7_75T_L%A1
x_PM_AO322X2_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_13_n N_A2_M10_g N_A2_c_14_n
+ N_A2_c_16_n N_A2_c_25_p A2 VSS PM_AO322X2_ASAP7_75T_L%A2
x_PM_AO322X2_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_31_n N_A3_M11_g A3 VSS
+ PM_AO322X2_ASAP7_75T_L%A3
x_PM_AO322X2_ASAP7_75T_L%B2 N_B2_M3_g N_B2_c_42_n N_B2_M12_g N_B2_c_43_n B2 VSS
+ PM_AO322X2_ASAP7_75T_L%B2
x_PM_AO322X2_ASAP7_75T_L%B1 N_B1_M4_g N_B1_c_53_n N_B1_M13_g B1 N_B1_c_59_p VSS
+ PM_AO322X2_ASAP7_75T_L%B1
x_PM_AO322X2_ASAP7_75T_L%C1 N_C1_M5_g N_C1_c_67_p N_C1_M14_g C1 VSS
+ PM_AO322X2_ASAP7_75T_L%C1
x_PM_AO322X2_ASAP7_75T_L%C2 N_C2_M6_g N_C2_c_75_n N_C2_M15_g N_C2_c_76_n C2 VSS
+ PM_AO322X2_ASAP7_75T_L%C2
x_PM_AO322X2_ASAP7_75T_L%10 N_10_M7_g N_10_M16_g N_10_M8_g N_10_c_127_p
+ N_10_M17_g N_10_M0_s N_10_M4_d N_10_c_93_n N_10_M5_s N_10_c_99_n N_10_M14_s
+ N_10_c_108_p N_10_M15_d N_10_c_115_p N_10_c_122_p N_10_c_82_n N_10_c_83_n
+ N_10_c_84_n N_10_c_87_n N_10_c_137_p N_10_c_89_n N_10_c_111_p N_10_c_91_n
+ N_10_c_112_p N_10_c_94_n N_10_c_113_p N_10_c_100_n N_10_c_96_n N_10_c_97_n
+ N_10_c_98_n N_10_c_110_p N_10_c_101_n N_10_c_116_p N_10_c_103_n N_10_c_105_n
+ N_10_c_106_n N_10_c_135_p N_10_c_128_p N_10_c_129_p VSS
+ PM_AO322X2_ASAP7_75T_L%10
x_PM_AO322X2_ASAP7_75T_L%Y N_Y_M7_s N_Y_M8_s N_Y_M16_s N_Y_c_139_n N_Y_M17_s
+ N_Y_c_138_n N_Y_c_141_n N_Y_c_146_n Y N_Y_c_150_n N_Y_c_152_n VSS
+ PM_AO322X2_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00335986f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_13_n 0.00120928f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A1 N_A2_c_14_n 9.90974e-19 $X=0.0505 $Y=0.1385 $X2=0.135 $Y2=0.135
cc_4 N_A1_c_4_p N_A2_c_14_n 8.78098e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_5 A1 N_A2_c_16_n 4.6841e-19 $X=0.0505 $Y=0.1385 $X2=0.135 $Y2=0.164
cc_6 N_A1_M0_g N_A3_M2_g 2.48122e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_7 A1 N_10_c_82_n 0.00119499f $X=0.0505 $Y=0.1385 $X2=0 $Y2=0
cc_8 A1 N_10_c_83_n 0.00208198f $X=0.0505 $Y=0.1385 $X2=0 $Y2=0
cc_9 N_A1_M0_g N_10_c_84_n 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_10 N_A1_c_4_p N_10_c_84_n 2.97176e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 VSS A1 5.24213e-19 $X=0.0505 $Y=0.1385 $X2=0.135 $Y2=0.171
cc_12 N_A2_M1_g N_A3_M2_g 0.00304756f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_13 N_A2_c_13_n N_A3_c_31_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 N_A2_c_14_n A3 0.00455283f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_15 N_A2_M1_g N_B2_M3_g 2.13359e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_A2_c_14_n N_10_c_83_n 0.00137201f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_17 N_A2_M1_g N_10_c_87_n 3.22844e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_18 N_A2_c_14_n N_10_c_87_n 0.00398146f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_19 VSS N_A2_c_16_n 9.20487e-19 $X=0.135 $Y=0.164 $X2=0.081 $Y2=0.135
cc_20 VSS N_A2_c_25_p 0.00119567f $X=0.135 $Y=0.198 $X2=0.081 $Y2=0.135
cc_21 VSS N_A2_M1_g 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_22 VSS N_A2_c_25_p 0.00372455f $X=0.135 $Y=0.198 $X2=0 $Y2=0
cc_23 VSS A2 7.4424e-19 $X=0.1355 $Y=0.1905 $X2=0 $Y2=0
cc_24 N_A3_M2_g N_B2_M3_g 0.00304756f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_25 N_A3_c_31_n N_B2_c_42_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_26 A3 N_B2_c_43_n 0.00406615f $X=0.1885 $Y=0.0905 $X2=0 $Y2=0
cc_27 N_A3_M2_g N_B1_M4_g 2.48122e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_28 N_A3_M2_g N_10_c_89_n 2.56935e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_29 A3 N_10_c_89_n 0.00123064f $X=0.1885 $Y=0.0905 $X2=0 $Y2=0
cc_30 VSS A3 0.00159458f $X=0.1885 $Y=0.0905 $X2=0 $Y2=0
cc_31 N_B2_M3_g N_B1_M4_g 0.00348334f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.0675
cc_32 N_B2_c_42_n N_B1_c_53_n 9.33263e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_33 N_B2_c_43_n B1 0.00460879f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_34 N_B2_M3_g N_10_c_91_n 2.56935e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_35 N_B2_c_43_n N_10_c_91_n 0.00123064f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_36 VSS N_B2_M3_g 3.62029e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_37 VSS N_B2_c_43_n 0.0012322f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_38 B1 N_10_c_93_n 0.00178959f $X=0.2995 $Y=0.0865 $X2=0 $Y2=0
cc_39 N_B1_M4_g N_10_c_94_n 2.34993e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_40 B1 N_10_c_94_n 0.00374072f $X=0.2995 $Y=0.0865 $X2=0 $Y2=0
cc_41 B1 N_10_c_96_n 0.00125528f $X=0.2995 $Y=0.0865 $X2=0 $Y2=0
cc_42 N_B1_c_59_p N_10_c_97_n 2.02971e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_43 N_B1_c_59_p N_10_c_98_n 2.02971e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_44 VSS N_B1_c_59_p 9.98224e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_45 VSS N_B1_M4_g 2.52885e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_46 VSS N_B1_c_59_p 0.0037392f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_47 VSS N_B1_c_59_p 3.03401e-19 $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.135
cc_48 VSS N_B1_M4_g 2.38303e-19 $X=0.297 $Y=0.054 $X2=0.135 $Y2=0.171
cc_49 N_C1_M5_g N_C2_M6_g 0.00353416f $X=0.459 $Y=0.054 $X2=0.513 $Y2=0.054
cc_50 N_C1_c_67_p N_C2_c_75_n 9.79748e-19 $X=0.459 $Y=0.135 $X2=0.513 $Y2=0.135
cc_51 C1 N_C2_c_76_n 0.00473083f $X=0.4585 $Y=0.0825 $X2=0.513 $Y2=0.135
cc_52 C1 N_10_c_99_n 3.87865e-19 $X=0.4585 $Y=0.0825 $X2=0 $Y2=0
cc_53 C1 N_10_c_100_n 0.00440084f $X=0.4585 $Y=0.0825 $X2=0 $Y2=0
cc_54 N_C1_M5_g N_10_c_101_n 2.68514e-19 $X=0.459 $Y=0.054 $X2=0 $Y2=0
cc_55 C1 N_10_c_101_n 0.00121543f $X=0.4585 $Y=0.0825 $X2=0 $Y2=0
cc_56 VSS N_C1_M5_g 2.38303e-19 $X=0.459 $Y=0.054 $X2=0.5145 $Y2=0.1515
cc_57 N_C2_M6_g N_10_c_103_n 3.62029e-19 $X=0.513 $Y=0.054 $X2=0 $Y2=0
cc_58 N_C2_c_76_n N_10_c_103_n 0.00123353f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_59 N_C2_c_76_n N_10_c_105_n 8.25345e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_60 N_C2_c_76_n N_10_c_106_n 8.25345e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_61 N_C2_c_76_n N_Y_c_138_n 5.10273e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_62 VSS N_10_c_93_n 7.03295e-19 $X=0.322 $Y=0.054 $X2=0 $Y2=0
cc_63 VSS N_10_c_108_p 0.00138601f $X=0.434 $Y=0.2025 $X2=0 $Y2=0
cc_64 VSS N_10_c_97_n 3.57339e-19 $X=0.405 $Y=0.164 $X2=0 $Y2=0
cc_65 VSS N_10_c_110_p 7.29421e-19 $X=0.414 $Y=0.198 $X2=0 $Y2=0
cc_66 VSS N_10_c_111_p 2.24129e-19 $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_67 VSS N_10_c_112_p 2.24129e-19 $X=0.288 $Y=0.036 $X2=0 $Y2=0
cc_68 VSS N_10_c_113_p 2.24129e-19 $X=0.338 $Y=0.036 $X2=0 $Y2=0
cc_69 VSS N_10_c_108_p 0.00385141f $X=0.434 $Y=0.2025 $X2=0 $Y2=0
cc_70 VSS N_10_c_115_p 0.00353266f $X=0.538 $Y=0.2025 $X2=0 $Y2=0
cc_71 VSS N_10_c_116_p 0.00239497f $X=0.5 $Y=0.198 $X2=0 $Y2=0
cc_72 VSS N_10_M14_s 3.13602e-19 $X=0.449 $Y=0.2025 $X2=0.0505 $Y2=0.135
cc_73 VSS N_10_c_108_p 0.00279124f $X=0.434 $Y=0.2025 $X2=0.0505 $Y2=0.135
cc_74 VSS N_10_c_115_p 5.10383e-19 $X=0.538 $Y=0.2025 $X2=0.0505 $Y2=0.135
cc_75 VSS N_10_c_110_p 0.00915527f $X=0.414 $Y=0.198 $X2=0.0505 $Y2=0.135
cc_76 VSS N_10_c_113_p 3.36552e-19 $X=0.338 $Y=0.036 $X2=0 $Y2=0
cc_77 VSS N_10_c_122_p 3.36552e-19 $X=0.396 $Y=0.036 $X2=0 $Y2=0
cc_78 N_10_c_115_p N_Y_c_139_n 0.00161971f $X=0.538 $Y=0.2025 $X2=0 $Y2=0
cc_79 N_10_c_105_n N_Y_c_139_n 8.72414e-19 $X=0.567 $Y=0.164 $X2=0 $Y2=0
cc_80 N_10_M7_g N_Y_c_141_n 4.28653e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_81 N_10_M8_g N_Y_c_141_n 4.28653e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_82 N_10_c_127_p N_Y_c_141_n 2.72752e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_83 N_10_c_128_p N_Y_c_141_n 0.00178689f $X=0.6545 $Y=0.135 $X2=0 $Y2=0
cc_84 N_10_c_129_p N_Y_c_141_n 2.07029e-19 $X=0.432 $Y=0.036 $X2=0 $Y2=0
cc_85 N_10_M7_g N_Y_c_146_n 4.28653e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_86 N_10_M8_g N_Y_c_146_n 4.28653e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_87 N_10_c_127_p N_Y_c_146_n 2.72752e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_88 N_10_c_128_p N_Y_c_146_n 0.0017263f $X=0.6545 $Y=0.135 $X2=0 $Y2=0
cc_89 N_10_c_127_p N_Y_c_150_n 5.06061e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_90 N_10_c_135_p N_Y_c_150_n 0.00103954f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_91 N_10_c_105_n N_Y_c_152_n 2.14189e-19 $X=0.567 $Y=0.164 $X2=0 $Y2=0
cc_92 VSS N_10_c_137_p 3.56327e-19 $X=0.18 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_93 VSS N_Y_c_146_n 2.63455e-19 $X=0.486 $Y=0.234 $X2=0 $Y2=0

* END of "./AO322x2_ASAP7_75t_L.pex.sp.AO322X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO32x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:06:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO32x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO32x1_ASAP7_75t_L.pex.sp.pex"
* File: AO32x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:06:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO32X1_ASAP7_75T_L%3 2 5 7 10 11 18 19 22 24 26 28 31 33 35 36 37 38
+ 42 45 51 52 53 58 60 VSS
c33 66 VSS 6.49054e-19 $X=0.09 $Y=0.135
c34 65 VSS 7.57725e-19 $X=0.099 $Y=0.135
c35 60 VSS 2.18493e-19 $X=0.076 $Y=0.135
c36 58 VSS 0.00420379f $X=0.405 $Y=0.164
c37 57 VSS 0.00114479f $X=0.405 $Y=0.07
c38 56 VSS 0.00132122f $X=0.405 $Y=0.189
c39 54 VSS 1.7098e-19 $X=0.394 $Y=0.198
c40 53 VSS 6.15718e-19 $X=0.392 $Y=0.198
c41 52 VSS 8.46035e-21 $X=0.36 $Y=0.198
c42 51 VSS 5.02599e-19 $X=0.342 $Y=0.198
c43 46 VSS 0.00201526f $X=0.396 $Y=0.198
c44 45 VSS 0.00146362f $X=0.36 $Y=0.036
c45 44 VSS 0.0030651f $X=0.342 $Y=0.036
c46 43 VSS 5.63812e-19 $X=0.31 $Y=0.036
c47 42 VSS 0.00142296f $X=0.306 $Y=0.036
c48 41 VSS 0.00131785f $X=0.288 $Y=0.036
c49 40 VSS 0.00142154f $X=0.276 $Y=0.036
c50 39 VSS 0.00103073f $X=0.261 $Y=0.036
c51 38 VSS 0.00142296f $X=0.252 $Y=0.036
c52 37 VSS 0.00350351f $X=0.234 $Y=0.036
c53 36 VSS 0.00142296f $X=0.198 $Y=0.036
c54 35 VSS 0.00312443f $X=0.18 $Y=0.036
c55 34 VSS 3.78291e-19 $X=0.148 $Y=0.036
c56 33 VSS 0.00146362f $X=0.144 $Y=0.036
c57 32 VSS 0.00294815f $X=0.126 $Y=0.036
c58 31 VSS 0.00316377f $X=0.27 $Y=0.036
c59 28 VSS 0.00270205f $X=0.108 $Y=0.036
c60 27 VSS 0.00907412f $X=0.396 $Y=0.036
c61 26 VSS 2.58269e-19 $X=0.099 $Y=0.081
c62 25 VSS 0.00127834f $X=0.099 $Y=0.07
c63 24 VSS 0.00134156f $X=0.099 $Y=0.126
c64 22 VSS 0.00221162f $X=0.324 $Y=0.216
c65 18 VSS 5.70405e-19 $X=0.341 $Y=0.216
c66 12 VSS 5.36031e-19 $X=0.27 $Y=0.0455
c67 5 VSS 0.00418456f $X=0.081 $Y=0.135
c68 2 VSS 0.0658735f $X=0.081 $Y=0.0675
r69 66 67 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.135 $X2=0.0945 $Y2=0.135
r70 65 67 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.135 $X2=0.0945 $Y2=0.135
r71 60 66 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.076
+ $Y=0.135 $X2=0.09 $Y2=0.135
r72 57 58 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.07 $X2=0.405 $Y2=0.164
r73 56 58 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.164
r74 55 57 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.07
r75 53 54 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.392
+ $Y=0.198 $X2=0.394 $Y2=0.198
r76 52 53 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.198 $X2=0.392 $Y2=0.198
r77 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r78 48 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.342 $Y2=0.198
r79 46 56 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.198 $X2=0.405 $Y2=0.189
r80 46 54 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.394 $Y2=0.198
r81 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r82 43 44 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.31
+ $Y=0.036 $X2=0.342 $Y2=0.036
r83 42 43 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.31 $Y2=0.036
r84 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r85 40 41 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.276
+ $Y=0.036 $X2=0.288 $Y2=0.036
r86 38 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.261 $Y2=0.036
r87 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r88 36 37 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.234 $Y2=0.036
r89 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r90 34 35 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.036 $X2=0.18 $Y2=0.036
r91 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.148 $Y2=0.036
r92 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r93 30 40 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.276 $Y2=0.036
r94 30 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.261 $Y2=0.036
r95 30 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r96 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r97 27 55 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r98 27 45 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.36 $Y2=0.036
r99 25 26 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.07 $X2=0.099 $Y2=0.081
r100 24 65 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.126 $X2=0.099 $Y2=0.135
r101 24 26 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.126 $X2=0.099 $Y2=0.081
r102 23 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.099 $Y=0.045 $X2=0.108 $Y2=0.036
r103 23 25 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.045 $X2=0.099 $Y2=0.07
r104 22 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198
+ $X2=0.324 $Y2=0.198
r105 19 22 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.216 $X2=0.324 $Y2=0.216
r106 18 22 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.216 $X2=0.324 $Y2=0.216
r107 17 31 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r108 11 12 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0455 $X2=0.27 $Y2=0.0455
r109 10 12 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0455 $X2=0.27 $Y2=0.0455
r110 9 17 3.12934 $w=6.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.27 $Y=0.064 $X2=0.253 $Y2=0.064
r111 9 12 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.27 $Y=0.064 $X2=0.27 $Y2=0.0455
r112 5 60 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.076 $Y=0.135 $X2=0.076
+ $Y2=0.135
r113 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r114 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO32X1_ASAP7_75T_L%A3 2 5 7 10 14 16 VSS
c11 16 VSS 1.37595e-19 $X=0.135 $Y=0.15975
c12 14 VSS 0.00155051f $X=0.137 $Y=0.1755
c13 10 VSS 2.70559e-19 $X=0.135 $Y=0.135
c14 5 VSS 0.001283f $X=0.135 $Y=0.135
c15 2 VSS 0.0598272f $X=0.135 $Y=0.0675
r16 15 16 1.06944 $w=1.8e-08 $l=1.575e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.15975
r17 14 16 1.06944 $w=1.8e-08 $l=1.575e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.1755 $X2=0.135 $Y2=0.15975
r18 10 15 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r19 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r20 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r21 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO32X1_ASAP7_75T_L%A2 2 5 7 10 VSS
c13 10 VSS 8.20834e-19 $X=0.189 $Y=0.1295
c14 5 VSS 0.00106592f $X=0.189 $Y=0.135
c15 2 VSS 0.059998f $X=0.189 $Y=0.0675
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO32X1_ASAP7_75T_L%A1 2 5 7 11 15 VSS
c15 17 VSS 1.49585e-19 $X=0.243 $Y=0.17025
c16 15 VSS 0.00172294f $X=0.248 $Y=0.1765
c17 11 VSS 3.33833e-19 $X=0.243 $Y=0.135
c18 5 VSS 0.0010782f $X=0.243 $Y=0.135
c19 2 VSS 0.0608182f $X=0.243 $Y=0.0675
r20 16 17 0.424383 $w=1.8e-08 $l=6.25e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.164 $X2=0.243 $Y2=0.17025
r21 15 17 0.424383 $w=1.8e-08 $l=6.25e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.1765 $X2=0.243 $Y2=0.17025
r22 11 16 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.164
r23 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r24 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r25 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO32X1_ASAP7_75T_L%B1 2 5 7 10 VSS
c12 10 VSS 5.05734e-19 $X=0.297 $Y=0.1195
c13 5 VSS 0.00113686f $X=0.297 $Y=0.135
c14 2 VSS 0.0621713f $X=0.297 $Y=0.054
r15 10 13 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1195 $X2=0.297 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO32X1_ASAP7_75T_L%B2 2 5 7 13 VSS
c10 13 VSS 8.26297e-19 $X=0.354 $Y=0.1345
c11 5 VSS 0.00170409f $X=0.351 $Y=0.135
c12 2 VSS 0.0655438f $X=0.351 $Y=0.054
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.216
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.054 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AO32X1_ASAP7_75T_L%Y 1 6 14 15 16 21 25 28 VSS
c6 28 VSS 0.00526409f $X=0.054 $Y=0.049
c7 25 VSS 0.00524642f $X=0.018 $Y=0.063
c8 21 VSS 0.00537134f $X=0.054 $Y=0.234
c9 19 VSS 0.00316555f $X=0.027 $Y=0.234
c10 18 VSS 2.379e-19 $X=0.018 $Y=0.207
c11 16 VSS 7.35763e-19 $X=0.018 $Y=0.144
c12 15 VSS 0.00212552f $X=0.018 $Y=0.126
c13 14 VSS 0.00265661f $X=0.017 $Y=0.1755
c14 12 VSS 5.9475e-19 $X=0.018 $Y=0.225
c15 9 VSS 0.00581009f $X=0.056 $Y=0.2025
c16 6 VSS 4.92917e-19 $X=0.071 $Y=0.2025
c17 1 VSS 5.15148e-19 $X=0.071 $Y=0.0675
r18 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.049 $X2=0.054
+ $Y2=0.049
r19 25 27 1.6 $w=2.75e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.054 $Y2=0.063
r20 19 21 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.054 $Y2=0.234
r21 17 18 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.207
r22 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.144
r23 14 17 1.66358 $w=1.8e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1755 $X2=0.018 $Y2=0.2
r24 14 16 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1755 $X2=0.018 $Y2=0.144
r25 12 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r26 12 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.207
r27 11 25 0.322338 $w=2.75e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.063
r28 11 15 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.126
r29 9 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r30 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
r31 4 28 15.9673 $w=2.4e-08 $l=1.85e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.049
r32 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./AO32x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO32x1_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 Y
* 
* Y	Y
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 VSS N_3_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 noxref_11 N_A3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_12 N_A2_M2_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_3_M3_d N_A1_M3_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_13 N_B1_M4_g N_3_M4_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.027
M5 VSS N_B2_M5_g noxref_13 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341
+ $Y=0.027
M6 VDD N_3_M6_g N_Y_M6_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M7 noxref_10 N_A3_M7_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M8 VDD N_A2_M8_g noxref_10 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M9 noxref_10 N_A1_M9_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M10 N_3_M10_d N_B1_M10_g noxref_10 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.287 $Y=0.189
M11 noxref_10 N_B2_M11_g N_3_M11_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.341 $Y=0.189
*
* 
* .include "AO32x1_ASAP7_75t_L.pex.sp.AO32X1_ASAP7_75T_L.pxi"
* BEGIN of "./AO32x1_ASAP7_75t_L.pex.sp.AO32X1_ASAP7_75T_L.pxi"
* File: AO32x1_ASAP7_75t_L.pex.sp.AO32X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:06:11 2017
* 
x_PM_AO32X1_ASAP7_75T_L%3 N_3_M0_g N_3_c_3_p N_3_M6_g N_3_M4_s N_3_M3_d
+ N_3_M11_s N_3_M10_d N_3_c_25_p N_3_c_21_p N_3_c_4_p N_3_c_23_p N_3_c_10_p
+ N_3_c_2_p N_3_c_32_p N_3_c_7_p N_3_c_33_p N_3_c_9_p N_3_c_13_p N_3_c_16_p
+ N_3_c_12_p N_3_c_17_p N_3_c_29_p N_3_c_20_p N_3_c_22_p VSS
+ PM_AO32X1_ASAP7_75T_L%3
x_PM_AO32X1_ASAP7_75T_L%A3 N_A3_M1_g N_A3_c_36_n N_A3_M7_g N_A3_c_37_n A3
+ N_A3_c_43_p VSS PM_AO32X1_ASAP7_75T_L%A3
x_PM_AO32X1_ASAP7_75T_L%A2 N_A2_M2_g N_A2_c_49_n N_A2_M8_g A2 VSS
+ PM_AO32X1_ASAP7_75T_L%A2
x_PM_AO32X1_ASAP7_75T_L%A1 N_A1_M3_g N_A1_c_64_n N_A1_M9_g N_A1_c_59_n A1 VSS
+ PM_AO32X1_ASAP7_75T_L%A1
x_PM_AO32X1_ASAP7_75T_L%B1 N_B1_M4_g N_B1_c_78_n N_B1_M10_g B1 VSS
+ PM_AO32X1_ASAP7_75T_L%B1
x_PM_AO32X1_ASAP7_75T_L%B2 N_B2_M5_g N_B2_c_92_n N_B2_M11_g B2 VSS
+ PM_AO32X1_ASAP7_75T_L%B2
x_PM_AO32X1_ASAP7_75T_L%Y N_Y_M0_s N_Y_M6_s Y N_Y_c_95_n N_Y_c_96_n N_Y_c_100_p
+ N_Y_c_97_n N_Y_c_98_n VSS PM_AO32X1_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M1_g 0.00287079f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_3_c_2_p N_A3_M1_g 2.64276e-19 $X=0.144 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_3 N_3_c_3_p N_A3_c_36_n 0.0011052f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_3_c_4_p N_A3_c_37_n 0.00612129f $X=0.099 $Y=0.081 $X2=0.135 $Y2=0.135
cc_5 N_3_c_2_p N_A3_c_37_n 0.00125352f $X=0.144 $Y=0.036 $X2=0.135 $Y2=0.135
cc_6 N_3_M0_g N_A2_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_7 N_3_c_7_p N_A2_M2_g 3.38929e-19 $X=0.198 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_8 N_3_c_7_p A2 0.00123604f $X=0.198 $Y=0.036 $X2=0.135 $Y2=0.135
cc_9 N_3_c_9_p N_A1_M3_g 2.56935e-19 $X=0.252 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_10 N_3_c_10_p N_A1_c_59_n 0.0013295f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.135
cc_11 N_3_c_9_p N_A1_c_59_n 0.00123678f $X=0.252 $Y=0.036 $X2=0.135 $Y2=0.135
cc_12 N_3_c_12_p A1 7.93475e-19 $X=0.342 $Y=0.198 $X2=0.135 $Y2=0.144
cc_13 N_3_c_13_p N_B1_M4_g 2.56935e-19 $X=0.306 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_14 N_3_c_10_p B1 0.00133251f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.135
cc_15 N_3_c_13_p B1 0.00123064f $X=0.306 $Y=0.036 $X2=0.135 $Y2=0.135
cc_16 N_3_c_16_p N_B2_M5_g 2.64276e-19 $X=0.36 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_17 N_3_c_17_p N_B2_M5_g 2.76185e-19 $X=0.36 $Y=0.198 $X2=0.135 $Y2=0.0675
cc_18 N_3_c_16_p B2 0.00124805f $X=0.36 $Y=0.036 $X2=0.135 $Y2=0.1755
cc_19 N_3_c_17_p B2 0.0012322f $X=0.36 $Y=0.198 $X2=0.135 $Y2=0.1755
cc_20 N_3_c_20_p B2 0.00446403f $X=0.405 $Y=0.164 $X2=0.135 $Y2=0.1755
cc_21 N_3_c_21_p N_Y_c_95_n 9.26167e-19 $X=0.099 $Y=0.126 $X2=0.135 $Y2=0.144
cc_22 N_3_c_22_p N_Y_c_96_n 7.90121e-19 $X=0.076 $Y=0.135 $X2=0.135 $Y2=0.15975
cc_23 N_3_c_23_p N_Y_c_97_n 0.00274492f $X=0.108 $Y=0.036 $X2=0 $Y2=0
cc_24 N_3_c_23_p N_Y_c_98_n 0.00135917f $X=0.108 $Y=0.036 $X2=0 $Y2=0
cc_25 VSS N_3_c_25_p 0.00288888f $X=0.324 $Y=0.216 $X2=0.135 $Y2=0.135
cc_26 VSS N_3_c_10_p 7.32217e-19 $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.135
cc_27 VSS N_3_c_12_p 2.56435e-19 $X=0.342 $Y=0.198 $X2=0.135 $Y2=0.135
cc_28 VSS N_3_c_25_p 0.00302498f $X=0.324 $Y=0.216 $X2=0.137 $Y2=0.1755
cc_29 VSS N_3_c_29_p 0.00393556f $X=0.392 $Y=0.198 $X2=0.137 $Y2=0.1755
cc_30 VSS N_3_c_25_p 0.00250965f $X=0.324 $Y=0.216 $X2=0 $Y2=0
cc_31 VSS N_3_c_12_p 0.0070721f $X=0.342 $Y=0.198 $X2=0 $Y2=0
cc_32 VSS N_3_c_32_p 4.57078e-19 $X=0.18 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_33 VSS N_3_c_33_p 4.8755e-19 $X=0.234 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_34 N_A3_M1_g N_A2_M2_g 0.00347357f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_35 N_A3_c_36_n N_A2_c_49_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_36 N_A3_c_37_n A2 0.00628398f $X=0.135 $Y=0.135 $X2=0.287 $Y2=0.0455
cc_37 N_A3_M1_g N_A1_M3_g 2.69148e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_38 N_A3_c_43_p Y 5.55023e-19 $X=0.135 $Y=0.15975 $X2=0 $Y2=0
cc_39 VSS A3 3.31541e-19 $X=0.137 $Y=0.1755 $X2=0.081 $Y2=0.135
cc_40 N_A2_M2_g N_A1_M3_g 0.00330657f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_41 N_A2_c_49_n N_A1_c_64_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_42 A2 N_A1_c_59_n 0.00625269f $X=0.189 $Y=0.1295 $X2=0.253 $Y2=0.0455
cc_43 N_A2_M2_g N_B1_M4_g 2.74891e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_44 VSS A2 3.31541e-19 $X=0.189 $Y=0.1295 $X2=0.081 $Y2=0.135
cc_45 VSS N_A2_M2_g 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0.099 $Y2=0.126
cc_46 VSS A2 0.00125352f $X=0.189 $Y=0.1295 $X2=0.099 $Y2=0.126
cc_47 N_A1_M3_g N_B1_M4_g 0.0036697f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_48 N_A1_c_64_n N_B1_c_78_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_49 N_A1_c_59_n B1 0.00383317f $X=0.243 $Y=0.135 $X2=0.287 $Y2=0.0455
cc_50 N_A1_M3_g N_B2_M5_g 3.03912e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_51 VSS A1 0.00221632f $X=0.248 $Y=0.1765 $X2=0.287 $Y2=0.0455
cc_52 VSS N_A1_M3_g 2.38303e-19 $X=0.243 $Y=0.0675 $X2=0.099 $Y2=0.081
cc_53 VSS A1 0.00413343f $X=0.248 $Y=0.1765 $X2=0.099 $Y2=0.081
cc_54 N_B1_M4_g N_B2_M5_g 0.0036697f $X=0.297 $Y=0.054 $X2=0.081 $Y2=0.0675
cc_55 N_B1_c_78_n N_B2_c_92_n 9.33263e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_56 B1 B2 0.00487321f $X=0.297 $Y=0.1195 $X2=0 $Y2=0
cc_57 VSS N_B1_M4_g 3.47199e-19 $X=0.297 $Y=0.054 $X2=0.126 $Y2=0.036
cc_58 VSS B1 5.30079e-19 $X=0.297 $Y=0.1195 $X2=0.126 $Y2=0.036
cc_59 VSS N_B2_M5_g 2.38303e-19 $X=0.351 $Y=0.054 $X2=0.108 $Y2=0.036
cc_60 VSS N_Y_c_100_p 2.79945e-19 $X=0.054 $Y=0.234 $X2=0.099 $Y2=0.045

* END of "./AO32x1_ASAP7_75t_L.pex.sp.AO32X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO32x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:06:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO32x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO32x2_ASAP7_75t_L.pex.sp.pex"
* File: AO32x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:06:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO32X2_ASAP7_75T_L%3 2 7 10 13 15 18 19 26 27 30 36 37 39 40 41 43 46
+ 48 50 51 52 53 57 60 66 67 68 73 VSS
c46 73 VSS 0.00420379f $X=0.459 $Y=0.164
c47 72 VSS 0.00114479f $X=0.459 $Y=0.07
c48 71 VSS 0.00132122f $X=0.459 $Y=0.189
c49 69 VSS 1.7098e-19 $X=0.448 $Y=0.198
c50 68 VSS 6.15718e-19 $X=0.446 $Y=0.198
c51 67 VSS 8.46035e-21 $X=0.414 $Y=0.198
c52 66 VSS 5.02599e-19 $X=0.396 $Y=0.198
c53 61 VSS 0.00201526f $X=0.45 $Y=0.198
c54 60 VSS 0.00146362f $X=0.414 $Y=0.036
c55 59 VSS 0.0030651f $X=0.396 $Y=0.036
c56 58 VSS 5.63812e-19 $X=0.364 $Y=0.036
c57 57 VSS 0.00142296f $X=0.36 $Y=0.036
c58 56 VSS 0.00131785f $X=0.342 $Y=0.036
c59 55 VSS 0.00142154f $X=0.33 $Y=0.036
c60 54 VSS 0.00103073f $X=0.315 $Y=0.036
c61 53 VSS 0.00142296f $X=0.306 $Y=0.036
c62 52 VSS 0.00350351f $X=0.288 $Y=0.036
c63 51 VSS 0.00142296f $X=0.252 $Y=0.036
c64 50 VSS 0.00312443f $X=0.234 $Y=0.036
c65 49 VSS 3.78291e-19 $X=0.202 $Y=0.036
c66 48 VSS 0.00146362f $X=0.198 $Y=0.036
c67 47 VSS 0.00294815f $X=0.18 $Y=0.036
c68 46 VSS 0.00316377f $X=0.324 $Y=0.036
c69 43 VSS 0.00270205f $X=0.162 $Y=0.036
c70 42 VSS 0.00907412f $X=0.45 $Y=0.036
c71 41 VSS 2.58269e-19 $X=0.153 $Y=0.081
c72 40 VSS 0.00127834f $X=0.153 $Y=0.07
c73 39 VSS 0.00123094f $X=0.153 $Y=0.126
c74 37 VSS 4.68643e-20 $X=0.122 $Y=0.135
c75 36 VSS 2.4063e-21 $X=0.117 $Y=0.135
c76 31 VSS 0.00151931f $X=0.144 $Y=0.135
c77 30 VSS 0.00221162f $X=0.378 $Y=0.216
c78 26 VSS 5.70405e-19 $X=0.395 $Y=0.216
c79 20 VSS 5.36031e-19 $X=0.324 $Y=0.0455
c80 13 VSS 0.00440286f $X=0.135 $Y=0.135
c81 10 VSS 0.0618812f $X=0.135 $Y=0.0675
c82 2 VSS 0.0645183f $X=0.081 $Y=0.0675
r83 72 73 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.07 $X2=0.459 $Y2=0.164
r84 71 73 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.189 $X2=0.459 $Y2=0.164
r85 70 72 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.07
r86 68 69 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.446
+ $Y=0.198 $X2=0.448 $Y2=0.198
r87 67 68 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.446 $Y2=0.198
r88 66 67 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.414 $Y2=0.198
r89 63 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.198 $X2=0.396 $Y2=0.198
r90 61 71 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.198 $X2=0.459 $Y2=0.189
r91 61 69 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.198 $X2=0.448 $Y2=0.198
r92 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r93 58 59 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.364
+ $Y=0.036 $X2=0.396 $Y2=0.036
r94 57 58 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.364 $Y2=0.036
r95 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r96 55 56 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.33
+ $Y=0.036 $X2=0.342 $Y2=0.036
r97 53 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.315 $Y2=0.036
r98 52 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r99 51 52 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r100 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r101 49 50 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.036 $X2=0.234 $Y2=0.036
r102 48 49 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.202 $Y2=0.036
r103 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r104 45 55 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.33 $Y2=0.036
r105 45 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.315 $Y2=0.036
r106 45 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r107 43 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r108 42 70 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r109 42 60 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.414 $Y2=0.036
r110 40 41 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.07 $X2=0.153 $Y2=0.081
r111 39 41 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.126 $X2=0.153 $Y2=0.081
r112 38 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.153 $Y=0.045 $X2=0.162 $Y2=0.036
r113 38 40 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.045 $X2=0.153 $Y2=0.07
r114 36 37 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.135 $X2=0.122 $Y2=0.135
r115 33 36 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.117 $Y2=0.135
r116 31 39 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.144 $Y=0.135 $X2=0.153 $Y2=0.126
r117 31 37 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.122 $Y2=0.135
r118 30 63 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.198
+ $X2=0.378 $Y2=0.198
r119 27 30 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.216 $X2=0.378 $Y2=0.216
r120 26 30 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.216 $X2=0.378 $Y2=0.216
r121 25 46 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r122 19 20 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0455 $X2=0.324 $Y2=0.0455
r123 18 20 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0455 $X2=0.324 $Y2=0.0455
r124 17 25 3.12934 $w=6.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.324 $Y=0.064 $X2=0.307 $Y2=0.064
r125 17 20 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.324 $Y=0.064 $X2=0.324 $Y2=0.0455
r126 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r127 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r128 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r129 5 33 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r130 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r131 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO32X2_ASAP7_75T_L%A3 2 5 7 10 14 16 VSS
c12 16 VSS 2.02574e-19 $X=0.189 $Y=0.15975
c13 14 VSS 0.00176071f $X=0.191 $Y=0.1755
c14 10 VSS 3.03777e-19 $X=0.189 $Y=0.135
c15 5 VSS 0.0011642f $X=0.189 $Y=0.135
c16 2 VSS 0.0590549f $X=0.189 $Y=0.0675
r17 15 16 1.06944 $w=1.8e-08 $l=1.575e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.15975
r18 14 16 1.06944 $w=1.8e-08 $l=1.575e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.1755 $X2=0.189 $Y2=0.15975
r19 10 15 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.144
r20 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r21 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO32X2_ASAP7_75T_L%A2 2 5 7 10 VSS
c13 10 VSS 8.20834e-19 $X=0.243 $Y=0.1295
c14 5 VSS 0.00106612f $X=0.243 $Y=0.135
c15 2 VSS 0.059998f $X=0.243 $Y=0.0675
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO32X2_ASAP7_75T_L%A1 2 5 7 11 15 VSS
c15 17 VSS 1.49585e-19 $X=0.297 $Y=0.17025
c16 15 VSS 0.00172294f $X=0.302 $Y=0.1765
c17 11 VSS 3.33833e-19 $X=0.297 $Y=0.135
c18 5 VSS 0.0010782f $X=0.297 $Y=0.135
c19 2 VSS 0.0608182f $X=0.297 $Y=0.0675
r20 16 17 0.424383 $w=1.8e-08 $l=6.25e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.164 $X2=0.297 $Y2=0.17025
r21 15 17 0.424383 $w=1.8e-08 $l=6.25e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1765 $X2=0.297 $Y2=0.17025
r22 11 16 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.164
r23 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r24 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r25 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO32X2_ASAP7_75T_L%B1 2 5 7 10 VSS
c12 10 VSS 5.05734e-19 $X=0.351 $Y=0.1195
c13 5 VSS 0.00113686f $X=0.351 $Y=0.135
c14 2 VSS 0.0621713f $X=0.351 $Y=0.054
r15 10 13 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1195 $X2=0.351 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.216
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.054 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AO32X2_ASAP7_75T_L%B2 2 5 7 13 VSS
c10 13 VSS 8.26297e-19 $X=0.408 $Y=0.1345
c11 5 VSS 0.00170409f $X=0.405 $Y=0.135
c12 2 VSS 0.0655438f $X=0.405 $Y=0.054
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.216
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.054 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO32X2_ASAP7_75T_L%Y 1 2 5 6 7 14 15 16 19 22 25 28 35 VSS
c18 35 VSS 0.00756933f $X=0.108 $Y=0.054
c19 28 VSS 0.00146362f $X=0.09 $Y=0.234
c20 27 VSS 0.00784882f $X=0.072 $Y=0.234
c21 25 VSS 0.00352975f $X=0.108 $Y=0.234
c22 23 VSS 0.00319564f $X=0.027 $Y=0.234
c23 22 VSS 7.72418e-19 $X=0.072 $Y=0.072
c24 21 VSS 0.0042436f $X=0.062 $Y=0.072
c25 20 VSS 0.00165989f $X=0.027 $Y=0.072
c26 19 VSS 1.63855e-19 $X=0.099 $Y=0.072
c27 18 VSS 4.40073e-19 $X=0.018 $Y=0.207
c28 16 VSS 7.45746e-19 $X=0.018 $Y=0.144
c29 15 VSS 0.00229372f $X=0.018 $Y=0.126
c30 14 VSS 0.00315626f $X=0.017 $Y=0.1755
c31 12 VSS 8.29409e-19 $X=0.018 $Y=0.225
c32 10 VSS 0.00916119f $X=0.108 $Y=0.2025
c33 6 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c34 5 VSS 0.0105145f $X=0.108 $Y=0.0675
c35 1 VSS 5.945e-19 $X=0.125 $Y=0.0675
r36 33 35 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.063 $X2=0.108 $Y2=0.054
r37 27 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r38 25 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.09 $Y2=0.234
r39 23 27 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.072 $Y2=0.234
r40 21 22 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.062
+ $Y=0.072 $X2=0.072 $Y2=0.072
r41 20 21 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.072 $X2=0.062 $Y2=0.072
r42 19 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.099 $Y=0.072 $X2=0.108 $Y2=0.063
r43 19 22 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.072 $X2=0.072 $Y2=0.072
r44 17 18 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.207
r45 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.144
r46 14 17 1.66358 $w=1.8e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1755 $X2=0.018 $Y2=0.2
r47 14 16 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1755 $X2=0.018 $Y2=0.144
r48 12 23 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r49 12 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.207
r50 11 20 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.081 $X2=0.027 $Y2=0.072
r51 11 15 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.126
r52 10 25 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r53 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r54 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r55 5 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.054 $X2=0.108
+ $Y2=0.054
r56 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r57 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./AO32x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO32x2_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 Y
* 
* Y	Y
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_11 N_A3_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_12 N_A2_M3_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_3_M4_d N_A1_M4_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_13 N_B1_M5_g N_3_M5_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341
+ $Y=0.027
M6 VSS N_B2_M6_g noxref_13 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.395
+ $Y=0.027
M7 N_Y_M7_d N_3_M7_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M8 N_Y_M8_d N_3_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M9 noxref_10 N_A3_M9_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M10 VDD N_A2_M10_g noxref_10 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M11 noxref_10 N_A1_M11_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.189
M12 N_3_M12_d N_B1_M12_g noxref_10 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.341 $Y=0.189
M13 noxref_10 N_B2_M13_g N_3_M13_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.395 $Y=0.189
*
* 
* .include "AO32x2_ASAP7_75t_L.pex.sp.AO32X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO32x2_ASAP7_75t_L.pex.sp.AO32X2_ASAP7_75T_L.pxi"
* File: AO32x2_ASAP7_75t_L.pex.sp.AO32X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:06:34 2017
* 
x_PM_AO32X2_ASAP7_75T_L%3 N_3_M0_g N_3_M7_g N_3_M1_g N_3_c_4_p N_3_M8_g N_3_M5_s
+ N_3_M4_d N_3_M13_s N_3_M12_d N_3_c_38_p N_3_c_27_p N_3_c_32_p N_3_c_26_p
+ N_3_c_36_p N_3_c_5_p N_3_c_23_p N_3_c_11_p N_3_c_3_p N_3_c_45_p N_3_c_8_p
+ N_3_c_46_p N_3_c_10_p N_3_c_14_p N_3_c_17_p N_3_c_13_p N_3_c_18_p N_3_c_42_p
+ N_3_c_21_p VSS PM_AO32X2_ASAP7_75T_L%3
x_PM_AO32X2_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_50_n N_A3_M9_g N_A3_c_51_n A3
+ N_A3_c_57_p VSS PM_AO32X2_ASAP7_75T_L%A3
x_PM_AO32X2_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_63_n N_A2_M10_g A2 VSS
+ PM_AO32X2_ASAP7_75T_L%A2
x_PM_AO32X2_ASAP7_75T_L%A1 N_A1_M4_g N_A1_c_78_n N_A1_M11_g N_A1_c_73_n A1 VSS
+ PM_AO32X2_ASAP7_75T_L%A1
x_PM_AO32X2_ASAP7_75T_L%B1 N_B1_M5_g N_B1_c_92_n N_B1_M12_g B1 VSS
+ PM_AO32X2_ASAP7_75T_L%B1
x_PM_AO32X2_ASAP7_75T_L%B2 N_B2_M6_g N_B2_c_106_n N_B2_M13_g B2 VSS
+ PM_AO32X2_ASAP7_75T_L%B2
x_PM_AO32X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_c_110_n N_Y_M8_d N_Y_M7_d Y
+ N_Y_c_112_n N_Y_c_114_n N_Y_c_115_n N_Y_c_118_n N_Y_c_119_n N_Y_c_120_n
+ N_Y_c_122_n VSS PM_AO32X2_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_A3_M2_g 0.00287079f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_A3_M2_g 2.64276e-19 $X=0.198 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_4 N_3_c_4_p N_A3_c_50_n 0.00108551f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_5 N_3_c_5_p N_A3_c_51_n 0.00611191f $X=0.153 $Y=0.081 $X2=0.189 $Y2=0.135
cc_6 N_3_c_3_p N_A3_c_51_n 0.00125352f $X=0.198 $Y=0.036 $X2=0.189 $Y2=0.135
cc_7 N_3_M1_g N_A2_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_8 N_3_c_8_p N_A2_M3_g 3.38929e-19 $X=0.252 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_9 N_3_c_8_p A2 0.00123604f $X=0.252 $Y=0.036 $X2=0.189 $Y2=0.135
cc_10 N_3_c_10_p N_A1_M4_g 2.56935e-19 $X=0.306 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_11 N_3_c_11_p N_A1_c_73_n 0.0013295f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.135
cc_12 N_3_c_10_p N_A1_c_73_n 0.00123678f $X=0.306 $Y=0.036 $X2=0.189 $Y2=0.135
cc_13 N_3_c_13_p A1 7.93475e-19 $X=0.396 $Y=0.198 $X2=0.189 $Y2=0.144
cc_14 N_3_c_14_p N_B1_M5_g 2.56935e-19 $X=0.36 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_15 N_3_c_11_p B1 0.00133251f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.135
cc_16 N_3_c_14_p B1 0.00123064f $X=0.36 $Y=0.036 $X2=0.189 $Y2=0.135
cc_17 N_3_c_17_p N_B2_M6_g 2.64276e-19 $X=0.414 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_18 N_3_c_18_p N_B2_M6_g 2.76185e-19 $X=0.414 $Y=0.198 $X2=0.189 $Y2=0.0675
cc_19 N_3_c_17_p B2 0.00124805f $X=0.414 $Y=0.036 $X2=0.189 $Y2=0.1755
cc_20 N_3_c_18_p B2 0.0012322f $X=0.414 $Y=0.198 $X2=0.189 $Y2=0.1755
cc_21 N_3_c_21_p B2 0.00446403f $X=0.459 $Y=0.164 $X2=0.189 $Y2=0.1755
cc_22 N_3_c_4_p N_Y_M1_d 3.8044e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_23 N_3_c_23_p N_Y_c_110_n 0.00123132f $X=0.162 $Y=0.036 $X2=0.189 $Y2=0.135
cc_24 N_3_c_4_p N_Y_M8_d 3.80218e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.216
cc_25 N_3_c_4_p N_Y_c_112_n 3.67406e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.144
cc_26 N_3_c_26_p N_Y_c_112_n 2.98624e-19 $X=0.153 $Y=0.126 $X2=0.189 $Y2=0.144
cc_27 N_3_c_27_p N_Y_c_114_n 5.88274e-19 $X=0.117 $Y=0.135 $X2=0.189 $Y2=0.15975
cc_28 N_3_M0_g N_Y_c_115_n 2.94632e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_29 N_3_c_27_p N_Y_c_115_n 0.00124156f $X=0.117 $Y=0.135 $X2=0 $Y2=0
cc_30 N_3_c_5_p N_Y_c_115_n 0.00110218f $X=0.153 $Y=0.081 $X2=0 $Y2=0
cc_31 N_3_c_4_p N_Y_c_118_n 2.00665e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_32 N_3_c_32_p N_Y_c_119_n 3.54274e-19 $X=0.122 $Y=0.135 $X2=0 $Y2=0
cc_33 N_3_M0_g N_Y_c_120_n 3.85788e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_34 N_3_c_27_p N_Y_c_120_n 3.54274e-19 $X=0.117 $Y=0.135 $X2=0 $Y2=0
cc_35 N_3_M0_g N_Y_c_122_n 2.24173e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_3_c_36_p N_Y_c_122_n 0.00110218f $X=0.153 $Y=0.07 $X2=0 $Y2=0
cc_37 N_3_c_23_p N_Y_c_122_n 0.00110218f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_38 VSS N_3_c_38_p 0.00288888f $X=0.378 $Y=0.216 $X2=0.189 $Y2=0.135
cc_39 VSS N_3_c_11_p 7.32217e-19 $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.135
cc_40 VSS N_3_c_13_p 2.56435e-19 $X=0.396 $Y=0.198 $X2=0.189 $Y2=0.135
cc_41 VSS N_3_c_38_p 0.00302498f $X=0.378 $Y=0.216 $X2=0.191 $Y2=0.1755
cc_42 VSS N_3_c_42_p 0.00393556f $X=0.446 $Y=0.198 $X2=0.191 $Y2=0.1755
cc_43 VSS N_3_c_38_p 0.00250965f $X=0.378 $Y=0.216 $X2=0 $Y2=0
cc_44 VSS N_3_c_13_p 0.0070721f $X=0.396 $Y=0.198 $X2=0 $Y2=0
cc_45 VSS N_3_c_45_p 4.57078e-19 $X=0.234 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_46 VSS N_3_c_46_p 4.8755e-19 $X=0.288 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_47 N_A3_M2_g N_A2_M3_g 0.00347357f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_48 N_A3_c_50_n N_A2_c_63_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_49 N_A3_c_51_n A2 0.00628398f $X=0.189 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_50 N_A3_M2_g N_A1_M4_g 2.69148e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_51 N_A3_c_57_p Y 2.86312e-19 $X=0.189 $Y=0.15975 $X2=0.135 $Y2=0.2025
cc_52 VSS A3 3.31541e-19 $X=0.191 $Y=0.1755 $X2=0.081 $Y2=0.135
cc_53 N_A2_M3_g N_A1_M4_g 0.00330657f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_54 N_A2_c_63_n N_A1_c_78_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_55 A2 N_A1_c_73_n 0.00625269f $X=0.243 $Y=0.1295 $X2=0 $Y2=0
cc_56 N_A2_M3_g N_B1_M5_g 2.74891e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_57 VSS A2 3.31541e-19 $X=0.243 $Y=0.1295 $X2=0.081 $Y2=0.135
cc_58 VSS N_A2_M3_g 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_59 VSS A2 0.00125352f $X=0.243 $Y=0.1295 $X2=0 $Y2=0
cc_60 N_A1_M4_g N_B1_M5_g 0.0036697f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_61 N_A1_c_78_n N_B1_c_92_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_62 N_A1_c_73_n B1 0.00383317f $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_63 N_A1_M4_g N_B2_M6_g 3.03912e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_64 VSS A1 0.00221632f $X=0.302 $Y=0.1765 $X2=0.135 $Y2=0.0675
cc_65 VSS N_A1_M4_g 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0.395 $Y2=0.216
cc_66 VSS A1 0.00413343f $X=0.302 $Y=0.1765 $X2=0.395 $Y2=0.216
cc_67 N_B1_M5_g N_B2_M6_g 0.0036697f $X=0.351 $Y=0.054 $X2=0.081 $Y2=0.0675
cc_68 N_B1_c_92_n N_B2_c_106_n 9.33263e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_69 B1 B2 0.00487321f $X=0.351 $Y=0.1195 $X2=0.135 $Y2=0.135
cc_70 VSS N_B1_M5_g 3.47199e-19 $X=0.351 $Y=0.054 $X2=0.081 $Y2=0.135
cc_71 VSS B1 5.30079e-19 $X=0.351 $Y=0.1195 $X2=0.081 $Y2=0.135
cc_72 VSS N_B2_M6_g 2.38303e-19 $X=0.405 $Y=0.054 $X2=0.378 $Y2=0.216
cc_73 VSS N_Y_c_119_n 2.92912e-19 $X=0.108 $Y=0.234 $X2=0.307 $Y2=0.064

* END of "./AO32x2_ASAP7_75t_L.pex.sp.AO32X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO331x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:06:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO331x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO331x1_ASAP7_75t_L.pex.sp.pex"
* File: AO331x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:06:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO331X1_ASAP7_75T_L%3 2 5 7 9 10 14 19 22 28 29 31 32 36 39 41 42 43
+ 44 48 50 52 53 54 55 56 58 64 66 72 VSS
c43 72 VSS 0.00385307f $X=0.504 $Y=0.234
c44 71 VSS 0.00278591f $X=0.513 $Y=0.234
c45 66 VSS 6.85875e-19 $X=0.513 $Y=0.207
c46 65 VSS 0.00104083f $X=0.513 $Y=0.189
c47 64 VSS 0.00414953f $X=0.513 $Y=0.164
c48 63 VSS 8.11244e-19 $X=0.513 $Y=0.07
c49 62 VSS 0.00102822f $X=0.513 $Y=0.225
c50 60 VSS 6.9735e-19 $X=0.4785 $Y=0.036
c51 59 VSS 2.39163e-19 $X=0.471 $Y=0.036
c52 58 VSS 0.00146362f $X=0.468 $Y=0.036
c53 57 VSS 2.39163e-19 $X=0.45 $Y=0.036
c54 56 VSS 0.00606761f $X=0.447 $Y=0.036
c55 55 VSS 0.00142296f $X=0.414 $Y=0.036
c56 54 VSS 0.00343941f $X=0.396 $Y=0.036
c57 53 VSS 0.00142296f $X=0.36 $Y=0.036
c58 52 VSS 0.00325376f $X=0.342 $Y=0.036
c59 51 VSS 1.47784e-19 $X=0.308 $Y=0.036
c60 50 VSS 0.00146362f $X=0.306 $Y=0.036
c61 49 VSS 0.00274887f $X=0.288 $Y=0.036
c62 48 VSS 0.00676142f $X=0.486 $Y=0.036
c63 45 VSS 0.00106181f $X=0.261 $Y=0.036
c64 44 VSS 0.00142296f $X=0.252 $Y=0.036
c65 43 VSS 0.0037673f $X=0.234 $Y=0.036
c66 42 VSS 0.00142296f $X=0.198 $Y=0.036
c67 41 VSS 0.00347922f $X=0.18 $Y=0.036
c68 40 VSS 1.51923e-19 $X=0.146 $Y=0.036
c69 39 VSS 0.00218387f $X=0.27 $Y=0.036
c70 36 VSS 0.00238538f $X=0.144 $Y=0.036
c71 35 VSS 0.00596382f $X=0.504 $Y=0.036
c72 34 VSS 4.29035e-19 $X=0.135 $Y=0.063
c73 32 VSS 3.49137e-19 $X=0.09 $Y=0.072
c74 31 VSS 0.00381214f $X=0.126 $Y=0.072
c75 29 VSS 1.65557e-19 $X=0.081 $Y=0.1205
c76 28 VSS 9.91953e-19 $X=0.081 $Y=0.106
c77 26 VSS 4.0436e-19 $X=0.081 $Y=0.135
c78 22 VSS 0.00259367f $X=0.484 $Y=0.2025
c79 17 VSS 2.55988e-19 $X=0.484 $Y=0.0675
c80 9 VSS 5.38922e-19 $X=0.287 $Y=0.0675
c81 5 VSS 0.00237091f $X=0.081 $Y=0.135
c82 2 VSS 0.0648622f $X=0.081 $Y=0.0675
r83 72 73 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.5085 $Y2=0.234
r84 71 73 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.234 $X2=0.5085 $Y2=0.234
r85 68 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.504 $Y2=0.234
r86 65 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.513 $Y2=0.207
r87 64 65 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.164 $X2=0.513 $Y2=0.189
r88 63 64 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.07 $X2=0.513 $Y2=0.164
r89 62 71 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.234
r90 62 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.207
r91 61 63 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.07
r92 59 60 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.471
+ $Y=0.036 $X2=0.4785 $Y2=0.036
r93 58 59 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.471 $Y2=0.036
r94 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r95 56 57 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.036 $X2=0.45 $Y2=0.036
r96 55 56 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.447 $Y2=0.036
r97 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r98 53 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.396 $Y2=0.036
r99 52 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r100 51 52 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.308
+ $Y=0.036 $X2=0.342 $Y2=0.036
r101 50 51 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.308 $Y2=0.036
r102 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r103 47 60 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.4785 $Y2=0.036
r104 47 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036
+ $X2=0.486 $Y2=0.036
r105 44 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.261 $Y2=0.036
r106 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r107 42 43 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.234 $Y2=0.036
r108 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r109 40 41 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.146
+ $Y=0.036 $X2=0.18 $Y2=0.036
r110 38 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.288 $Y2=0.036
r111 38 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.261 $Y2=0.036
r112 38 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r113 36 40 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.146 $Y2=0.036
r114 35 61 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.036 $X2=0.513 $Y2=0.045
r115 35 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.486 $Y2=0.036
r116 33 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.045 $X2=0.144 $Y2=0.036
r117 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.063
r118 31 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.063
r119 31 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.09 $Y2=0.072
r120 28 29 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.106 $X2=0.081 $Y2=0.1205
r121 26 29 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1205
r122 24 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.081 $X2=0.09 $Y2=0.072
r123 24 28 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.081 $X2=0.081 $Y2=0.106
r124 22 68 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234
+ $X2=0.486 $Y2=0.234
r125 19 22 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.484 $Y2=0.2025
r126 17 48 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.486 $Y=0.0675 $X2=0.486 $Y2=0.036
r127 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.484 $Y2=0.0675
r128 13 39 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r129 10 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r130 9 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r131 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r132 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r133 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO331X1_ASAP7_75T_L%A3 2 5 7 10 13 VSS
c10 13 VSS 0.00221897f $X=0.135 $Y=0.135
c11 10 VSS 2.57666e-19 $X=0.135 $Y=0.115
c12 5 VSS 0.00122791f $X=0.135 $Y=0.135
c13 2 VSS 0.0596882f $X=0.135 $Y=0.0675
r14 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.115 $X2=0.135 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO331X1_ASAP7_75T_L%A2 2 5 7 10 VSS
c16 10 VSS 0.00193643f $X=0.189 $Y=0.115
c17 5 VSS 0.00110916f $X=0.189 $Y=0.135
c18 2 VSS 0.059482f $X=0.189 $Y=0.0675
r19 10 15 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r20 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r21 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO331X1_ASAP7_75T_L%A1 2 5 7 10 13 VSS
c16 13 VSS 0.00115482f $X=0.243 $Y=0.135
c17 10 VSS 3.80937e-19 $X=0.243 $Y=0.115
c18 5 VSS 0.00110907f $X=0.243 $Y=0.135
c19 2 VSS 0.060543f $X=0.243 $Y=0.0675
r20 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.115 $X2=0.243 $Y2=0.135
r21 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO331X1_ASAP7_75T_L%B1 2 5 7 10 VSS
c13 10 VSS 5.08499e-19 $X=0.297 $Y=0.116
c14 5 VSS 0.00110017f $X=0.297 $Y=0.135
c15 2 VSS 0.0616432f $X=0.297 $Y=0.0675
r16 10 13 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.116 $X2=0.297 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO331X1_ASAP7_75T_L%B2 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.35 $Y=0.115
c14 5 VSS 0.00112057f $X=0.351 $Y=0.135
c15 2 VSS 0.0616432f $X=0.351 $Y=0.0675
r16 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.115 $X2=0.351 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AO331X1_ASAP7_75T_L%B3 2 5 7 10 VSS
c11 10 VSS 6.93937e-19 $X=0.403 $Y=0.115
c12 5 VSS 0.00114932f $X=0.405 $Y=0.135
c13 2 VSS 0.0619365f $X=0.405 $Y=0.0675
r14 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.115 $X2=0.405 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO331X1_ASAP7_75T_L%C 2 5 7 10 VSS
c8 10 VSS 0.00201948f $X=0.457 $Y=0.115
c9 5 VSS 0.00178699f $X=0.459 $Y=0.135
c10 2 VSS 0.0660367f $X=0.459 $Y=0.0675
r11 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.115 $X2=0.459 $Y2=0.135
r12 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AO331X1_ASAP7_75T_L%Y 1 6 9 14 16 18 23 24 31 VSS
c9 34 VSS 9.17717e-19 $X=0.045 $Y=0.234
c10 33 VSS 0.0032947f $X=0.036 $Y=0.234
c11 31 VSS 0.00327598f $X=0.054 $Y=0.234
c12 24 VSS 0.00651756f $X=0.054 $Y=0.036
c13 23 VSS 0.0053018f $X=0.054 $Y=0.036
c14 21 VSS 0.0033063f $X=0.036 $Y=0.036
c15 20 VSS 2.98008e-19 $X=0.027 $Y=0.216
c16 19 VSS 2.15228e-19 $X=0.027 $Y=0.207
c17 18 VSS 0.00217784f $X=0.027 $Y=0.2
c18 16 VSS 0.00169414f $X=0.027 $Y=0.10525
c19 15 VSS 7.23378e-19 $X=0.027 $Y=0.063
c20 14 VSS 0.00209763f $X=0.03 $Y=0.1475
c21 12 VSS 2.81452e-19 $X=0.027 $Y=0.225
c22 9 VSS 0.00636217f $X=0.056 $Y=0.2025
c23 6 VSS 3.7894e-19 $X=0.071 $Y=0.2025
c24 1 VSS 3.3212e-19 $X=0.071 $Y=0.0675
r25 33 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.045 $Y2=0.234
r26 31 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.045 $Y2=0.234
r27 28 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.036 $Y2=0.234
r28 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r29 21 23 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.054 $Y2=0.036
r30 19 20 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.207 $X2=0.027 $Y2=0.216
r31 18 19 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.2 $X2=0.027 $Y2=0.207
r32 17 18 3.25926 $w=1.8e-08 $l=4.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.152 $X2=0.027 $Y2=0.2
r33 15 16 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.063 $X2=0.027 $Y2=0.10525
r34 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.1475 $X2=0.027 $Y2=0.152
r35 14 16 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.1475 $X2=0.027 $Y2=0.10525
r36 12 28 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.234
r37 12 20 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.216
r38 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r39 11 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.063
r40 9 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r41 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
r42 4 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r43 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./AO331x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO331x1_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C Y
* 
* Y	Y
* C	C
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 VSS N_3_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 noxref_14 N_A3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_15 N_A2_M2_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_3_M3_d N_A1_M3_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_16 N_B1_M4_g N_3_M4_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_17 N_B2_M5_g noxref_16 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 VSS N_B3_M6_g noxref_17 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_3_M7_d N_C_M7_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 VDD N_3_M8_g N_Y_M8_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M9 noxref_12 N_A3_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M10 VDD N_A2_M10_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M11 noxref_12 N_A1_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M12 noxref_13 N_B1_M12_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M13 noxref_12 N_B2_M13_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M14 noxref_13 N_B3_M14_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M15 N_3_M15_d N_C_M15_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "AO331x1_ASAP7_75t_L.pex.sp.AO331X1_ASAP7_75T_L.pxi"
* BEGIN of "./AO331x1_ASAP7_75t_L.pex.sp.AO331X1_ASAP7_75T_L.pxi"
* File: AO331x1_ASAP7_75t_L.pex.sp.AO331X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:06:56 2017
* 
x_PM_AO331X1_ASAP7_75T_L%3 N_3_M0_g N_3_c_2_p N_3_M8_g N_3_M4_s N_3_M3_d
+ N_3_M7_d N_3_M15_d N_3_c_31_p N_3_c_7_p N_3_c_3_p N_3_c_4_p N_3_c_25_p
+ N_3_c_28_p N_3_c_11_p N_3_c_40_p N_3_c_6_p N_3_c_41_p N_3_c_10_p N_3_c_21_p
+ N_3_c_13_p N_3_c_37_p N_3_c_16_p N_3_c_38_p N_3_c_18_p N_3_c_39_p N_3_c_20_p
+ N_3_c_23_p N_3_c_36_p N_3_c_32_p VSS PM_AO331X1_ASAP7_75T_L%3
x_PM_AO331X1_ASAP7_75T_L%A3 N_A3_M1_g N_A3_c_45_n N_A3_M9_g A3 N_A3_c_52_p VSS
+ PM_AO331X1_ASAP7_75T_L%A3
x_PM_AO331X1_ASAP7_75T_L%A2 N_A2_M2_g N_A2_c_60_n N_A2_M10_g A2 VSS
+ PM_AO331X1_ASAP7_75T_L%A2
x_PM_AO331X1_ASAP7_75T_L%A1 N_A1_M3_g N_A1_c_75_n N_A1_M11_g A1 N_A1_c_77_n VSS
+ PM_AO331X1_ASAP7_75T_L%A1
x_PM_AO331X1_ASAP7_75T_L%B1 N_B1_M4_g N_B1_c_91_n N_B1_M12_g B1 VSS
+ PM_AO331X1_ASAP7_75T_L%B1
x_PM_AO331X1_ASAP7_75T_L%B2 N_B2_M5_g N_B2_c_103_n N_B2_M13_g B2 VSS
+ PM_AO331X1_ASAP7_75T_L%B2
x_PM_AO331X1_ASAP7_75T_L%B3 N_B3_M6_g N_B3_c_116_n N_B3_M14_g B3 VSS
+ PM_AO331X1_ASAP7_75T_L%B3
x_PM_AO331X1_ASAP7_75T_L%C N_C_M7_g N_C_c_129_n N_C_M15_g C VSS
+ PM_AO331X1_ASAP7_75T_L%C
x_PM_AO331X1_ASAP7_75T_L%Y N_Y_M0_s N_Y_M8_s N_Y_c_138_p Y N_Y_c_132_n
+ N_Y_c_137_n N_Y_c_133_n N_Y_c_136_n N_Y_c_139_p VSS PM_AO331X1_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M1_g 0.00284417f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_3_c_2_p N_A3_c_45_n 9.34529e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_3_c_3_p A3 0.00200929f $X=0.081 $Y=0.1205 $X2=0.135 $Y2=0.115
cc_4 N_3_c_4_p A3 0.00133324f $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.115
cc_5 N_3_M0_g N_A2_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 N_3_c_6_p N_A2_M2_g 3.38929e-19 $X=0.198 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_7 N_3_c_7_p A2 2.69033e-19 $X=0.081 $Y=0.106 $X2=0.135 $Y2=0.115
cc_8 N_3_c_4_p A2 7.10035e-19 $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.115
cc_9 N_3_c_6_p A2 0.00123604f $X=0.198 $Y=0.036 $X2=0.135 $Y2=0.115
cc_10 N_3_c_10_p N_A1_M3_g 2.56935e-19 $X=0.252 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_11 N_3_c_11_p A1 0.0013295f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.115
cc_12 N_3_c_10_p A1 0.00123604f $X=0.252 $Y=0.036 $X2=0.135 $Y2=0.115
cc_13 N_3_c_13_p N_B1_M4_g 2.64276e-19 $X=0.306 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_14 N_3_c_11_p B1 0.0013295f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.115
cc_15 N_3_c_13_p B1 0.00124805f $X=0.306 $Y=0.036 $X2=0.135 $Y2=0.115
cc_16 N_3_c_16_p N_B2_M5_g 3.38929e-19 $X=0.36 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_17 N_3_c_16_p B2 0.00123064f $X=0.36 $Y=0.036 $X2=0.135 $Y2=0.115
cc_18 N_3_c_18_p N_B3_M6_g 2.56935e-19 $X=0.414 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_19 N_3_c_18_p B3 0.00123064f $X=0.414 $Y=0.036 $X2=0.135 $Y2=0.115
cc_20 N_3_c_20_p N_C_M7_g 2.64276e-19 $X=0.468 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_21 N_3_c_21_p C 0.00114532f $X=0.486 $Y=0.036 $X2=0.135 $Y2=0.115
cc_22 N_3_c_20_p C 0.00124805f $X=0.468 $Y=0.036 $X2=0.135 $Y2=0.115
cc_23 N_3_c_23_p C 0.00392202f $X=0.513 $Y=0.164 $X2=0.135 $Y2=0.115
cc_24 N_3_c_3_p Y 0.00179201f $X=0.081 $Y=0.1205 $X2=0.135 $Y2=0.135
cc_25 N_3_c_25_p N_Y_c_132_n 0.00179201f $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_26 N_3_M0_g N_Y_c_133_n 2.49235e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_3_c_25_p N_Y_c_133_n 8.16832e-19 $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_28 N_3_c_28_p N_Y_c_133_n 4.96595e-19 $X=0.144 $Y=0.036 $X2=0 $Y2=0
cc_29 N_3_c_25_p N_Y_c_136_n 0.00135457f $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_30 VSS N_3_c_11_p 0.00107252f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.115
cc_31 VSS N_3_c_31_p 2.24644e-19 $X=0.484 $Y=0.2025 $X2=0 $Y2=0
cc_32 VSS N_3_c_32_p 2.83845e-19 $X=0.504 $Y=0.234 $X2=0 $Y2=0
cc_33 VSS N_3_c_31_p 0.0036142f $X=0.484 $Y=0.2025 $X2=0.135 $Y2=0.115
cc_34 VSS N_3_c_32_p 4.47506e-19 $X=0.504 $Y=0.234 $X2=0.135 $Y2=0.115
cc_35 VSS N_3_c_31_p 3.99913e-19 $X=0.484 $Y=0.2025 $X2=0 $Y2=0
cc_36 VSS N_3_c_36_p 3.53514e-19 $X=0.513 $Y=0.207 $X2=0 $Y2=0
cc_37 VSS N_3_c_37_p 3.03225e-19 $X=0.342 $Y=0.036 $X2=0 $Y2=0
cc_38 VSS N_3_c_38_p 3.03225e-19 $X=0.396 $Y=0.036 $X2=0 $Y2=0
cc_39 VSS N_3_c_39_p 3.03225e-19 $X=0.447 $Y=0.036 $X2=0 $Y2=0
cc_40 VSS N_3_c_40_p 3.56327e-19 $X=0.18 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_41 VSS N_3_c_41_p 3.56327e-19 $X=0.234 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_42 VSS N_3_c_37_p 3.48201e-19 $X=0.342 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_43 VSS N_3_c_38_p 3.34078e-19 $X=0.396 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_44 N_A3_M1_g N_A2_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_45 N_A3_c_45_n N_A2_c_60_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_46 A3 A2 0.00393501f $X=0.135 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_47 N_A3_M1_g N_A1_M3_g 2.66145e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_48 N_A3_c_52_p N_Y_c_137_n 4.90507e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_49 VSS N_A3_c_52_p 0.00114532f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_50 N_A2_M2_g N_A1_M3_g 0.00327995f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_51 N_A2_c_60_n N_A1_c_75_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_52 A2 A1 0.00193488f $X=0.189 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_53 A2 N_A1_c_77_n 0.00386975f $X=0.189 $Y=0.115 $X2=0.27 $Y2=0.0675
cc_54 N_A2_M2_g N_B1_M4_g 2.71887e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_55 VSS A2 0.00114532f $X=0.189 $Y=0.115 $X2=0.081 $Y2=0.135
cc_56 VSS N_A2_M2_g 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.081
cc_57 VSS A2 0.00125352f $X=0.189 $Y=0.115 $X2=0.081 $Y2=0.081
cc_58 N_A1_M3_g N_B1_M4_g 0.0036939f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_59 N_A1_c_75_n N_B1_c_91_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_60 A1 B1 0.00389755f $X=0.243 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_61 N_A1_M3_g N_B2_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_62 VSS A1 8.72546e-19 $X=0.243 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_63 VSS N_A1_M3_g 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_64 VSS N_A1_c_77_n 0.00125352f $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_65 VSS N_A1_c_77_n 2.75021e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_66 N_B1_M4_g N_B2_M5_g 0.00371573f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_67 N_B1_c_91_n N_B2_c_103_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_68 B1 B2 0.00483372f $X=0.297 $Y=0.116 $X2=0.253 $Y2=0.0675
cc_69 N_B1_M4_g N_B3_M6_g 3.06651e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_70 VSS N_B1_M4_g 3.57119e-19 $X=0.297 $Y=0.0675 $X2=0.126 $Y2=0.072
cc_71 VSS B1 5.37372e-19 $X=0.297 $Y=0.116 $X2=0.126 $Y2=0.072
cc_72 N_B2_M5_g N_B3_M6_g 0.0036939f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_73 N_B2_c_103_n N_B3_c_116_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_74 B2 B3 0.00483372f $X=0.35 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_75 N_B2_M5_g N_C_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_76 VSS N_B2_M5_g 2.21754e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.106
cc_77 VSS N_B2_M5_g 2.76185e-19 $X=0.351 $Y=0.0675 $X2=0.469 $Y2=0.2025
cc_78 VSS B2 0.0012322f $X=0.35 $Y=0.115 $X2=0.469 $Y2=0.2025
cc_79 N_B3_M6_g N_C_M7_g 0.00333077f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_80 N_B3_c_116_n N_C_c_129_n 9.33263e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_81 B3 C 0.00406322f $X=0.403 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_82 VSS N_B3_M6_g 3.51973e-19 $X=0.405 $Y=0.0675 $X2=0.484 $Y2=0.2025
cc_83 VSS B3 0.00121543f $X=0.403 $Y=0.115 $X2=0.484 $Y2=0.2025
cc_84 VSS N_Y_c_138_p 2.87474e-19 $X=0.056 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_85 VSS N_Y_c_139_p 2.83353e-19 $X=0.054 $Y=0.234 $X2=0 $Y2=0

* END of "./AO331x1_ASAP7_75t_L.pex.sp.AO331X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO331x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:07:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO331x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO331x2_ASAP7_75t_L.pex.sp.pex"
* File: AO331x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:07:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO331X2_ASAP7_75T_L%3 2 7 10 13 15 17 18 22 27 30 36 37 39 40 44 47
+ 49 50 51 52 56 58 60 61 62 63 64 66 72 74 80 VSS
c52 80 VSS 0.00385307f $X=0.558 $Y=0.234
c53 79 VSS 0.00278591f $X=0.567 $Y=0.234
c54 74 VSS 6.85875e-19 $X=0.567 $Y=0.207
c55 73 VSS 0.00104083f $X=0.567 $Y=0.189
c56 72 VSS 0.00414953f $X=0.567 $Y=0.164
c57 71 VSS 8.11244e-19 $X=0.567 $Y=0.07
c58 70 VSS 0.00102822f $X=0.567 $Y=0.225
c59 68 VSS 6.9735e-19 $X=0.5325 $Y=0.036
c60 67 VSS 2.39163e-19 $X=0.525 $Y=0.036
c61 66 VSS 0.00146362f $X=0.522 $Y=0.036
c62 65 VSS 2.39163e-19 $X=0.504 $Y=0.036
c63 64 VSS 0.00606761f $X=0.501 $Y=0.036
c64 63 VSS 0.00142296f $X=0.468 $Y=0.036
c65 62 VSS 0.00343941f $X=0.45 $Y=0.036
c66 61 VSS 0.00142296f $X=0.414 $Y=0.036
c67 60 VSS 0.00325376f $X=0.396 $Y=0.036
c68 59 VSS 1.47784e-19 $X=0.362 $Y=0.036
c69 58 VSS 0.00146362f $X=0.36 $Y=0.036
c70 57 VSS 0.00274887f $X=0.342 $Y=0.036
c71 56 VSS 0.00676142f $X=0.54 $Y=0.036
c72 53 VSS 0.00106181f $X=0.315 $Y=0.036
c73 52 VSS 0.00142296f $X=0.306 $Y=0.036
c74 51 VSS 0.0037673f $X=0.288 $Y=0.036
c75 50 VSS 0.00142296f $X=0.252 $Y=0.036
c76 49 VSS 0.00347922f $X=0.234 $Y=0.036
c77 48 VSS 1.51923e-19 $X=0.2 $Y=0.036
c78 47 VSS 0.00218387f $X=0.324 $Y=0.036
c79 44 VSS 0.00238538f $X=0.198 $Y=0.036
c80 43 VSS 0.00596382f $X=0.558 $Y=0.036
c81 42 VSS 9.0336e-19 $X=0.189 $Y=0.063
c82 40 VSS 3.49137e-19 $X=0.144 $Y=0.072
c83 39 VSS 0.00381214f $X=0.18 $Y=0.072
c84 37 VSS 1.33309e-19 $X=0.135 $Y=0.1205
c85 36 VSS 9.91953e-19 $X=0.135 $Y=0.106
c86 34 VSS 4.03627e-19 $X=0.135 $Y=0.135
c87 30 VSS 0.00259367f $X=0.538 $Y=0.2025
c88 25 VSS 2.55988e-19 $X=0.538 $Y=0.0675
c89 17 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c90 13 VSS 0.00426847f $X=0.135 $Y=0.135
c91 10 VSS 0.0608921f $X=0.135 $Y=0.0675
c92 2 VSS 0.0639847f $X=0.081 $Y=0.0675
r93 80 81 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.5625 $Y2=0.234
r94 79 81 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.234 $X2=0.5625 $Y2=0.234
r95 76 80 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.558 $Y2=0.234
r96 73 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.567 $Y2=0.207
r97 72 73 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.164 $X2=0.567 $Y2=0.189
r98 71 72 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.07 $X2=0.567 $Y2=0.164
r99 70 79 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.225 $X2=0.567 $Y2=0.234
r100 70 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.225 $X2=0.567 $Y2=0.207
r101 69 71 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.045 $X2=0.567 $Y2=0.07
r102 67 68 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.525
+ $Y=0.036 $X2=0.5325 $Y2=0.036
r103 66 67 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.525 $Y2=0.036
r104 65 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.522 $Y2=0.036
r105 64 65 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.501
+ $Y=0.036 $X2=0.504 $Y2=0.036
r106 63 64 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.501 $Y2=0.036
r107 62 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r108 61 62 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.45 $Y2=0.036
r109 60 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r110 59 60 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.362
+ $Y=0.036 $X2=0.396 $Y2=0.036
r111 58 59 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.362 $Y2=0.036
r112 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r113 55 68 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.5325 $Y2=0.036
r114 55 56 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r115 52 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.315 $Y2=0.036
r116 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r117 50 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r118 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r119 48 49 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2
+ $Y=0.036 $X2=0.234 $Y2=0.036
r120 46 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r121 46 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.315 $Y2=0.036
r122 46 47 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r123 44 48 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.2 $Y2=0.036
r124 43 69 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.036 $X2=0.567 $Y2=0.045
r125 43 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.54 $Y2=0.036
r126 41 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.045 $X2=0.198 $Y2=0.036
r127 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r128 39 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.072 $X2=0.189 $Y2=0.063
r129 39 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.072 $X2=0.144 $Y2=0.072
r130 36 37 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.106 $X2=0.135 $Y2=0.1205
r131 34 37 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.1205
r132 32 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.081 $X2=0.144 $Y2=0.072
r133 32 36 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.081 $X2=0.135 $Y2=0.106
r134 30 76 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r135 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.538 $Y2=0.2025
r136 25 56 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r137 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.538 $Y2=0.0675
r138 21 47 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r139 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r140 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r141 13 34 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r142 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r143 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r144 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r145 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r146 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO331X2_ASAP7_75T_L%A3 2 5 7 10 13 VSS
c11 13 VSS 0.0023342f $X=0.189 $Y=0.135
c12 10 VSS 3.21887e-19 $X=0.189 $Y=0.115
c13 5 VSS 0.0011078f $X=0.189 $Y=0.135
c14 2 VSS 0.0588951f $X=0.189 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO331X2_ASAP7_75T_L%A2 2 5 7 10 VSS
c16 10 VSS 0.00193643f $X=0.243 $Y=0.115
c17 5 VSS 0.0011122f $X=0.243 $Y=0.135
c18 2 VSS 0.059482f $X=0.243 $Y=0.0675
r19 10 15 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.115 $X2=0.243 $Y2=0.135
r20 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r21 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO331X2_ASAP7_75T_L%A1 2 5 7 10 13 VSS
c16 13 VSS 0.00115482f $X=0.297 $Y=0.135
c17 10 VSS 3.80937e-19 $X=0.297 $Y=0.115
c18 5 VSS 0.00110907f $X=0.297 $Y=0.135
c19 2 VSS 0.060543f $X=0.297 $Y=0.0675
r20 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.115 $X2=0.297 $Y2=0.135
r21 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO331X2_ASAP7_75T_L%B1 2 5 7 10 VSS
c13 10 VSS 5.08499e-19 $X=0.351 $Y=0.116
c14 5 VSS 0.00110017f $X=0.351 $Y=0.135
c15 2 VSS 0.0616432f $X=0.351 $Y=0.0675
r16 10 13 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.116 $X2=0.351 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AO331X2_ASAP7_75T_L%B2 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.404 $Y=0.115
c14 5 VSS 0.00112057f $X=0.405 $Y=0.135
c15 2 VSS 0.0616432f $X=0.405 $Y=0.0675
r16 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.115 $X2=0.405 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO331X2_ASAP7_75T_L%B3 2 5 7 10 VSS
c11 10 VSS 6.93937e-19 $X=0.457 $Y=0.115
c12 5 VSS 0.00114932f $X=0.459 $Y=0.135
c13 2 VSS 0.0619365f $X=0.459 $Y=0.0675
r14 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.115 $X2=0.459 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AO331X2_ASAP7_75T_L%C 2 5 7 10 VSS
c8 10 VSS 0.00201948f $X=0.511 $Y=0.115
c9 5 VSS 0.00178699f $X=0.513 $Y=0.135
c10 2 VSS 0.0660367f $X=0.513 $Y=0.0675
r11 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.115 $X2=0.513 $Y2=0.135
r12 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AO331X2_ASAP7_75T_L%Y 1 2 6 7 10 14 16 23 24 30 VSS
c17 30 VSS 0.00681666f $X=0.108 $Y=0.234
c18 28 VSS 0.00385179f $X=0.063 $Y=0.234
c19 24 VSS 0.0102944f $X=0.108 $Y=0.036
c20 23 VSS 0.00783831f $X=0.108 $Y=0.036
c21 21 VSS 0.00386107f $X=0.063 $Y=0.036
c22 20 VSS 8.50351e-19 $X=0.054 $Y=0.216
c23 19 VSS 4.97402e-19 $X=0.054 $Y=0.207
c24 18 VSS 0.00434529f $X=0.054 $Y=0.2
c25 16 VSS 0.00372228f $X=0.054 $Y=0.10525
c26 15 VSS 0.00165346f $X=0.054 $Y=0.063
c27 14 VSS 0.00242602f $X=0.057 $Y=0.1475
c28 12 VSS 8.0311e-19 $X=0.054 $Y=0.225
c29 10 VSS 0.00894851f $X=0.108 $Y=0.2025
c30 6 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c31 1 VSS 5.25448e-19 $X=0.125 $Y=0.0675
r32 28 30 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.234 $X2=0.108 $Y2=0.234
r33 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r34 21 23 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.036 $X2=0.108 $Y2=0.036
r35 19 20 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.207 $X2=0.054 $Y2=0.216
r36 18 19 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.2 $X2=0.054 $Y2=0.207
r37 17 18 3.25926 $w=1.8e-08 $l=4.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.152 $X2=0.054 $Y2=0.2
r38 15 16 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.063 $X2=0.054 $Y2=0.10525
r39 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.1475 $X2=0.054 $Y2=0.152
r40 14 16 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.1475 $X2=0.054 $Y2=0.10525
r41 12 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.054 $Y=0.225 $X2=0.063 $Y2=0.234
r42 12 20 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.225 $X2=0.054 $Y2=0.216
r43 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.054 $Y=0.045 $X2=0.063 $Y2=0.036
r44 11 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.045 $X2=0.054 $Y2=0.063
r45 10 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r46 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r47 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r48 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r49 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r50 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./AO331x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO331x2_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C Y
* 
* Y	Y
* C	C
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_14 N_A3_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_15 N_A2_M3_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_3_M4_d N_A1_M4_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_16 N_B1_M5_g N_3_M5_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_17 N_B2_M6_g noxref_16 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 VSS N_B3_M7_g noxref_17 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_3_M8_d N_C_M8_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_3_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M10 N_Y_M10_d N_3_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M11 noxref_12 N_A3_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M12 VDD N_A2_M12_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M13 noxref_12 N_A1_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M14 noxref_13 N_B1_M14_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M15 noxref_12 N_B2_M15_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M16 noxref_13 N_B3_M16_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M17 N_3_M17_d N_C_M17_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
*
* 
* .include "AO331x2_ASAP7_75t_L.pex.sp.AO331X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO331x2_ASAP7_75t_L.pex.sp.AO331X2_ASAP7_75T_L.pxi"
* File: AO331x2_ASAP7_75t_L.pex.sp.AO331X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:07:18 2017
* 
x_PM_AO331X2_ASAP7_75T_L%3 N_3_M0_g N_3_M9_g N_3_M1_g N_3_c_3_p N_3_M10_g
+ N_3_M5_s N_3_M4_d N_3_M8_d N_3_M17_d N_3_c_40_p N_3_c_8_p N_3_c_4_p N_3_c_5_p
+ N_3_c_29_p N_3_c_34_p N_3_c_12_p N_3_c_49_p N_3_c_7_p N_3_c_50_p N_3_c_11_p
+ N_3_c_22_p N_3_c_14_p N_3_c_46_p N_3_c_17_p N_3_c_47_p N_3_c_19_p N_3_c_48_p
+ N_3_c_21_p N_3_c_24_p N_3_c_45_p N_3_c_41_p VSS PM_AO331X2_ASAP7_75T_L%3
x_PM_AO331X2_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_55_n N_A3_M11_g A3 N_A3_c_62_p VSS
+ PM_AO331X2_ASAP7_75T_L%A3
x_PM_AO331X2_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_70_n N_A2_M12_g A2 VSS
+ PM_AO331X2_ASAP7_75T_L%A2
x_PM_AO331X2_ASAP7_75T_L%A1 N_A1_M4_g N_A1_c_85_n N_A1_M13_g A1 N_A1_c_87_n VSS
+ PM_AO331X2_ASAP7_75T_L%A1
x_PM_AO331X2_ASAP7_75T_L%B1 N_B1_M5_g N_B1_c_101_n N_B1_M14_g B1 VSS
+ PM_AO331X2_ASAP7_75T_L%B1
x_PM_AO331X2_ASAP7_75T_L%B2 N_B2_M6_g N_B2_c_113_n N_B2_M15_g B2 VSS
+ PM_AO331X2_ASAP7_75T_L%B2
x_PM_AO331X2_ASAP7_75T_L%B3 N_B3_M7_g N_B3_c_126_n N_B3_M16_g B3 VSS
+ PM_AO331X2_ASAP7_75T_L%B3
x_PM_AO331X2_ASAP7_75T_L%C N_C_M8_g N_C_c_139_n N_C_M17_g C VSS
+ PM_AO331X2_ASAP7_75T_L%C
x_PM_AO331X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_M10_d N_Y_M9_d N_Y_c_143_n Y
+ N_Y_c_145_n N_Y_c_146_n N_Y_c_151_n N_Y_c_153_n VSS PM_AO331X2_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_A3_M2_g 0.00284417f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_A3_c_55_n 9.59383e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_4 N_3_c_4_p A3 0.0020116f $X=0.135 $Y=0.1205 $X2=0.189 $Y2=0.115
cc_5 N_3_c_5_p A3 0.00133324f $X=0.18 $Y=0.072 $X2=0.189 $Y2=0.115
cc_6 N_3_M1_g N_A2_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_7 N_3_c_7_p N_A2_M3_g 3.38929e-19 $X=0.252 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_8 N_3_c_8_p A2 2.69033e-19 $X=0.135 $Y=0.106 $X2=0.189 $Y2=0.115
cc_9 N_3_c_5_p A2 7.10035e-19 $X=0.18 $Y=0.072 $X2=0.189 $Y2=0.115
cc_10 N_3_c_7_p A2 0.00123604f $X=0.252 $Y=0.036 $X2=0.189 $Y2=0.115
cc_11 N_3_c_11_p N_A1_M4_g 2.56935e-19 $X=0.306 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_12 N_3_c_12_p A1 0.0013295f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.115
cc_13 N_3_c_11_p A1 0.00123604f $X=0.306 $Y=0.036 $X2=0.189 $Y2=0.115
cc_14 N_3_c_14_p N_B1_M5_g 2.64276e-19 $X=0.36 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_15 N_3_c_12_p B1 0.0013295f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.115
cc_16 N_3_c_14_p B1 0.00124805f $X=0.36 $Y=0.036 $X2=0.189 $Y2=0.115
cc_17 N_3_c_17_p N_B2_M6_g 3.38929e-19 $X=0.414 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_18 N_3_c_17_p B2 0.00123064f $X=0.414 $Y=0.036 $X2=0.189 $Y2=0.115
cc_19 N_3_c_19_p N_B3_M7_g 2.56935e-19 $X=0.468 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_20 N_3_c_19_p B3 0.00123064f $X=0.468 $Y=0.036 $X2=0.189 $Y2=0.115
cc_21 N_3_c_21_p N_C_M8_g 2.64276e-19 $X=0.522 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_22 N_3_c_22_p C 0.00114532f $X=0.54 $Y=0.036 $X2=0.189 $Y2=0.115
cc_23 N_3_c_21_p C 0.00124805f $X=0.522 $Y=0.036 $X2=0.189 $Y2=0.115
cc_24 N_3_c_24_p C 0.00392202f $X=0.567 $Y=0.164 $X2=0.189 $Y2=0.115
cc_25 N_3_c_3_p N_Y_M1_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_26 N_3_c_3_p N_Y_M10_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_27 N_3_c_3_p N_Y_c_143_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.115
cc_28 N_3_c_4_p Y 9.40908e-19 $X=0.135 $Y=0.1205 $X2=0.189 $Y2=0.135
cc_29 N_3_c_29_p N_Y_c_145_n 9.40908e-19 $X=0.144 $Y=0.072 $X2=0 $Y2=0
cc_30 N_3_M0_g N_Y_c_146_n 4.59284e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_3_M1_g N_Y_c_146_n 2.51294e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_32 N_3_c_3_p N_Y_c_146_n 6.10804e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_33 N_3_c_29_p N_Y_c_146_n 8.16832e-19 $X=0.144 $Y=0.072 $X2=0 $Y2=0
cc_34 N_3_c_34_p N_Y_c_146_n 5.0963e-19 $X=0.198 $Y=0.036 $X2=0 $Y2=0
cc_35 N_3_c_3_p N_Y_c_151_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_36 N_3_c_29_p N_Y_c_151_n 0.00152998f $X=0.144 $Y=0.072 $X2=0 $Y2=0
cc_37 N_3_M0_g N_Y_c_153_n 4.59284e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_38 N_3_c_3_p N_Y_c_153_n 5.51214e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_39 VSS N_3_c_12_p 0.00107252f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.115
cc_40 VSS N_3_c_40_p 2.24644e-19 $X=0.538 $Y=0.2025 $X2=0 $Y2=0
cc_41 VSS N_3_c_41_p 2.83845e-19 $X=0.558 $Y=0.234 $X2=0 $Y2=0
cc_42 VSS N_3_c_40_p 0.0036142f $X=0.538 $Y=0.2025 $X2=0.189 $Y2=0.115
cc_43 VSS N_3_c_41_p 4.47506e-19 $X=0.558 $Y=0.234 $X2=0.189 $Y2=0.115
cc_44 VSS N_3_c_40_p 3.99913e-19 $X=0.538 $Y=0.2025 $X2=0 $Y2=0
cc_45 VSS N_3_c_45_p 3.53514e-19 $X=0.567 $Y=0.207 $X2=0 $Y2=0
cc_46 VSS N_3_c_46_p 3.03225e-19 $X=0.396 $Y=0.036 $X2=0 $Y2=0
cc_47 VSS N_3_c_47_p 3.03225e-19 $X=0.45 $Y=0.036 $X2=0 $Y2=0
cc_48 VSS N_3_c_48_p 3.03225e-19 $X=0.501 $Y=0.036 $X2=0 $Y2=0
cc_49 VSS N_3_c_49_p 3.56327e-19 $X=0.234 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_50 VSS N_3_c_50_p 3.56327e-19 $X=0.288 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_51 VSS N_3_c_46_p 3.48201e-19 $X=0.396 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_52 VSS N_3_c_47_p 3.34078e-19 $X=0.45 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_53 N_A3_M2_g N_A2_M3_g 0.00344695f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_54 N_A3_c_55_n N_A2_c_70_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_55 A3 A2 0.00393501f $X=0.189 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_56 N_A3_M2_g N_A1_M4_g 2.66145e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_57 N_A3_c_62_p Y 4.07379e-19 $X=0.189 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_58 VSS N_A3_c_62_p 0.00114532f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_59 N_A2_M3_g N_A1_M4_g 0.00327995f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_60 N_A2_c_70_n N_A1_c_85_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_61 A2 A1 0.00193488f $X=0.243 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_62 A2 N_A1_c_87_n 0.00386975f $X=0.243 $Y=0.115 $X2=0.135 $Y2=0.135
cc_63 N_A2_M3_g N_B1_M5_g 2.71887e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_64 VSS A2 0.00114532f $X=0.243 $Y=0.115 $X2=0.081 $Y2=0.135
cc_65 VSS N_A2_M3_g 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_66 VSS A2 0.00125352f $X=0.243 $Y=0.115 $X2=0 $Y2=0
cc_67 N_A1_M4_g N_B1_M5_g 0.0036939f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_68 N_A1_c_85_n N_B1_c_101_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_69 A1 B1 0.00389755f $X=0.297 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_70 N_A1_M4_g N_B2_M6_g 3.06651e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_71 VSS A1 8.72546e-19 $X=0.297 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_72 VSS N_A1_M4_g 2.64276e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_73 VSS N_A1_c_87_n 0.00125352f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_74 VSS N_A1_c_87_n 2.75021e-19 $X=0.297 $Y=0.135 $X2=0.307 $Y2=0.0675
cc_75 N_B1_M5_g N_B2_M6_g 0.00371573f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_76 N_B1_c_101_n N_B2_c_113_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_77 B1 B2 0.00483372f $X=0.351 $Y=0.116 $X2=0.135 $Y2=0.0675
cc_78 N_B1_M5_g N_B3_M7_g 3.06651e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_79 VSS N_B1_M5_g 3.57119e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_80 VSS B1 5.37372e-19 $X=0.351 $Y=0.116 $X2=0 $Y2=0
cc_81 N_B2_M6_g N_B3_M7_g 0.0036939f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_82 N_B2_c_113_n N_B3_c_126_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_83 B2 B3 0.00483372f $X=0.404 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_84 N_B2_M6_g N_C_M8_g 2.71887e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_85 VSS N_B2_M6_g 2.21754e-19 $X=0.405 $Y=0.0675 $X2=0.538 $Y2=0.2025
cc_86 VSS N_B2_M6_g 2.76185e-19 $X=0.405 $Y=0.0675 $X2=0.324 $Y2=0.0675
cc_87 VSS B2 0.0012322f $X=0.404 $Y=0.115 $X2=0.324 $Y2=0.0675
cc_88 N_B3_M7_g N_C_M8_g 0.00333077f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_89 N_B3_c_126_n N_C_c_139_n 9.33263e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.135
cc_90 B3 C 0.00406322f $X=0.457 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_91 VSS N_B3_M7_g 3.51973e-19 $X=0.459 $Y=0.0675 $X2=0.523 $Y2=0.0675
cc_92 VSS B3 0.00121543f $X=0.457 $Y=0.115 $X2=0.523 $Y2=0.0675
cc_93 VSS N_Y_c_143_n 2.23372e-19 $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_94 VSS N_Y_c_153_n 2.92759e-19 $X=0.108 $Y=0.234 $X2=0.538 $Y2=0.0675

* END of "./AO331x2_ASAP7_75t_L.pex.sp.AO331X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO332x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:07:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO332x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO332x1_ASAP7_75t_L.pex.sp.pex"
* File: AO332x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:07:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO332X1_ASAP7_75T_L%3 2 5 7 9 10 14 19 20 23 28 29 31 32 38 41 43 44
+ 45 46 47 50 51 52 53 54 55 57 59 61 62 68 69 70 75 VSS
c55 75 VSS 0.00412141f $X=0.567 $Y=0.164
c56 74 VSS 9.6701e-19 $X=0.567 $Y=0.07
c57 73 VSS 0.00112176f $X=0.567 $Y=0.189
c58 71 VSS 4.93718e-20 $X=0.557 $Y=0.198
c59 70 VSS 4.1269e-19 $X=0.556 $Y=0.198
c60 69 VSS 8.46035e-21 $X=0.522 $Y=0.198
c61 68 VSS 4.70878e-19 $X=0.504 $Y=0.198
c62 63 VSS 0.0019286f $X=0.558 $Y=0.198
c63 62 VSS 0.00146362f $X=0.522 $Y=0.036
c64 61 VSS 0.00296425f $X=0.504 $Y=0.036
c65 60 VSS 3.35992e-19 $X=0.471 $Y=0.036
c66 59 VSS 0.00142296f $X=0.468 $Y=0.036
c67 58 VSS 0.00672869f $X=0.45 $Y=0.036
c68 57 VSS 0.00142296f $X=0.414 $Y=0.036
c69 56 VSS 3.35992e-19 $X=0.396 $Y=0.036
c70 55 VSS 0.00311761f $X=0.393 $Y=0.036
c71 54 VSS 0.00146362f $X=0.36 $Y=0.036
c72 53 VSS 0.00340162f $X=0.342 $Y=0.036
c73 52 VSS 0.00146362f $X=0.306 $Y=0.036
c74 51 VSS 0.00256536f $X=0.288 $Y=0.036
c75 50 VSS 0.00357414f $X=0.54 $Y=0.036
c76 47 VSS 8.84964e-19 $X=0.261 $Y=0.036
c77 46 VSS 0.00142296f $X=0.252 $Y=0.036
c78 45 VSS 0.00360252f $X=0.234 $Y=0.036
c79 44 VSS 0.00142296f $X=0.198 $Y=0.036
c80 43 VSS 0.00331443f $X=0.18 $Y=0.036
c81 42 VSS 1.51923e-19 $X=0.146 $Y=0.036
c82 41 VSS 0.00220219f $X=0.27 $Y=0.036
c83 38 VSS 0.00233672f $X=0.144 $Y=0.036
c84 37 VSS 0.00702647f $X=0.558 $Y=0.036
c85 36 VSS 9.0336e-19 $X=0.135 $Y=0.063
c86 34 VSS 0.00182969f $X=0.11 $Y=0.072
c87 33 VSS 8.41473e-20 $X=0.094 $Y=0.072
c88 32 VSS 4.67384e-20 $X=0.09 $Y=0.072
c89 31 VSS 0.00174552f $X=0.126 $Y=0.072
c90 29 VSS 1.71139e-19 $X=0.081 $Y=0.1205
c91 28 VSS 9.91953e-19 $X=0.081 $Y=0.106
c92 26 VSS 3.54713e-19 $X=0.081 $Y=0.135
c93 23 VSS 0.0023085f $X=0.486 $Y=0.2025
c94 19 VSS 5.70099e-19 $X=0.503 $Y=0.2025
c95 17 VSS 2.69461e-19 $X=0.538 $Y=0.0675
c96 9 VSS 5.38922e-19 $X=0.287 $Y=0.0675
c97 5 VSS 0.00176753f $X=0.081 $Y=0.135
c98 2 VSS 0.0645889f $X=0.081 $Y=0.0675
r99 74 75 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.07 $X2=0.567 $Y2=0.164
r100 73 75 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.567 $Y2=0.164
r101 72 74 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.045 $X2=0.567 $Y2=0.07
r102 70 71 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.556
+ $Y=0.198 $X2=0.557 $Y2=0.198
r103 69 70 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.198 $X2=0.556 $Y2=0.198
r104 68 69 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.198 $X2=0.522 $Y2=0.198
r105 65 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.198 $X2=0.504 $Y2=0.198
r106 63 73 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.198 $X2=0.567 $Y2=0.189
r107 63 71 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.198 $X2=0.557 $Y2=0.198
r108 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.522 $Y2=0.036
r109 60 61 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.471
+ $Y=0.036 $X2=0.504 $Y2=0.036
r110 59 60 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.471 $Y2=0.036
r111 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r112 57 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.45 $Y2=0.036
r113 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r114 55 56 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.393
+ $Y=0.036 $X2=0.396 $Y2=0.036
r115 54 55 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.393 $Y2=0.036
r116 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r117 52 53 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.342 $Y2=0.036
r118 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r119 49 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.522 $Y2=0.036
r120 49 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r121 46 47 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.261 $Y2=0.036
r122 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r123 44 45 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.234 $Y2=0.036
r124 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r125 42 43 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.146
+ $Y=0.036 $X2=0.18 $Y2=0.036
r126 40 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.288 $Y2=0.036
r127 40 47 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.261 $Y2=0.036
r128 40 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r129 38 42 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.146 $Y2=0.036
r130 37 72 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.036 $X2=0.567 $Y2=0.045
r131 37 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.54 $Y2=0.036
r132 35 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.045 $X2=0.144 $Y2=0.036
r133 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.063
r134 33 34 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.072 $X2=0.11 $Y2=0.072
r135 32 33 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.094 $Y2=0.072
r136 31 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.063
r137 31 34 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.11 $Y2=0.072
r138 28 29 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.106 $X2=0.081 $Y2=0.1205
r139 26 29 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1205
r140 24 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.081 $X2=0.09 $Y2=0.072
r141 24 28 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.081 $X2=0.081 $Y2=0.106
r142 23 65 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.198
+ $X2=0.486 $Y2=0.198
r143 20 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.486 $Y2=0.2025
r144 19 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.2025 $X2=0.486 $Y2=0.2025
r145 17 50 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r146 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.538 $Y2=0.0675
r147 13 41 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r148 10 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r149 9 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r150 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r151 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r152 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO332X1_ASAP7_75T_L%A3 2 5 7 10 13 VSS
c11 13 VSS 0.00226375f $X=0.135 $Y=0.135
c12 10 VSS 2.53832e-19 $X=0.135 $Y=0.115
c13 5 VSS 0.00122791f $X=0.135 $Y=0.135
c14 2 VSS 0.0596346f $X=0.135 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.115 $X2=0.135 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO332X1_ASAP7_75T_L%A2 2 5 7 10 15 VSS
c17 15 VSS 0.00159343f $X=0.189 $Y=0.135
c18 10 VSS 7.68637e-19 $X=0.189 $Y=0.115
c19 5 VSS 0.00110907f $X=0.189 $Y=0.135
c20 2 VSS 0.059482f $X=0.189 $Y=0.0675
r21 10 15 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r22 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r23 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r24 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO332X1_ASAP7_75T_L%A1 2 5 7 10 VSS
c12 10 VSS 4.82288e-19 $X=0.243 $Y=0.115
c13 5 VSS 0.00111383f $X=0.243 $Y=0.135
c14 2 VSS 0.0608471f $X=0.243 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.115 $X2=0.243 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO332X1_ASAP7_75T_L%B1 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.297 $Y=0.116
c14 5 VSS 0.00111336f $X=0.297 $Y=0.135
c15 2 VSS 0.0617786f $X=0.297 $Y=0.0675
r16 10 13 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.116 $X2=0.297 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO332X1_ASAP7_75T_L%B2 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.35 $Y=0.115
c14 5 VSS 0.00112198f $X=0.351 $Y=0.135
c15 2 VSS 0.0616432f $X=0.351 $Y=0.0675
r16 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.115 $X2=0.351 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AO332X1_ASAP7_75T_L%B3 2 5 7 10 VSS
c12 10 VSS 7.27237e-19 $X=0.403 $Y=0.115
c13 5 VSS 0.00111185f $X=0.405 $Y=0.135
c14 2 VSS 0.0615515f $X=0.405 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.115 $X2=0.405 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO332X1_ASAP7_75T_L%C2 2 5 7 10 VSS
c11 10 VSS 0.00167719f $X=0.46 $Y=0.114
c12 5 VSS 0.00113407f $X=0.459 $Y=0.135
c13 2 VSS 0.0618699f $X=0.459 $Y=0.0675
r14 10 13 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.114 $X2=0.459 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AO332X1_ASAP7_75T_L%C1 2 5 7 10 VSS
c11 10 VSS 4.90626e-19 $X=0.513 $Y=0.115
c12 5 VSS 0.00170409f $X=0.513 $Y=0.135
c13 2 VSS 0.0662985f $X=0.513 $Y=0.0675
r14 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.115 $X2=0.513 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AO332X1_ASAP7_75T_L%Y 1 6 9 14 16 18 21 22 28 VSS
c9 28 VSS 0.00548172f $X=0.054 $Y=0.234
c10 26 VSS 0.00317012f $X=0.027 $Y=0.234
c11 22 VSS 0.00568786f $X=0.054 $Y=0.036
c12 21 VSS 0.0078719f $X=0.054 $Y=0.036
c13 19 VSS 0.00318685f $X=0.027 $Y=0.036
c14 18 VSS 0.00230477f $X=0.018 $Y=0.2
c15 16 VSS 0.00161505f $X=0.018 $Y=0.10125
c16 15 VSS 8.29409e-19 $X=0.018 $Y=0.063
c17 14 VSS 0.00231798f $X=0.0195 $Y=0.1395
c18 12 VSS 0.00107066f $X=0.018 $Y=0.225
c19 9 VSS 0.00525295f $X=0.056 $Y=0.2025
c20 6 VSS 3.02808e-19 $X=0.071 $Y=0.2025
c21 1 VSS 2.55988e-19 $X=0.071 $Y=0.0675
r22 26 28 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.054 $Y2=0.234
r23 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r24 19 21 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.054 $Y2=0.036
r25 17 18 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.151 $X2=0.018 $Y2=0.2
r26 15 16 2.59722 $w=1.8e-08 $l=3.825e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.10125
r27 14 17 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.151
r28 14 16 2.59722 $w=1.8e-08 $l=3.825e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.10125
r29 12 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r30 12 18 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2
r31 11 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r32 11 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r33 9 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r34 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
r35 4 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r36 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./AO332x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO332x1_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 VSS N_3_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 noxref_15 N_A3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_16 N_A2_M2_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_3_M3_d N_A1_M3_g noxref_16 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_17 N_B1_M4_g N_3_M4_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_18 N_B2_M5_g noxref_17 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 VSS N_B3_M6_g noxref_18 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_19 N_C2_M7_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_3_M8_d N_C1_M8_g noxref_19 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 VDD N_3_M9_g N_Y_M9_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M10 noxref_13 N_A3_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M11 VDD N_A2_M11_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M12 noxref_13 N_A1_M12_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M13 noxref_14 N_B1_M13_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M14 noxref_13 N_B2_M14_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M15 noxref_14 N_B3_M15_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M16 N_3_M16_d N_C2_M16_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M17 noxref_14 N_C1_M17_g N_3_M17_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
*
* 
* .include "AO332x1_ASAP7_75t_L.pex.sp.AO332X1_ASAP7_75T_L.pxi"
* BEGIN of "./AO332x1_ASAP7_75t_L.pex.sp.AO332X1_ASAP7_75T_L.pxi"
* File: AO332x1_ASAP7_75t_L.pex.sp.AO332X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:07:41 2017
* 
x_PM_AO332X1_ASAP7_75T_L%3 N_3_M0_g N_3_c_2_p N_3_M9_g N_3_M4_s N_3_M3_d
+ N_3_M8_d N_3_M17_s N_3_M16_d N_3_c_42_p N_3_c_7_p N_3_c_3_p N_3_c_4_p
+ N_3_c_29_p N_3_c_32_p N_3_c_11_p N_3_c_36_p N_3_c_6_p N_3_c_35_p N_3_c_10_p
+ N_3_c_38_p N_3_c_24_p N_3_c_39_p N_3_c_13_p N_3_c_40_p N_3_c_16_p N_3_c_41_p
+ N_3_c_18_p N_3_c_20_p N_3_c_55_p N_3_c_22_p N_3_c_37_p N_3_c_23_p N_3_c_46_p
+ N_3_c_27_p VSS PM_AO332X1_ASAP7_75T_L%3
x_PM_AO332X1_ASAP7_75T_L%A3 N_A3_M1_g N_A3_c_57_n N_A3_M10_g A3 N_A3_c_63_p VSS
+ PM_AO332X1_ASAP7_75T_L%A3
x_PM_AO332X1_ASAP7_75T_L%A2 N_A2_M2_g N_A2_c_73_n N_A2_M11_g A2 N_A2_c_75_n VSS
+ PM_AO332X1_ASAP7_75T_L%A2
x_PM_AO332X1_ASAP7_75T_L%A1 N_A1_M3_g N_A1_c_89_n N_A1_M12_g A1 VSS
+ PM_AO332X1_ASAP7_75T_L%A1
x_PM_AO332X1_ASAP7_75T_L%B1 N_B1_M4_g N_B1_c_101_n N_B1_M13_g B1 VSS
+ PM_AO332X1_ASAP7_75T_L%B1
x_PM_AO332X1_ASAP7_75T_L%B2 N_B2_M5_g N_B2_c_113_n N_B2_M14_g B2 VSS
+ PM_AO332X1_ASAP7_75T_L%B2
x_PM_AO332X1_ASAP7_75T_L%B3 N_B3_M6_g N_B3_c_126_n N_B3_M15_g B3 VSS
+ PM_AO332X1_ASAP7_75T_L%B3
x_PM_AO332X1_ASAP7_75T_L%C2 N_C2_M7_g N_C2_c_138_n N_C2_M16_g C2 VSS
+ PM_AO332X1_ASAP7_75T_L%C2
x_PM_AO332X1_ASAP7_75T_L%C1 N_C1_M8_g N_C1_c_153_n N_C1_M17_g C1 VSS
+ PM_AO332X1_ASAP7_75T_L%C1
x_PM_AO332X1_ASAP7_75T_L%Y N_Y_M0_s N_Y_M9_s N_Y_c_163_p Y N_Y_c_157_n
+ N_Y_c_162_n N_Y_c_158_n N_Y_c_161_n N_Y_c_164_p VSS PM_AO332X1_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M1_g 0.00286002f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_3_c_2_p N_A3_c_57_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_3_c_3_p A3 0.00196039f $X=0.081 $Y=0.1205 $X2=0.135 $Y2=0.115
cc_4 N_3_c_4_p A3 0.00133324f $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.115
cc_5 N_3_M0_g N_A2_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 N_3_c_6_p N_A2_M2_g 3.38929e-19 $X=0.198 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_7 N_3_c_7_p A2 2.69033e-19 $X=0.081 $Y=0.106 $X2=0.135 $Y2=0.115
cc_8 N_3_c_4_p A2 7.10035e-19 $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.115
cc_9 N_3_c_6_p A2 0.00123604f $X=0.198 $Y=0.036 $X2=0.135 $Y2=0.115
cc_10 N_3_c_10_p N_A1_M3_g 2.56935e-19 $X=0.252 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_11 N_3_c_11_p A1 0.0013295f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.115
cc_12 N_3_c_10_p A1 0.00123064f $X=0.252 $Y=0.036 $X2=0.135 $Y2=0.115
cc_13 N_3_c_13_p N_B1_M4_g 2.64276e-19 $X=0.306 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_14 N_3_c_11_p B1 0.0013295f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.115
cc_15 N_3_c_13_p B1 0.00124805f $X=0.306 $Y=0.036 $X2=0.135 $Y2=0.115
cc_16 N_3_c_16_p N_B2_M5_g 3.48613e-19 $X=0.36 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_17 N_3_c_16_p B2 0.00124805f $X=0.36 $Y=0.036 $X2=0.135 $Y2=0.115
cc_18 N_3_c_18_p N_B3_M6_g 2.56935e-19 $X=0.414 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_19 N_3_c_18_p B3 0.00123064f $X=0.414 $Y=0.036 $X2=0.135 $Y2=0.115
cc_20 N_3_c_20_p N_C2_M7_g 2.56935e-19 $X=0.468 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_21 N_3_c_20_p C2 0.00123064f $X=0.468 $Y=0.036 $X2=0.135 $Y2=0.115
cc_22 N_3_c_22_p N_C1_M8_g 2.64276e-19 $X=0.522 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_23 N_3_c_23_p N_C1_M8_g 2.76185e-19 $X=0.522 $Y=0.198 $X2=0.135 $Y2=0.0675
cc_24 N_3_c_24_p C1 0.0013399f $X=0.54 $Y=0.036 $X2=0.135 $Y2=0.115
cc_25 N_3_c_22_p C1 0.00124805f $X=0.522 $Y=0.036 $X2=0.135 $Y2=0.115
cc_26 N_3_c_23_p C1 0.0012322f $X=0.522 $Y=0.198 $X2=0.135 $Y2=0.115
cc_27 N_3_c_27_p C1 0.00392202f $X=0.567 $Y=0.164 $X2=0.135 $Y2=0.115
cc_28 N_3_c_3_p Y 0.00139016f $X=0.081 $Y=0.1205 $X2=0.135 $Y2=0.135
cc_29 N_3_c_29_p N_Y_c_157_n 0.00139016f $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_30 N_3_M0_g N_Y_c_158_n 2.34993e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_3_c_29_p N_Y_c_158_n 0.00197676f $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_32 N_3_c_32_p N_Y_c_158_n 7.93849e-19 $X=0.144 $Y=0.036 $X2=0 $Y2=0
cc_33 N_3_c_29_p N_Y_c_161_n 0.00143805f $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_34 VSS N_3_c_11_p 0.00138157f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.115
cc_35 VSS N_3_c_35_p 2.30767e-19 $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_36 VSS N_3_c_36_p 2.30767e-19 $X=0.18 $Y=0.036 $X2=0 $Y2=0
cc_37 VSS N_3_c_37_p 2.9669e-19 $X=0.504 $Y=0.198 $X2=0 $Y2=0
cc_38 VSS N_3_c_38_p 2.23188e-19 $X=0.261 $Y=0.036 $X2=0 $Y2=0
cc_39 VSS N_3_c_39_p 2.23188e-19 $X=0.288 $Y=0.036 $X2=0 $Y2=0
cc_40 VSS N_3_c_40_p 2.23188e-19 $X=0.342 $Y=0.036 $X2=0 $Y2=0
cc_41 VSS N_3_c_41_p 2.23188e-19 $X=0.393 $Y=0.036 $X2=0 $Y2=0
cc_42 VSS N_3_c_42_p 0.00333582f $X=0.486 $Y=0.2025 $X2=0.135 $Y2=0.115
cc_43 VSS N_3_c_37_p 4.54465e-19 $X=0.504 $Y=0.198 $X2=0.135 $Y2=0.115
cc_44 VSS N_3_c_42_p 0.00371671f $X=0.486 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_45 VSS N_3_c_24_p 0.00138157f $X=0.54 $Y=0.036 $X2=0.135 $Y2=0.135
cc_46 VSS N_3_c_46_p 0.00284922f $X=0.556 $Y=0.198 $X2=0.135 $Y2=0.135
cc_47 VSS N_3_c_27_p 3.97918e-19 $X=0.567 $Y=0.164 $X2=0.135 $Y2=0.135
cc_48 VSS N_3_c_23_p 0.00365373f $X=0.522 $Y=0.198 $X2=0 $Y2=0
cc_49 VSS N_3_c_42_p 0.00250965f $X=0.486 $Y=0.2025 $X2=0 $Y2=0
cc_50 VSS N_3_c_37_p 0.00365373f $X=0.504 $Y=0.198 $X2=0 $Y2=0
cc_51 VSS N_3_c_36_p 3.56327e-19 $X=0.18 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_52 VSS N_3_c_35_p 3.56327e-19 $X=0.234 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_53 VSS N_3_c_40_p 3.48201e-19 $X=0.342 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_54 VSS N_3_c_41_p 3.30547e-19 $X=0.393 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_55 VSS N_3_c_55_p 3.30547e-19 $X=0.504 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_56 N_A3_M1_g N_A2_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_57 N_A3_c_57_n N_A2_c_73_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_58 A3 A2 0.00196244f $X=0.135 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_59 N_A3_c_63_p N_A2_c_75_n 0.00196244f $X=0.135 $Y=0.135 $X2=0.538 $Y2=0.0675
cc_60 N_A3_M1_g N_A1_M3_g 2.66145e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_61 N_A3_c_63_p N_Y_c_162_n 4.56551e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_62 VSS N_A3_c_63_p 0.00114532f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_63 N_A2_M2_g N_A1_M3_g 0.00327995f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_64 N_A2_c_73_n N_A1_c_89_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_65 A2 A1 0.00464977f $X=0.189 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_66 N_A2_M2_g N_B1_M4_g 2.71887e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_67 VSS A2 0.0011319f $X=0.189 $Y=0.115 $X2=0.081 $Y2=0.135
cc_68 VSS N_A2_M2_g 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_69 VSS N_A2_c_75_n 0.00125352f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_70 VSS N_A2_c_75_n 4.64812e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_71 N_A1_M3_g N_B1_M4_g 0.0036939f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_72 N_A1_c_89_n N_B1_c_101_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_73 A1 B1 0.00406615f $X=0.243 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_74 N_A1_M3_g N_B2_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_75 VSS A1 0.00159458f $X=0.243 $Y=0.115 $X2=0.081 $Y2=0.135
cc_76 N_B1_M4_g N_B2_M5_g 0.00371573f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_77 N_B1_c_101_n N_B2_c_113_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_78 B1 B2 0.00483372f $X=0.297 $Y=0.116 $X2=0.253 $Y2=0.0675
cc_79 N_B1_M4_g N_B3_M6_g 3.06651e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_80 VSS N_B1_M4_g 3.62029e-19 $X=0.297 $Y=0.0675 $X2=0.094 $Y2=0.072
cc_81 VSS B1 0.0012322f $X=0.297 $Y=0.116 $X2=0.094 $Y2=0.072
cc_82 N_B2_M5_g N_B3_M6_g 0.0036939f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_83 N_B2_c_113_n N_B3_c_126_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_84 B2 B3 0.00483372f $X=0.35 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_85 N_B2_M5_g N_C2_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_86 VSS N_B2_M5_g 2.68514e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.063
cc_87 VSS B2 0.00121543f $X=0.35 $Y=0.115 $X2=0.135 $Y2=0.063
cc_88 VSS N_B2_M5_g 2.38303e-19 $X=0.351 $Y=0.0675 $X2=0.486 $Y2=0.2025
cc_89 N_B3_M6_g N_C2_M7_g 0.00333077f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_90 N_B3_c_126_n N_C2_c_138_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_91 B3 C2 0.00406615f $X=0.403 $Y=0.115 $X2=0.253 $Y2=0.0675
cc_92 N_B3_M6_g N_C1_M8_g 2.71887e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_93 VSS N_B3_M6_g 3.47199e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_94 VSS B3 5.30079e-19 $X=0.403 $Y=0.115 $X2=0.081 $Y2=0.135
cc_95 N_C2_M7_g N_C1_M8_g 0.0036939f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_96 N_C2_c_138_n N_C1_c_153_n 9.33263e-19 $X=0.459 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_97 C2 C1 0.00477924f $X=0.46 $Y=0.114 $X2=0.253 $Y2=0.0675
cc_98 VSS N_C2_M7_g 3.57119e-19 $X=0.459 $Y=0.0675 $X2=0.126 $Y2=0.072
cc_99 VSS C2 5.37372e-19 $X=0.46 $Y=0.114 $X2=0.126 $Y2=0.072
cc_100 VSS N_C1_M8_g 2.15135e-19 $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.106
cc_101 VSS N_Y_c_163_p 2.2337e-19 $X=0.056 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_102 VSS N_Y_c_164_p 2.82839e-19 $X=0.054 $Y=0.234 $X2=0.486 $Y2=0.2025

* END of "./AO332x1_ASAP7_75t_L.pex.sp.AO332X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO332x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:08:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO332x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO332x2_ASAP7_75t_L.pex.sp.pex"
* File: AO332x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:08:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO332X2_ASAP7_75T_L%3 2 7 10 13 15 17 18 22 27 28 31 36 37 39 40 46
+ 49 51 52 53 54 55 58 59 60 61 62 63 65 67 69 70 76 77 78 83 VSS
c65 83 VSS 0.00412141f $X=0.621 $Y=0.164
c66 82 VSS 9.6701e-19 $X=0.621 $Y=0.07
c67 81 VSS 0.00112176f $X=0.621 $Y=0.189
c68 79 VSS 4.93718e-20 $X=0.611 $Y=0.198
c69 78 VSS 4.1269e-19 $X=0.61 $Y=0.198
c70 77 VSS 8.46035e-21 $X=0.576 $Y=0.198
c71 76 VSS 4.70878e-19 $X=0.558 $Y=0.198
c72 71 VSS 0.0019286f $X=0.612 $Y=0.198
c73 70 VSS 0.00146362f $X=0.576 $Y=0.036
c74 69 VSS 0.00296425f $X=0.558 $Y=0.036
c75 68 VSS 3.35992e-19 $X=0.525 $Y=0.036
c76 67 VSS 0.00142296f $X=0.522 $Y=0.036
c77 66 VSS 0.00672869f $X=0.504 $Y=0.036
c78 65 VSS 0.00142296f $X=0.468 $Y=0.036
c79 64 VSS 3.35992e-19 $X=0.45 $Y=0.036
c80 63 VSS 0.00311761f $X=0.447 $Y=0.036
c81 62 VSS 0.00146362f $X=0.414 $Y=0.036
c82 61 VSS 0.00340162f $X=0.396 $Y=0.036
c83 60 VSS 0.00146362f $X=0.36 $Y=0.036
c84 59 VSS 0.00256536f $X=0.342 $Y=0.036
c85 58 VSS 0.00357414f $X=0.594 $Y=0.036
c86 55 VSS 8.84964e-19 $X=0.315 $Y=0.036
c87 54 VSS 0.00142296f $X=0.306 $Y=0.036
c88 53 VSS 0.00360252f $X=0.288 $Y=0.036
c89 52 VSS 0.00142296f $X=0.252 $Y=0.036
c90 51 VSS 0.00331443f $X=0.234 $Y=0.036
c91 50 VSS 1.51923e-19 $X=0.2 $Y=0.036
c92 49 VSS 0.00220219f $X=0.324 $Y=0.036
c93 46 VSS 0.00233672f $X=0.198 $Y=0.036
c94 45 VSS 0.00702647f $X=0.612 $Y=0.036
c95 44 VSS 9.0336e-19 $X=0.189 $Y=0.063
c96 42 VSS 0.00182969f $X=0.164 $Y=0.072
c97 41 VSS 8.41473e-20 $X=0.148 $Y=0.072
c98 40 VSS 4.67384e-20 $X=0.144 $Y=0.072
c99 39 VSS 0.00174552f $X=0.18 $Y=0.072
c100 37 VSS 1.76256e-19 $X=0.135 $Y=0.1205
c101 36 VSS 9.91953e-19 $X=0.135 $Y=0.106
c102 34 VSS 4.07276e-19 $X=0.135 $Y=0.135
c103 31 VSS 0.0023085f $X=0.54 $Y=0.2025
c104 27 VSS 5.70099e-19 $X=0.557 $Y=0.2025
c105 25 VSS 2.69461e-19 $X=0.592 $Y=0.0675
c106 17 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c107 13 VSS 0.00397026f $X=0.135 $Y=0.135
c108 10 VSS 0.0608916f $X=0.135 $Y=0.0675
c109 2 VSS 0.0615048f $X=0.081 $Y=0.0675
r110 82 83 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.07 $X2=0.621 $Y2=0.164
r111 81 83 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.189 $X2=0.621 $Y2=0.164
r112 80 82 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.07
r113 78 79 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.61
+ $Y=0.198 $X2=0.611 $Y2=0.198
r114 77 78 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.198 $X2=0.61 $Y2=0.198
r115 76 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.198 $X2=0.576 $Y2=0.198
r116 73 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.198 $X2=0.558 $Y2=0.198
r117 71 81 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.198 $X2=0.621 $Y2=0.189
r118 71 79 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.198 $X2=0.611 $Y2=0.198
r119 69 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.576 $Y2=0.036
r120 68 69 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.525
+ $Y=0.036 $X2=0.558 $Y2=0.036
r121 67 68 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.525 $Y2=0.036
r122 66 67 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.522 $Y2=0.036
r123 65 66 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.504 $Y2=0.036
r124 64 65 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r125 63 64 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.036 $X2=0.45 $Y2=0.036
r126 62 63 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.447 $Y2=0.036
r127 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r128 60 61 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.396 $Y2=0.036
r129 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r130 57 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.576 $Y2=0.036
r131 57 58 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036
+ $X2=0.594 $Y2=0.036
r132 54 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.315 $Y2=0.036
r133 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r134 52 53 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r135 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r136 50 51 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2
+ $Y=0.036 $X2=0.234 $Y2=0.036
r137 48 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r138 48 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.315 $Y2=0.036
r139 48 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r140 46 50 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.2 $Y2=0.036
r141 45 80 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r142 45 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.594 $Y2=0.036
r143 43 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.045 $X2=0.198 $Y2=0.036
r144 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r145 41 42 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.072 $X2=0.164 $Y2=0.072
r146 40 41 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.148 $Y2=0.072
r147 39 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.072 $X2=0.189 $Y2=0.063
r148 39 42 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.072 $X2=0.164 $Y2=0.072
r149 36 37 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.106 $X2=0.135 $Y2=0.1205
r150 34 37 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.1205
r151 32 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.081 $X2=0.144 $Y2=0.072
r152 32 36 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.081 $X2=0.135 $Y2=0.106
r153 31 73 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.198 $X2=0.54
+ $Y2=0.198
r154 28 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r155 27 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r156 25 58 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.594 $Y=0.0675 $X2=0.594 $Y2=0.036
r157 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0675 $X2=0.592 $Y2=0.0675
r158 21 49 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r159 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r160 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r161 13 34 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r162 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r163 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r164 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r165 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r166 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO332X2_ASAP7_75T_L%A3 2 5 7 10 13 VSS
c12 13 VSS 0.00246747f $X=0.189 $Y=0.135
c13 10 VSS 3.14219e-19 $X=0.189 $Y=0.115
c14 5 VSS 0.0011078f $X=0.189 $Y=0.135
c15 2 VSS 0.0588833f $X=0.189 $Y=0.0675
r16 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO332X2_ASAP7_75T_L%A2 2 5 7 10 15 VSS
c17 15 VSS 0.00159343f $X=0.243 $Y=0.135
c18 10 VSS 7.68637e-19 $X=0.243 $Y=0.115
c19 5 VSS 0.00111216f $X=0.243 $Y=0.135
c20 2 VSS 0.059482f $X=0.243 $Y=0.0675
r21 10 15 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.115 $X2=0.243 $Y2=0.135
r22 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r23 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r24 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO332X2_ASAP7_75T_L%A1 2 5 7 10 VSS
c12 10 VSS 4.82288e-19 $X=0.297 $Y=0.115
c13 5 VSS 0.00111383f $X=0.297 $Y=0.135
c14 2 VSS 0.0608471f $X=0.297 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.115 $X2=0.297 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO332X2_ASAP7_75T_L%B1 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.351 $Y=0.116
c14 5 VSS 0.00111336f $X=0.351 $Y=0.135
c15 2 VSS 0.0617786f $X=0.351 $Y=0.0675
r16 10 13 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.116 $X2=0.351 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AO332X2_ASAP7_75T_L%B2 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.404 $Y=0.115
c14 5 VSS 0.00112198f $X=0.405 $Y=0.135
c15 2 VSS 0.0616432f $X=0.405 $Y=0.0675
r16 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.115 $X2=0.405 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO332X2_ASAP7_75T_L%B3 2 5 7 10 VSS
c12 10 VSS 7.27237e-19 $X=0.457 $Y=0.115
c13 5 VSS 0.00111185f $X=0.459 $Y=0.135
c14 2 VSS 0.0615515f $X=0.459 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.115 $X2=0.459 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AO332X2_ASAP7_75T_L%C2 2 5 7 10 VSS
c11 10 VSS 0.00167719f $X=0.514 $Y=0.114
c12 5 VSS 0.00113407f $X=0.513 $Y=0.135
c13 2 VSS 0.0618699f $X=0.513 $Y=0.0675
r14 10 13 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.114 $X2=0.513 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AO332X2_ASAP7_75T_L%C1 2 5 7 10 VSS
c11 10 VSS 4.90626e-19 $X=0.567 $Y=0.115
c12 5 VSS 0.00170409f $X=0.567 $Y=0.135
c13 2 VSS 0.0662985f $X=0.567 $Y=0.0675
r14 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.115 $X2=0.567 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
.ends

.subckt PM_AO332X2_ASAP7_75T_L%Y 1 2 6 7 10 14 16 18 21 22 28 VSS
c18 28 VSS 0.0131561f $X=0.108 $Y=0.234
c19 26 VSS 0.00320021f $X=0.027 $Y=0.234
c20 22 VSS 0.0102944f $X=0.108 $Y=0.036
c21 21 VSS 0.0154624f $X=0.108 $Y=0.036
c22 19 VSS 0.0032101f $X=0.027 $Y=0.036
c23 18 VSS 0.00278197f $X=0.018 $Y=0.2
c24 16 VSS 0.00196447f $X=0.018 $Y=0.10125
c25 15 VSS 8.29409e-19 $X=0.018 $Y=0.063
c26 14 VSS 0.0025255f $X=0.0195 $Y=0.1395
c27 12 VSS 0.00126561f $X=0.018 $Y=0.225
c28 10 VSS 0.00902033f $X=0.108 $Y=0.2025
c29 6 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c30 1 VSS 5.25448e-19 $X=0.125 $Y=0.0675
r31 26 28 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.108 $Y2=0.234
r32 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r33 19 21 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.108 $Y2=0.036
r34 17 18 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.151 $X2=0.018 $Y2=0.2
r35 15 16 2.59722 $w=1.8e-08 $l=3.825e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.10125
r36 14 17 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.151
r37 14 16 2.59722 $w=1.8e-08 $l=3.825e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.10125
r38 12 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r39 12 18 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2
r40 11 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r41 11 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r42 10 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r43 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r44 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r45 5 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r46 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r47 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./AO332x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO332x2_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_15 N_A3_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_16 N_A2_M3_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_3_M4_d N_A1_M4_g noxref_16 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_17 N_B1_M5_g N_3_M5_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_18 N_B2_M6_g noxref_17 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 VSS N_B3_M7_g noxref_18 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 noxref_19 N_C2_M8_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 N_3_M9_d N_C1_M9_g noxref_19 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M10 N_Y_M10_d N_3_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M11 N_Y_M11_d N_3_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M12 noxref_13 N_A3_M12_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M13 VDD N_A2_M13_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M14 noxref_13 N_A1_M14_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M15 noxref_14 N_B1_M15_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M16 noxref_13 N_B2_M16_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M17 noxref_14 N_B3_M17_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M18 N_3_M18_d N_C2_M18_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
M19 noxref_14 N_C1_M19_g N_3_M19_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
*
* 
* .include "AO332x2_ASAP7_75t_L.pex.sp.AO332X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO332x2_ASAP7_75t_L.pex.sp.AO332X2_ASAP7_75T_L.pxi"
* File: AO332x2_ASAP7_75t_L.pex.sp.AO332X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:08:03 2017
* 
x_PM_AO332X2_ASAP7_75T_L%3 N_3_M0_g N_3_M10_g N_3_M1_g N_3_c_3_p N_3_M11_g
+ N_3_M5_s N_3_M4_d N_3_M9_d N_3_M19_s N_3_M18_d N_3_c_52_p N_3_c_8_p N_3_c_4_p
+ N_3_c_5_p N_3_c_34_p N_3_c_39_p N_3_c_12_p N_3_c_46_p N_3_c_7_p N_3_c_45_p
+ N_3_c_11_p N_3_c_48_p N_3_c_25_p N_3_c_49_p N_3_c_14_p N_3_c_50_p N_3_c_17_p
+ N_3_c_51_p N_3_c_19_p N_3_c_21_p N_3_c_65_p N_3_c_23_p N_3_c_47_p N_3_c_24_p
+ N_3_c_56_p N_3_c_28_p VSS PM_AO332X2_ASAP7_75T_L%3
x_PM_AO332X2_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_68_n N_A3_M12_g A3 N_A3_c_74_p VSS
+ PM_AO332X2_ASAP7_75T_L%A3
x_PM_AO332X2_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_84_n N_A2_M13_g A2 N_A2_c_86_n VSS
+ PM_AO332X2_ASAP7_75T_L%A2
x_PM_AO332X2_ASAP7_75T_L%A1 N_A1_M4_g N_A1_c_100_n N_A1_M14_g A1 VSS
+ PM_AO332X2_ASAP7_75T_L%A1
x_PM_AO332X2_ASAP7_75T_L%B1 N_B1_M5_g N_B1_c_112_n N_B1_M15_g B1 VSS
+ PM_AO332X2_ASAP7_75T_L%B1
x_PM_AO332X2_ASAP7_75T_L%B2 N_B2_M6_g N_B2_c_124_n N_B2_M16_g B2 VSS
+ PM_AO332X2_ASAP7_75T_L%B2
x_PM_AO332X2_ASAP7_75T_L%B3 N_B3_M7_g N_B3_c_137_n N_B3_M17_g B3 VSS
+ PM_AO332X2_ASAP7_75T_L%B3
x_PM_AO332X2_ASAP7_75T_L%C2 N_C2_M8_g N_C2_c_149_n N_C2_M18_g C2 VSS
+ PM_AO332X2_ASAP7_75T_L%C2
x_PM_AO332X2_ASAP7_75T_L%C1 N_C1_M9_g N_C1_c_164_n N_C1_M19_g C1 VSS
+ PM_AO332X2_ASAP7_75T_L%C1
x_PM_AO332X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_M11_d N_Y_M10_d N_Y_c_169_n Y
+ N_Y_c_172_n N_Y_c_182_n N_Y_c_173_n N_Y_c_178_n N_Y_c_180_n VSS
+ PM_AO332X2_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M2_g 2.13359e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_A3_M2_g 0.00286002f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_A3_c_68_n 9.59209e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_4 N_3_c_4_p A3 0.00196257f $X=0.135 $Y=0.1205 $X2=0.189 $Y2=0.115
cc_5 N_3_c_5_p A3 0.00133324f $X=0.18 $Y=0.072 $X2=0.189 $Y2=0.115
cc_6 N_3_M1_g N_A2_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_7 N_3_c_7_p N_A2_M3_g 3.38929e-19 $X=0.252 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_8 N_3_c_8_p A2 2.69033e-19 $X=0.135 $Y=0.106 $X2=0.189 $Y2=0.115
cc_9 N_3_c_5_p A2 7.10035e-19 $X=0.18 $Y=0.072 $X2=0.189 $Y2=0.115
cc_10 N_3_c_7_p A2 0.00123604f $X=0.252 $Y=0.036 $X2=0.189 $Y2=0.115
cc_11 N_3_c_11_p N_A1_M4_g 2.56935e-19 $X=0.306 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_12 N_3_c_12_p A1 0.0013295f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.115
cc_13 N_3_c_11_p A1 0.00123064f $X=0.306 $Y=0.036 $X2=0.189 $Y2=0.115
cc_14 N_3_c_14_p N_B1_M5_g 2.64276e-19 $X=0.36 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_15 N_3_c_12_p B1 0.0013295f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.115
cc_16 N_3_c_14_p B1 0.00124805f $X=0.36 $Y=0.036 $X2=0.189 $Y2=0.115
cc_17 N_3_c_17_p N_B2_M6_g 3.48613e-19 $X=0.414 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_18 N_3_c_17_p B2 0.00124805f $X=0.414 $Y=0.036 $X2=0.189 $Y2=0.115
cc_19 N_3_c_19_p N_B3_M7_g 2.56935e-19 $X=0.468 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_20 N_3_c_19_p B3 0.00123064f $X=0.468 $Y=0.036 $X2=0.189 $Y2=0.115
cc_21 N_3_c_21_p N_C2_M8_g 2.56935e-19 $X=0.522 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_22 N_3_c_21_p C2 0.00123064f $X=0.522 $Y=0.036 $X2=0.189 $Y2=0.115
cc_23 N_3_c_23_p N_C1_M9_g 2.64276e-19 $X=0.576 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_24 N_3_c_24_p N_C1_M9_g 2.76185e-19 $X=0.576 $Y=0.198 $X2=0.189 $Y2=0.0675
cc_25 N_3_c_25_p C1 0.0013399f $X=0.594 $Y=0.036 $X2=0.189 $Y2=0.115
cc_26 N_3_c_23_p C1 0.00124805f $X=0.576 $Y=0.036 $X2=0.189 $Y2=0.115
cc_27 N_3_c_24_p C1 0.0012322f $X=0.576 $Y=0.198 $X2=0.189 $Y2=0.115
cc_28 N_3_c_28_p C1 0.00392202f $X=0.621 $Y=0.164 $X2=0.189 $Y2=0.115
cc_29 N_3_c_3_p N_Y_M1_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_30 N_3_c_3_p N_Y_M11_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_31 N_3_c_3_p N_Y_c_169_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.115
cc_32 N_3_c_3_p Y 3.36333e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_33 N_3_c_4_p Y 4.74317e-19 $X=0.135 $Y=0.1205 $X2=0.189 $Y2=0.135
cc_34 N_3_c_34_p N_Y_c_172_n 4.74317e-19 $X=0.144 $Y=0.072 $X2=0 $Y2=0
cc_35 N_3_M0_g N_Y_c_173_n 4.59284e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_3_M1_g N_Y_c_173_n 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_3_c_3_p N_Y_c_173_n 5.94649e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_38 N_3_c_34_p N_Y_c_173_n 0.00197676f $X=0.144 $Y=0.072 $X2=0 $Y2=0
cc_39 N_3_c_39_p N_Y_c_173_n 8.21768e-19 $X=0.198 $Y=0.036 $X2=0 $Y2=0
cc_40 N_3_c_3_p N_Y_c_178_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_41 N_3_c_34_p N_Y_c_178_n 0.0015778f $X=0.144 $Y=0.072 $X2=0 $Y2=0
cc_42 N_3_M0_g N_Y_c_180_n 4.59284e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_3_c_3_p N_Y_c_180_n 5.35059e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_44 VSS N_3_c_12_p 0.00138157f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.115
cc_45 VSS N_3_c_45_p 2.30767e-19 $X=0.288 $Y=0.036 $X2=0 $Y2=0
cc_46 VSS N_3_c_46_p 2.30767e-19 $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_47 VSS N_3_c_47_p 2.9669e-19 $X=0.558 $Y=0.198 $X2=0 $Y2=0
cc_48 VSS N_3_c_48_p 2.23188e-19 $X=0.315 $Y=0.036 $X2=0 $Y2=0
cc_49 VSS N_3_c_49_p 2.23188e-19 $X=0.342 $Y=0.036 $X2=0 $Y2=0
cc_50 VSS N_3_c_50_p 2.23188e-19 $X=0.396 $Y=0.036 $X2=0 $Y2=0
cc_51 VSS N_3_c_51_p 2.23188e-19 $X=0.447 $Y=0.036 $X2=0 $Y2=0
cc_52 VSS N_3_c_52_p 0.00333582f $X=0.54 $Y=0.2025 $X2=0.189 $Y2=0.115
cc_53 VSS N_3_c_47_p 4.54465e-19 $X=0.558 $Y=0.198 $X2=0.189 $Y2=0.115
cc_54 VSS N_3_c_52_p 0.00371671f $X=0.54 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_55 VSS N_3_c_25_p 0.00138157f $X=0.594 $Y=0.036 $X2=0.189 $Y2=0.135
cc_56 VSS N_3_c_56_p 0.00284922f $X=0.61 $Y=0.198 $X2=0.189 $Y2=0.135
cc_57 VSS N_3_c_28_p 3.97918e-19 $X=0.621 $Y=0.164 $X2=0.189 $Y2=0.135
cc_58 VSS N_3_c_24_p 0.00365373f $X=0.576 $Y=0.198 $X2=0 $Y2=0
cc_59 VSS N_3_c_52_p 0.00250965f $X=0.54 $Y=0.2025 $X2=0 $Y2=0
cc_60 VSS N_3_c_47_p 0.00365373f $X=0.558 $Y=0.198 $X2=0 $Y2=0
cc_61 VSS N_3_c_46_p 3.56327e-19 $X=0.234 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_62 VSS N_3_c_45_p 3.56327e-19 $X=0.288 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_63 VSS N_3_c_50_p 3.48201e-19 $X=0.396 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_64 VSS N_3_c_51_p 3.30547e-19 $X=0.447 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_65 VSS N_3_c_65_p 3.30547e-19 $X=0.558 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_66 N_A3_M2_g N_A2_M3_g 0.00344695f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_67 N_A3_c_68_n N_A2_c_84_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_68 A3 A2 0.00196244f $X=0.189 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_69 N_A3_c_74_p N_A2_c_86_n 0.00196244f $X=0.189 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_70 N_A3_M2_g N_A1_M4_g 2.66145e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_71 N_A3_c_74_p N_Y_c_182_n 2.26084e-19 $X=0.189 $Y=0.135 $X2=0.307 $Y2=0.0675
cc_72 VSS N_A3_c_74_p 0.00114532f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_73 N_A2_M3_g N_A1_M4_g 0.00327995f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_74 N_A2_c_84_n N_A1_c_100_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_75 A2 A1 0.00464977f $X=0.243 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_76 N_A2_M3_g N_B1_M5_g 2.71887e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_77 VSS A2 0.0011319f $X=0.243 $Y=0.115 $X2=0.081 $Y2=0.135
cc_78 VSS N_A2_M3_g 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0.577 $Y2=0.0675
cc_79 VSS N_A2_c_86_n 0.00125352f $X=0.243 $Y=0.135 $X2=0.577 $Y2=0.0675
cc_80 VSS N_A2_c_86_n 4.64812e-19 $X=0.243 $Y=0.135 $X2=0.592 $Y2=0.0675
cc_81 N_A1_M4_g N_B1_M5_g 0.0036939f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_82 N_A1_c_100_n N_B1_c_112_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_83 A1 B1 0.00406615f $X=0.297 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_84 N_A1_M4_g N_B2_M6_g 3.06651e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_85 VSS A1 0.00159458f $X=0.297 $Y=0.115 $X2=0.592 $Y2=0.0675
cc_86 N_B1_M5_g N_B2_M6_g 0.00371573f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_87 N_B1_c_112_n N_B2_c_124_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_88 B1 B2 0.00483372f $X=0.351 $Y=0.116 $X2=0.135 $Y2=0.0675
cc_89 N_B1_M5_g N_B3_M7_g 3.06651e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_90 VSS N_B1_M5_g 3.62029e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_91 VSS B1 0.0012322f $X=0.351 $Y=0.116 $X2=0.135 $Y2=0.135
cc_92 N_B2_M6_g N_B3_M7_g 0.0036939f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_93 N_B2_c_124_n N_B3_c_137_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_94 B2 B3 0.00483372f $X=0.404 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_95 N_B2_M6_g N_C2_M8_g 2.71887e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_96 VSS N_B2_M6_g 2.68514e-19 $X=0.405 $Y=0.0675 $X2=0.135 $Y2=0.106
cc_97 VSS B2 0.00121543f $X=0.404 $Y=0.115 $X2=0.135 $Y2=0.106
cc_98 VSS N_B2_M6_g 2.38303e-19 $X=0.405 $Y=0.0675 $X2=0.592 $Y2=0.0675
cc_99 N_B3_M7_g N_C2_M8_g 0.00333077f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_100 N_B3_c_137_n N_C2_c_149_n 8.86777e-19 $X=0.459 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_101 B3 C2 0.00406615f $X=0.457 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_102 N_B3_M7_g N_C1_M9_g 2.71887e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_103 VSS N_B3_M7_g 3.47199e-19 $X=0.459 $Y=0.0675 $X2=0.592 $Y2=0.0675
cc_104 VSS B3 5.30079e-19 $X=0.457 $Y=0.115 $X2=0.592 $Y2=0.0675
cc_105 N_C2_M8_g N_C1_M9_g 0.0036939f $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_106 N_C2_c_149_n N_C1_c_164_n 9.33263e-19 $X=0.513 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_107 C2 C1 0.00477924f $X=0.514 $Y=0.114 $X2=0.135 $Y2=0.0675
cc_108 VSS N_C2_M8_g 3.57119e-19 $X=0.513 $Y=0.0675 $X2=0.54 $Y2=0.2025
cc_109 VSS C2 5.37372e-19 $X=0.514 $Y=0.114 $X2=0.54 $Y2=0.2025
cc_110 VSS N_C1_M9_g 2.15135e-19 $X=0.567 $Y=0.0675 $X2=0.523 $Y2=0.2025
cc_111 VSS N_Y_c_169_n 2.23372e-19 $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_112 VSS N_Y_c_180_n 2.93728e-19 $X=0.108 $Y=0.234 $X2=0.324 $Y2=0.0675

* END of "./AO332x2_ASAP7_75t_L.pex.sp.AO332X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO333x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:08:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO333x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO333x1_ASAP7_75t_L.pex.sp.pex"
* File: AO333x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:08:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO333X1_ASAP7_75T_L%3 2 5 7 9 10 14 19 20 23 24 27 33 34 36 37 41 44
+ 46 47 48 49 53 55 57 58 59 60 61 62 63 64 65 66 76 81 83 VSS
c57 83 VSS 6.70384e-19 $X=0.621 $Y=0.207
c58 82 VSS 0.00104083f $X=0.621 $Y=0.189
c59 81 VSS 0.00414971f $X=0.621 $Y=0.164
c60 80 VSS 9.73652e-19 $X=0.621 $Y=0.07
c61 79 VSS 8.85605e-19 $X=0.621 $Y=0.225
c62 77 VSS 8.42643e-19 $X=0.585 $Y=0.234
c63 76 VSS 0.00886015f $X=0.576 $Y=0.234
c64 68 VSS 0.00606021f $X=0.612 $Y=0.234
c65 67 VSS 8.42643e-19 $X=0.585 $Y=0.036
c66 66 VSS 0.00142296f $X=0.576 $Y=0.036
c67 65 VSS 0.00346807f $X=0.558 $Y=0.036
c68 64 VSS 0.00142296f $X=0.522 $Y=0.036
c69 63 VSS 0.00330791f $X=0.504 $Y=0.036
c70 62 VSS 0.00142296f $X=0.468 $Y=0.036
c71 61 VSS 0.0068014f $X=0.45 $Y=0.036
c72 60 VSS 0.00142296f $X=0.414 $Y=0.036
c73 59 VSS 0.00346807f $X=0.396 $Y=0.036
c74 58 VSS 0.00142296f $X=0.36 $Y=0.036
c75 57 VSS 0.00309345f $X=0.342 $Y=0.036
c76 56 VSS 3.54965e-19 $X=0.31 $Y=0.036
c77 55 VSS 0.00146362f $X=0.306 $Y=0.036
c78 54 VSS 0.00274772f $X=0.288 $Y=0.036
c79 53 VSS 0.00224055f $X=0.594 $Y=0.036
c80 50 VSS 0.00106066f $X=0.261 $Y=0.036
c81 49 VSS 0.00142296f $X=0.252 $Y=0.036
c82 48 VSS 0.00376615f $X=0.234 $Y=0.036
c83 47 VSS 0.00142296f $X=0.198 $Y=0.036
c84 46 VSS 0.00329341f $X=0.18 $Y=0.036
c85 45 VSS 3.78291e-19 $X=0.148 $Y=0.036
c86 44 VSS 0.00218387f $X=0.27 $Y=0.036
c87 41 VSS 0.00238558f $X=0.144 $Y=0.036
c88 40 VSS 0.00612605f $X=0.612 $Y=0.036
c89 39 VSS 9.0336e-19 $X=0.135 $Y=0.063
c90 37 VSS 3.49137e-19 $X=0.09 $Y=0.072
c91 36 VSS 0.00381214f $X=0.126 $Y=0.072
c92 34 VSS 1.71139e-19 $X=0.081 $Y=0.1205
c93 33 VSS 9.91953e-19 $X=0.081 $Y=0.106
c94 31 VSS 4.09835e-19 $X=0.081 $Y=0.135
c95 27 VSS 0.00257027f $X=0.592 $Y=0.2025
c96 23 VSS 0.00238723f $X=0.486 $Y=0.2025
c97 19 VSS 7.12337e-19 $X=0.503 $Y=0.2025
c98 17 VSS 2.69461e-19 $X=0.592 $Y=0.0675
c99 9 VSS 5.38922e-19 $X=0.287 $Y=0.0675
c100 5 VSS 0.00182168f $X=0.081 $Y=0.135
c101 2 VSS 0.0623882f $X=0.081 $Y=0.0675
r102 82 83 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.189 $X2=0.621 $Y2=0.207
r103 81 82 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.164 $X2=0.621 $Y2=0.189
r104 80 81 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.07 $X2=0.621 $Y2=0.164
r105 79 83 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.207
r106 78 80 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.07
r107 76 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.234 $X2=0.585 $Y2=0.234
r108 74 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.585 $Y2=0.234
r109 70 76 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.576 $Y2=0.234
r110 68 79 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r111 68 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r112 66 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.036 $X2=0.585 $Y2=0.036
r113 65 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.576 $Y2=0.036
r114 64 65 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.558 $Y2=0.036
r115 63 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.522 $Y2=0.036
r116 62 63 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.504 $Y2=0.036
r117 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r118 60 61 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.45 $Y2=0.036
r119 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r120 58 59 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.396 $Y2=0.036
r121 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r122 56 57 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.31
+ $Y=0.036 $X2=0.342 $Y2=0.036
r123 55 56 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.31 $Y2=0.036
r124 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r125 52 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.585 $Y2=0.036
r126 52 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036
+ $X2=0.594 $Y2=0.036
r127 49 50 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.261 $Y2=0.036
r128 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r129 47 48 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.234 $Y2=0.036
r130 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r131 45 46 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.036 $X2=0.18 $Y2=0.036
r132 43 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.288 $Y2=0.036
r133 43 50 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.261 $Y2=0.036
r134 43 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r135 41 45 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.148 $Y2=0.036
r136 40 78 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r137 40 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.594 $Y2=0.036
r138 38 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.045 $X2=0.144 $Y2=0.036
r139 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.063
r140 36 39 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.063
r141 36 37 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.09 $Y2=0.072
r142 33 34 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.106 $X2=0.081 $Y2=0.1205
r143 31 34 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1205
r144 29 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.081 $X2=0.09 $Y2=0.072
r145 29 33 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.081 $X2=0.081 $Y2=0.106
r146 27 74 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r147 24 27 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2025 $X2=0.592 $Y2=0.2025
r148 23 70 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234
+ $X2=0.486 $Y2=0.234
r149 20 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.486 $Y2=0.2025
r150 19 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.2025 $X2=0.486 $Y2=0.2025
r151 17 53 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.594 $Y=0.0675 $X2=0.594 $Y2=0.036
r152 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0675 $X2=0.592 $Y2=0.0675
r153 13 44 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r154 10 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r155 9 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r156 5 31 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r157 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r158 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO333X1_ASAP7_75T_L%A3 2 5 7 10 14 VSS
c10 14 VSS 0.00225541f $X=0.1365 $Y=0.1485
c11 10 VSS 2.57666e-19 $X=0.135 $Y=0.135
c12 5 VSS 0.00123086f $X=0.135 $Y=0.135
c13 2 VSS 0.057276f $X=0.135 $Y=0.0675
r14 10 14 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.1485
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AO333X1_ASAP7_75T_L%A2 2 5 7 10 16 VSS
c15 10 VSS 0.00193643f $X=0.189 $Y=0.135
c16 5 VSS 0.00110907f $X=0.189 $Y=0.135
c17 2 VSS 0.057046f $X=0.189 $Y=0.0675
r18 10 16 3.49691 $w=1.8e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.1865
r19 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r20 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r21 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO333X1_ASAP7_75T_L%A1 2 5 7 10 VSS
c15 10 VSS 0.00153576f $X=0.2435 $Y=0.1345
c16 5 VSS 0.00110983f $X=0.243 $Y=0.135
c17 2 VSS 0.058107f $X=0.243 $Y=0.0675
r18 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r19 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r20 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO333X1_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c13 10 VSS 5.08499e-19 $X=0.297 $Y=0.135
c14 5 VSS 0.0011055f $X=0.297 $Y=0.135
c15 2 VSS 0.0591416f $X=0.297 $Y=0.0675
r16 10 14 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.1545
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO333X1_ASAP7_75T_L%B2 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.3505 $Y=0.0845
c14 5 VSS 0.00164678f $X=0.351 $Y=0.135
c15 2 VSS 0.0591416f $X=0.351 $Y=0.0675
r16 10 13 3.42901 $w=1.8e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.0845 $X2=0.351 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AO333X1_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c12 10 VSS 6.96915e-19 $X=0.405 $Y=0.135
c13 5 VSS 0.00164704f $X=0.405 $Y=0.135
c14 2 VSS 0.0594389f $X=0.405 $Y=0.0675
r15 10 14 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.1555
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO333X1_ASAP7_75T_L%C3 2 5 7 10 VSS
c12 10 VSS 6.96915e-19 $X=0.4565 $Y=0.0835
c13 5 VSS 0.00160703f $X=0.459 $Y=0.135
c14 2 VSS 0.0592509f $X=0.459 $Y=0.0675
r15 10 13 3.49691 $w=1.8e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.0835 $X2=0.459 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AO333X1_ASAP7_75T_L%C2 2 5 7 10 14 VSS
c12 10 VSS 4.80429e-19 $X=0.513 $Y=0.135
c13 5 VSS 0.00167591f $X=0.513 $Y=0.135
c14 2 VSS 0.0598619f $X=0.513 $Y=0.0675
r15 10 14 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.1535
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AO333X1_ASAP7_75T_L%C1 2 5 7 10 VSS
c11 10 VSS 4.90626e-19 $X=0.5715 $Y=0.0815
c12 5 VSS 0.00223503f $X=0.567 $Y=0.135
c13 2 VSS 0.0638948f $X=0.567 $Y=0.0675
r14 10 13 3.63272 $w=1.8e-08 $l=5.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.0815 $X2=0.567 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
.ends

.subckt PM_AO333X1_ASAP7_75T_L%Y 1 6 9 14 16 18 23 24 30 VSS
c9 30 VSS 0.00559176f $X=0.054 $Y=0.234
c10 28 VSS 0.00317088f $X=0.027 $Y=0.234
c11 24 VSS 0.00568786f $X=0.054 $Y=0.036
c12 23 VSS 0.00654426f $X=0.054 $Y=0.036
c13 21 VSS 0.00317919f $X=0.027 $Y=0.036
c14 20 VSS 4.26553e-19 $X=0.018 $Y=0.216
c15 19 VSS 2.20907e-19 $X=0.018 $Y=0.207
c16 18 VSS 0.0022486f $X=0.018 $Y=0.2
c17 16 VSS 0.00161505f $X=0.018 $Y=0.10125
c18 15 VSS 8.29409e-19 $X=0.018 $Y=0.063
c19 14 VSS 0.00236945f $X=0.0195 $Y=0.1395
c20 12 VSS 4.02856e-19 $X=0.018 $Y=0.225
c21 9 VSS 0.00525308f $X=0.056 $Y=0.2025
c22 6 VSS 2.91692e-19 $X=0.071 $Y=0.2025
c23 1 VSS 2.55988e-19 $X=0.071 $Y=0.0675
r24 28 30 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.054 $Y2=0.234
r25 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r26 21 23 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.054 $Y2=0.036
r27 19 20 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.207 $X2=0.018 $Y2=0.216
r28 18 19 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.207
r29 17 18 3.25926 $w=1.8e-08 $l=4.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.152 $X2=0.018 $Y2=0.2
r30 15 16 2.59722 $w=1.8e-08 $l=3.825e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.10125
r31 14 17 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.152
r32 14 16 2.59722 $w=1.8e-08 $l=3.825e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.10125
r33 12 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r34 12 20 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.216
r35 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r36 11 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r37 9 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r38 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
r39 4 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r40 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./AO333x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO333x1_ASAP7_75t_L  VSS VDD A3 A2 A1 B3 B2 B1 C3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* C3	C3
* B1	B1
* B2	B2
* B3	B3
* A1	A1
* A2	A2
* A3	A3
M0 VSS N_3_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 noxref_16 N_A3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_17 N_A2_M2_g noxref_16 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_3_M3_d N_A1_M3_g noxref_17 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_18 N_B3_M4_g N_3_M4_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_19 N_B2_M5_g noxref_18 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 VSS N_B1_M6_g noxref_19 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_20 N_C3_M7_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 noxref_21 N_C2_M8_g noxref_20 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 N_3_M9_d N_C1_M9_g noxref_21 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M10 VDD N_3_M10_g N_Y_M10_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M11 noxref_14 N_A3_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M12 VDD N_A2_M12_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M13 noxref_14 N_A1_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M14 noxref_15 N_B3_M14_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M15 noxref_14 N_B2_M15_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M16 noxref_15 N_B1_M16_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M17 N_3_M17_d N_C3_M17_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M18 noxref_15 N_C2_M18_g N_3_M18_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
M19 N_3_M19_d N_C1_M19_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
*
* 
* .include "AO333x1_ASAP7_75t_L.pex.sp.AO333X1_ASAP7_75T_L.pxi"
* BEGIN of "./AO333x1_ASAP7_75t_L.pex.sp.AO333X1_ASAP7_75T_L.pxi"
* File: AO333x1_ASAP7_75t_L.pex.sp.AO333X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:08:26 2017
* 
x_PM_AO333X1_ASAP7_75T_L%3 N_3_M0_g N_3_c_2_p N_3_M10_g N_3_M4_s N_3_M3_d
+ N_3_M9_d N_3_M18_s N_3_M17_d N_3_c_38_p N_3_M19_d N_3_c_41_p N_3_c_7_p
+ N_3_c_3_p N_3_c_4_p N_3_c_31_p N_3_c_34_p N_3_c_11_p N_3_c_52_p N_3_c_6_p
+ N_3_c_53_p N_3_c_10_p N_3_c_27_p N_3_c_13_p N_3_c_43_p N_3_c_16_p N_3_c_44_p
+ N_3_c_18_p N_3_c_45_p N_3_c_20_p N_3_c_48_p N_3_c_22_p N_3_c_51_p N_3_c_25_p
+ N_3_c_23_p N_3_c_29_p N_3_c_47_p VSS PM_AO333X1_ASAP7_75T_L%3
x_PM_AO333X1_ASAP7_75T_L%A3 N_A3_M1_g N_A3_c_59_n N_A3_M11_g N_A3_c_60_n A3 VSS
+ PM_AO333X1_ASAP7_75T_L%A3
x_PM_AO333X1_ASAP7_75T_L%A2 N_A2_M2_g N_A2_c_74_n N_A2_M12_g N_A2_c_70_n A2 VSS
+ PM_AO333X1_ASAP7_75T_L%A2
x_PM_AO333X1_ASAP7_75T_L%A1 N_A1_M3_g N_A1_c_88_n N_A1_M13_g A1 VSS
+ PM_AO333X1_ASAP7_75T_L%A1
x_PM_AO333X1_ASAP7_75T_L%B3 N_B3_M4_g N_B3_c_103_n N_B3_M14_g N_B3_c_99_n B3 VSS
+ PM_AO333X1_ASAP7_75T_L%B3
x_PM_AO333X1_ASAP7_75T_L%B2 N_B2_M5_g N_B2_c_115_n N_B2_M15_g B2 VSS
+ PM_AO333X1_ASAP7_75T_L%B2
x_PM_AO333X1_ASAP7_75T_L%B1 N_B1_M6_g N_B1_c_128_n N_B1_M16_g N_B1_c_125_n B1
+ VSS PM_AO333X1_ASAP7_75T_L%B1
x_PM_AO333X1_ASAP7_75T_L%C3 N_C3_M7_g N_C3_c_140_n N_C3_M17_g C3 VSS
+ PM_AO333X1_ASAP7_75T_L%C3
x_PM_AO333X1_ASAP7_75T_L%C2 N_C2_M8_g N_C2_c_153_n N_C2_M18_g N_C2_c_150_n C2
+ VSS PM_AO333X1_ASAP7_75T_L%C2
x_PM_AO333X1_ASAP7_75T_L%C1 N_C1_M9_g N_C1_c_167_n N_C1_M19_g C1 VSS
+ PM_AO333X1_ASAP7_75T_L%C1
x_PM_AO333X1_ASAP7_75T_L%Y N_Y_M0_s N_Y_M10_s N_Y_c_178_p Y N_Y_c_172_n
+ N_Y_c_177_n N_Y_c_173_n N_Y_c_176_n N_Y_c_179_p VSS PM_AO333X1_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M1_g 0.00268443f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_3_c_2_p N_A3_c_59_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_3_c_3_p N_A3_c_60_n 0.00200929f $X=0.081 $Y=0.1205 $X2=0.135 $Y2=0.135
cc_4 N_3_c_4_p N_A3_c_60_n 0.00133324f $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.135
cc_5 N_3_M0_g N_A2_M2_g 2.13359e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 N_3_c_6_p N_A2_M2_g 3.38929e-19 $X=0.198 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_7 N_3_c_7_p N_A2_c_70_n 2.69033e-19 $X=0.081 $Y=0.106 $X2=0.135 $Y2=0.135
cc_8 N_3_c_4_p N_A2_c_70_n 7.10035e-19 $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.135
cc_9 N_3_c_6_p N_A2_c_70_n 0.00123604f $X=0.198 $Y=0.036 $X2=0.135 $Y2=0.135
cc_10 N_3_c_10_p N_A1_M3_g 2.56935e-19 $X=0.252 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_11 N_3_c_11_p A1 0.0013295f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.135
cc_12 N_3_c_10_p A1 0.00123604f $X=0.252 $Y=0.036 $X2=0.135 $Y2=0.135
cc_13 N_3_c_13_p N_B3_M4_g 2.64276e-19 $X=0.306 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_14 N_3_c_11_p N_B3_c_99_n 0.0013295f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.135
cc_15 N_3_c_13_p N_B3_c_99_n 0.00124805f $X=0.306 $Y=0.036 $X2=0.135 $Y2=0.135
cc_16 N_3_c_16_p N_B2_M5_g 3.38929e-19 $X=0.36 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_17 N_3_c_16_p B2 0.00123064f $X=0.36 $Y=0.036 $X2=0.135 $Y2=0.135
cc_18 N_3_c_18_p N_B1_M6_g 2.56935e-19 $X=0.414 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_19 N_3_c_18_p N_B1_c_125_n 0.00123064f $X=0.414 $Y=0.036 $X2=0.135 $Y2=0.135
cc_20 N_3_c_20_p N_C3_M7_g 2.56935e-19 $X=0.468 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_21 N_3_c_20_p C3 0.00123064f $X=0.468 $Y=0.036 $X2=0.135 $Y2=0.135
cc_22 N_3_c_22_p N_C2_M8_g 3.38929e-19 $X=0.522 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_23 N_3_c_23_p N_C2_M8_g 2.38303e-19 $X=0.576 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_24 N_3_c_22_p N_C2_c_150_n 0.00123064f $X=0.522 $Y=0.036 $X2=0.135 $Y2=0.135
cc_25 N_3_c_25_p N_C1_M9_g 2.56935e-19 $X=0.576 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_26 N_3_c_23_p N_C1_M9_g 2.34993e-19 $X=0.576 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_27 N_3_c_27_p C1 0.0013295f $X=0.594 $Y=0.036 $X2=0.135 $Y2=0.135
cc_28 N_3_c_25_p C1 0.00123064f $X=0.576 $Y=0.036 $X2=0.135 $Y2=0.135
cc_29 N_3_c_29_p C1 0.00392202f $X=0.621 $Y=0.164 $X2=0.135 $Y2=0.135
cc_30 N_3_c_3_p Y 0.00141141f $X=0.081 $Y=0.1205 $X2=0.1365 $Y2=0.1485
cc_31 N_3_c_31_p N_Y_c_172_n 0.00141141f $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_32 N_3_M0_g N_Y_c_173_n 2.50002e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_33 N_3_c_31_p N_Y_c_173_n 8.16832e-19 $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_34 N_3_c_34_p N_Y_c_173_n 5.02333e-19 $X=0.144 $Y=0.036 $X2=0 $Y2=0
cc_35 N_3_c_31_p N_Y_c_176_n 0.00143805f $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_36 VSS N_3_c_11_p 0.00107252f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.135
cc_37 VSS N_3_c_23_p 3.07534e-19 $X=0.576 $Y=0.234 $X2=0 $Y2=0
cc_38 VSS N_3_c_38_p 0.00323404f $X=0.486 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_39 VSS N_3_c_23_p 4.49076e-19 $X=0.576 $Y=0.234 $X2=0.135 $Y2=0.135
cc_40 VSS N_3_c_38_p 0.00355395f $X=0.486 $Y=0.2025 $X2=0 $Y2=0
cc_41 VSS N_3_c_41_p 0.00377613f $X=0.592 $Y=0.2025 $X2=0 $Y2=0
cc_42 VSS N_3_c_23_p 0.00250965f $X=0.576 $Y=0.234 $X2=0 $Y2=0
cc_43 VSS N_3_c_43_p 3.02632e-19 $X=0.342 $Y=0.036 $X2=0 $Y2=0
cc_44 VSS N_3_c_44_p 3.02632e-19 $X=0.396 $Y=0.036 $X2=0 $Y2=0
cc_45 VSS N_3_c_45_p 3.02632e-19 $X=0.45 $Y=0.036 $X2=0 $Y2=0
cc_46 VSS N_3_c_41_p 5.59317e-19 $X=0.592 $Y=0.2025 $X2=0 $Y2=0
cc_47 VSS N_3_c_47_p 5.85806e-19 $X=0.621 $Y=0.207 $X2=0 $Y2=0
cc_48 VSS N_3_c_48_p 3.02632e-19 $X=0.504 $Y=0.036 $X2=0 $Y2=0
cc_49 VSS N_3_c_38_p 0.00233206f $X=0.486 $Y=0.2025 $X2=0 $Y2=0
cc_50 VSS N_3_c_23_p 0.00880749f $X=0.576 $Y=0.234 $X2=0 $Y2=0
cc_51 VSS N_3_c_51_p 3.02632e-19 $X=0.558 $Y=0.036 $X2=0 $Y2=0
cc_52 VSS N_3_c_52_p 3.25855e-19 $X=0.18 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_53 VSS N_3_c_53_p 3.56327e-19 $X=0.234 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_54 VSS N_3_c_43_p 3.22747e-19 $X=0.342 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_55 VSS N_3_c_44_p 3.50993e-19 $X=0.396 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_56 VSS N_3_c_48_p 3.3687e-19 $X=0.504 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_57 VSS N_3_c_51_p 3.50993e-19 $X=0.558 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_58 N_A3_M1_g N_A2_M2_g 0.00328721f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_59 N_A3_c_59_n N_A2_c_74_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_60 N_A3_c_60_n N_A2_c_70_n 0.00393501f $X=0.135 $Y=0.135 $X2=0.253 $Y2=0.0675
cc_61 N_A3_M1_g N_A1_M3_g 2.48122e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_62 A3 N_Y_c_177_n 4.38883e-19 $X=0.1365 $Y=0.1485 $X2=0 $Y2=0
cc_63 VSS A3 0.00114532f $X=0.1365 $Y=0.1485 $X2=0.081 $Y2=0.135
cc_64 N_A2_M2_g N_A1_M3_g 0.00312021f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_65 N_A2_c_74_n N_A1_c_88_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_66 N_A2_c_70_n A1 0.00580463f $X=0.189 $Y=0.135 $X2=0.253 $Y2=0.0675
cc_67 N_A2_M2_g N_B3_M4_g 2.53865e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_68 VSS N_A2_c_70_n 0.00114532f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_69 VSS N_A2_M2_g 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0.577 $Y2=0.2025
cc_70 VSS N_A2_c_70_n 0.00125352f $X=0.189 $Y=0.135 $X2=0.577 $Y2=0.2025
cc_71 N_A1_M3_g N_B3_M4_g 0.00353416f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_72 N_A1_c_88_n N_B3_c_103_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_73 A1 N_B3_c_99_n 0.00389755f $X=0.2435 $Y=0.1345 $X2=0.253 $Y2=0.0675
cc_74 N_A1_M3_g N_B2_M5_g 2.88628e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_75 VSS A1 8.74436e-19 $X=0.2435 $Y=0.1345 $X2=0.253 $Y2=0.0675
cc_76 VSS N_A1_M3_g 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_77 VSS A1 0.00125352f $X=0.2435 $Y=0.1345 $X2=0 $Y2=0
cc_78 VSS A1 2.64861e-19 $X=0.2435 $Y=0.1345 $X2=0.486 $Y2=0.2025
cc_79 N_B3_M4_g N_B2_M5_g 0.00355599f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_80 N_B3_c_103_n N_B2_c_115_n 9.06722e-19 $X=0.297 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_81 N_B3_c_99_n B2 0.00483098f $X=0.297 $Y=0.135 $X2=0.253 $Y2=0.0675
cc_82 N_B3_M4_g N_B1_M6_g 2.88628e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_83 VSS N_B3_M4_g 3.57119e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_84 VSS N_B3_c_99_n 5.37372e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_85 N_B2_M5_g N_B1_M6_g 0.00353416f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_86 N_B2_c_115_n N_B1_c_128_n 9.07977e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_87 B2 N_B1_c_125_n 0.00483098f $X=0.3505 $Y=0.0845 $X2=0.253 $Y2=0.0675
cc_88 N_B2_M5_g N_C3_M7_g 2.53865e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_89 VSS N_B2_M5_g 2.08515e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_90 VSS N_B2_M5_g 2.76185e-19 $X=0.351 $Y=0.0675 $X2=0.577 $Y2=0.2025
cc_91 VSS B2 0.0012322f $X=0.3505 $Y=0.0845 $X2=0.577 $Y2=0.2025
cc_92 N_B1_M6_g N_C3_M7_g 0.00317103f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_93 N_B1_c_128_n N_C3_c_140_n 9.07977e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_94 N_B1_c_125_n C3 0.0040634f $X=0.405 $Y=0.135 $X2=0.253 $Y2=0.0675
cc_95 N_B1_M6_g N_C2_M8_g 2.53865e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_96 VSS N_B1_M6_g 3.51973e-19 $X=0.405 $Y=0.0675 $X2=0.592 $Y2=0.2025
cc_97 VSS N_B1_c_125_n 0.00121543f $X=0.405 $Y=0.135 $X2=0.592 $Y2=0.2025
cc_98 N_C3_M7_g N_C2_M8_g 0.00353416f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_99 N_C3_c_140_n N_C2_c_153_n 9.07977e-19 $X=0.459 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_100 C3 N_C2_c_150_n 0.00483098f $X=0.4565 $Y=0.0835 $X2=0.253 $Y2=0.0675
cc_101 N_C3_M7_g N_C1_M9_g 2.88628e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_102 VSS N_C3_M7_g 3.62029e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.106
cc_103 VSS C3 0.0012322f $X=0.4565 $Y=0.0835 $X2=0.081 $Y2=0.106
cc_104 N_C2_M8_g N_C1_M9_g 0.00360681f $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_105 N_C2_c_153_n N_C1_c_167_n 9.55934e-19 $X=0.513 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_106 N_C2_c_150_n C1 0.00482806f $X=0.513 $Y=0.135 $X2=0.253 $Y2=0.0675
cc_107 VSS N_C2_M8_g 2.68514e-19 $X=0.513 $Y=0.0675 $X2=0.126 $Y2=0.072
cc_108 VSS N_C2_c_150_n 0.00121543f $X=0.513 $Y=0.135 $X2=0.126 $Y2=0.072
cc_109 VSS N_C1_M9_g 2.83408e-19 $X=0.567 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_110 VSS C1 0.00147374f $X=0.5715 $Y=0.0815 $X2=0.081 $Y2=0.135
cc_111 VSS N_Y_c_178_p 2.2337e-19 $X=0.056 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_112 VSS N_Y_c_179_p 2.83875e-19 $X=0.054 $Y=0.234 $X2=0.486 $Y2=0.2025

* END of "./AO333x1_ASAP7_75t_L.pex.sp.AO333X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO333x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:08:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO333x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO333x2_ASAP7_75t_L.pex.sp.pex"
* File: AO333x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:08:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO333X2_ASAP7_75T_L%3 2 7 10 13 15 17 18 22 27 28 31 32 35 42 43 46
+ 47 49 52 54 56 57 58 59 63 65 67 68 69 70 71 72 73 74 75 76 86 91 93 VSS
c64 93 VSS 6.70384e-19 $X=0.675 $Y=0.207
c65 92 VSS 0.00104083f $X=0.675 $Y=0.189
c66 91 VSS 0.00414971f $X=0.675 $Y=0.164
c67 90 VSS 9.77725e-19 $X=0.675 $Y=0.07
c68 89 VSS 8.85605e-19 $X=0.675 $Y=0.225
c69 87 VSS 8.42643e-19 $X=0.639 $Y=0.234
c70 86 VSS 0.00886015f $X=0.63 $Y=0.234
c71 78 VSS 0.00618523f $X=0.666 $Y=0.234
c72 77 VSS 8.42643e-19 $X=0.639 $Y=0.036
c73 76 VSS 0.00142296f $X=0.63 $Y=0.036
c74 75 VSS 0.00346807f $X=0.612 $Y=0.036
c75 74 VSS 0.00142296f $X=0.576 $Y=0.036
c76 73 VSS 0.00330791f $X=0.558 $Y=0.036
c77 72 VSS 0.00142296f $X=0.522 $Y=0.036
c78 71 VSS 0.0068014f $X=0.504 $Y=0.036
c79 70 VSS 0.00142296f $X=0.468 $Y=0.036
c80 69 VSS 0.00346807f $X=0.45 $Y=0.036
c81 68 VSS 0.00142296f $X=0.414 $Y=0.036
c82 67 VSS 0.00309345f $X=0.396 $Y=0.036
c83 66 VSS 3.54965e-19 $X=0.364 $Y=0.036
c84 65 VSS 0.00146362f $X=0.36 $Y=0.036
c85 64 VSS 0.00274772f $X=0.342 $Y=0.036
c86 63 VSS 0.00224055f $X=0.648 $Y=0.036
c87 60 VSS 0.00106066f $X=0.315 $Y=0.036
c88 59 VSS 0.00142296f $X=0.306 $Y=0.036
c89 58 VSS 0.00376615f $X=0.288 $Y=0.036
c90 57 VSS 0.00142296f $X=0.252 $Y=0.036
c91 56 VSS 0.00329341f $X=0.234 $Y=0.036
c92 55 VSS 3.78291e-19 $X=0.202 $Y=0.036
c93 54 VSS 0.00146362f $X=0.198 $Y=0.036
c94 53 VSS 0.00294815f $X=0.18 $Y=0.036
c95 52 VSS 0.00218387f $X=0.324 $Y=0.036
c96 49 VSS 0.00270205f $X=0.162 $Y=0.036
c97 48 VSS 0.00607741f $X=0.666 $Y=0.036
c98 47 VSS 7.02432e-19 $X=0.153 $Y=0.099
c99 46 VSS 0.00127834f $X=0.153 $Y=0.07
c100 45 VSS 9.44693e-19 $X=0.153 $Y=0.126
c101 43 VSS 4.68643e-20 $X=0.122 $Y=0.135
c102 42 VSS 3.04954e-19 $X=0.117 $Y=0.135
c103 37 VSS 0.00151949f $X=0.144 $Y=0.135
c104 35 VSS 0.00257027f $X=0.646 $Y=0.2025
c105 31 VSS 0.00238723f $X=0.54 $Y=0.2025
c106 27 VSS 7.12337e-19 $X=0.557 $Y=0.2025
c107 25 VSS 2.69461e-19 $X=0.646 $Y=0.0675
c108 17 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c109 13 VSS 0.00520739f $X=0.135 $Y=0.135
c110 10 VSS 0.0590374f $X=0.135 $Y=0.0675
c111 2 VSS 0.0615998f $X=0.081 $Y=0.0675
r112 92 93 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.189 $X2=0.675 $Y2=0.207
r113 91 92 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.164 $X2=0.675 $Y2=0.189
r114 90 91 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.07 $X2=0.675 $Y2=0.164
r115 89 93 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.225 $X2=0.675 $Y2=0.207
r116 88 90 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.045 $X2=0.675 $Y2=0.07
r117 86 87 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.234 $X2=0.639 $Y2=0.234
r118 84 87 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.639 $Y2=0.234
r119 80 86 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.63 $Y2=0.234
r120 78 89 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.234 $X2=0.675 $Y2=0.225
r121 78 84 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.234 $X2=0.648 $Y2=0.234
r122 76 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.036 $X2=0.639 $Y2=0.036
r123 75 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.63 $Y2=0.036
r124 74 75 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.036 $X2=0.612 $Y2=0.036
r125 73 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.576 $Y2=0.036
r126 72 73 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.558 $Y2=0.036
r127 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.522 $Y2=0.036
r128 70 71 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.504 $Y2=0.036
r129 69 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r130 68 69 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.45 $Y2=0.036
r131 67 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r132 66 67 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.364
+ $Y=0.036 $X2=0.396 $Y2=0.036
r133 65 66 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.364 $Y2=0.036
r134 64 65 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r135 62 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.639 $Y2=0.036
r136 62 63 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r137 59 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.315 $Y2=0.036
r138 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r139 57 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r140 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r141 55 56 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.036 $X2=0.234 $Y2=0.036
r142 54 55 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.202 $Y2=0.036
r143 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r144 51 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r145 51 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.315 $Y2=0.036
r146 51 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r147 49 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r148 48 88 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.036 $X2=0.675 $Y2=0.045
r149 48 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.648 $Y2=0.036
r150 46 47 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.07 $X2=0.153 $Y2=0.099
r151 45 47 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.126 $X2=0.153 $Y2=0.099
r152 44 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.153 $Y=0.045 $X2=0.162 $Y2=0.036
r153 44 46 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.045 $X2=0.153 $Y2=0.07
r154 42 43 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.135 $X2=0.122 $Y2=0.135
r155 39 42 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.117 $Y2=0.135
r156 37 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.144 $Y=0.135 $X2=0.153 $Y2=0.126
r157 37 43 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.122 $Y2=0.135
r158 35 84 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234
+ $X2=0.648 $Y2=0.234
r159 32 35 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.646 $Y2=0.2025
r160 31 80 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r161 28 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r162 27 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r163 25 63 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r164 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.646 $Y2=0.0675
r165 21 52 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r166 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r167 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r168 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r169 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r170 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r171 5 39 3.03549 $a=6.48e-16 $layer=V0LIG $count=2 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r172 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r173 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AO333X2_ASAP7_75T_L%A3 2 5 7 10 13 VSS
c12 13 VSS 0.0025565f $X=0.189 $Y=0.135
c13 10 VSS 3.18228e-19 $X=0.1875 $Y=0.0925
c14 5 VSS 0.00116428f $X=0.189 $Y=0.135
c15 2 VSS 0.0561685f $X=0.189 $Y=0.0675
r16 10 13 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.0925 $X2=0.189 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO333X2_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c13 10 VSS 0.00154873f $X=0.243 $Y=0.135
c14 5 VSS 0.00106612f $X=0.243 $Y=0.135
c15 2 VSS 0.057046f $X=0.243 $Y=0.0675
r16 10 14 3.49691 $w=1.8e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.1865
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO333X2_ASAP7_75T_L%A1 2 5 7 10 VSS
c15 10 VSS 0.00153576f $X=0.2975 $Y=0.1345
c16 5 VSS 0.00110983f $X=0.297 $Y=0.135
c17 2 VSS 0.058107f $X=0.297 $Y=0.0675
r18 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r19 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r20 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO333X2_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c13 10 VSS 5.11375e-19 $X=0.351 $Y=0.135
c14 5 VSS 0.0011055f $X=0.351 $Y=0.135
c15 2 VSS 0.0591416f $X=0.351 $Y=0.0675
r16 10 14 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.1545
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AO333X2_ASAP7_75T_L%B2 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.4045 $Y=0.0845
c14 5 VSS 0.00164678f $X=0.405 $Y=0.135
c15 2 VSS 0.0591416f $X=0.405 $Y=0.0675
r16 10 13 3.42901 $w=1.8e-08 $l=5.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.0845 $X2=0.405 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO333X2_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c12 10 VSS 6.96915e-19 $X=0.459 $Y=0.135
c13 5 VSS 0.00164704f $X=0.459 $Y=0.135
c14 2 VSS 0.0594389f $X=0.459 $Y=0.0675
r15 10 14 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.1555
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AO333X2_ASAP7_75T_L%C3 2 5 7 10 VSS
c12 10 VSS 6.96915e-19 $X=0.5105 $Y=0.0835
c13 5 VSS 0.00160703f $X=0.513 $Y=0.135
c14 2 VSS 0.0592509f $X=0.513 $Y=0.0675
r15 10 13 3.49691 $w=1.8e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.0835 $X2=0.513 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AO333X2_ASAP7_75T_L%C2 2 5 7 10 14 VSS
c12 10 VSS 4.80429e-19 $X=0.567 $Y=0.135
c13 5 VSS 0.00167591f $X=0.567 $Y=0.135
c14 2 VSS 0.0598619f $X=0.567 $Y=0.0675
r15 10 14 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.1535
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
.ends

.subckt PM_AO333X2_ASAP7_75T_L%C1 2 5 7 10 VSS
c11 10 VSS 4.90626e-19 $X=0.6255 $Y=0.0815
c12 5 VSS 0.00223503f $X=0.621 $Y=0.135
c13 2 VSS 0.0638948f $X=0.621 $Y=0.0675
r14 10 13 3.63272 $w=1.8e-08 $l=5.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.0815 $X2=0.621 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
.ends

.subckt PM_AO333X2_ASAP7_75T_L%Y 1 2 5 6 7 10 14 16 18 19 25 28 35 VSS
c16 35 VSS 0.00511303f $X=0.108 $Y=0.072
c17 28 VSS 0.00187096f $X=0.0875 $Y=0.234
c18 27 VSS 0.00712235f $X=0.067 $Y=0.234
c19 25 VSS 0.00373949f $X=0.108 $Y=0.234
c20 23 VSS 0.00319268f $X=0.027 $Y=0.234
c21 22 VSS 7.10506e-19 $X=0.067 $Y=0.09
c22 21 VSS 0.00398742f $X=0.062 $Y=0.09
c23 20 VSS 0.00151603f $X=0.027 $Y=0.09
c24 19 VSS 4.07525e-19 $X=0.099 $Y=0.09
c25 18 VSS 0.00325596f $X=0.018 $Y=0.2
c26 16 VSS 2.72708e-19 $X=0.018 $Y=0.13275
c27 15 VSS 0.00146526f $X=0.018 $Y=0.126
c28 14 VSS 4.40771e-19 $X=0.0195 $Y=0.1395
c29 12 VSS 0.00126561f $X=0.018 $Y=0.225
c30 10 VSS 0.00902046f $X=0.108 $Y=0.2025
c31 6 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c32 5 VSS 0.00861358f $X=0.108 $Y=0.0675
c33 1 VSS 6.59976e-19 $X=0.125 $Y=0.0675
r34 33 35 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.081 $X2=0.108 $Y2=0.072
r35 27 28 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.067
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r36 25 28 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r37 23 27 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.067 $Y2=0.234
r38 21 22 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.062
+ $Y=0.09 $X2=0.067 $Y2=0.09
r39 20 21 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.09 $X2=0.062 $Y2=0.09
r40 19 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.099 $Y=0.09 $X2=0.108 $Y2=0.081
r41 19 22 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.09 $X2=0.067 $Y2=0.09
r42 17 18 3.80247 $w=1.8e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.2
r43 15 16 0.458333 $w=1.8e-08 $l=6.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.13275
r44 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.144
r45 14 16 0.458333 $w=1.8e-08 $l=6.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.13275
r46 12 23 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r47 12 18 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2
r48 11 20 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.099 $X2=0.027 $Y2=0.09
r49 11 15 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.099 $X2=0.018 $Y2=0.126
r50 10 25 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r51 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r52 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r53 5 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072 $X2=0.108
+ $Y2=0.072
r54 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r55 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./AO333x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO333x2_ASAP7_75t_L  VSS VDD A3 A2 A1 B3 B2 B1 C3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* C3	C3
* B1	B1
* B2	B2
* B3	B3
* A1	A1
* A2	A2
* A3	A3
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_16 N_A3_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_17 N_A2_M3_g noxref_16 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_3_M4_d N_A1_M4_g noxref_17 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_18 N_B3_M5_g N_3_M5_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_19 N_B2_M6_g noxref_18 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 VSS N_B1_M7_g noxref_19 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 noxref_20 N_C3_M8_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 noxref_21 N_C2_M9_g noxref_20 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M10 N_3_M10_d N_C1_M10_g noxref_21 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.611 $Y=0.027
M11 N_Y_M11_d N_3_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M12 N_Y_M12_d N_3_M12_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M13 noxref_14 N_A3_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M14 VDD N_A2_M14_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M15 noxref_14 N_A1_M15_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M16 noxref_15 N_B3_M16_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M17 noxref_14 N_B2_M17_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M18 noxref_15 N_B1_M18_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M19 N_3_M19_d N_C3_M19_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
M20 noxref_15 N_C2_M20_g N_3_M20_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M21 N_3_M21_d N_C1_M21_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.611 $Y=0.162
*
* 
* .include "AO333x2_ASAP7_75t_L.pex.sp.AO333X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO333x2_ASAP7_75t_L.pex.sp.AO333X2_ASAP7_75T_L.pxi"
* File: AO333x2_ASAP7_75t_L.pex.sp.AO333X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:08:48 2017
* 
x_PM_AO333X2_ASAP7_75T_L%3 N_3_M0_g N_3_M11_g N_3_M1_g N_3_c_4_p N_3_M12_g
+ N_3_M5_s N_3_M4_d N_3_M10_d N_3_M20_s N_3_M19_d N_3_c_45_p N_3_M21_d
+ N_3_c_48_p N_3_c_34_p N_3_c_37_p N_3_c_41_p N_3_c_5_p N_3_c_31_p N_3_c_11_p
+ N_3_c_3_p N_3_c_59_p N_3_c_8_p N_3_c_60_p N_3_c_10_p N_3_c_27_p N_3_c_13_p
+ N_3_c_50_p N_3_c_16_p N_3_c_51_p N_3_c_18_p N_3_c_52_p N_3_c_20_p N_3_c_55_p
+ N_3_c_22_p N_3_c_58_p N_3_c_25_p N_3_c_23_p N_3_c_29_p N_3_c_54_p VSS
+ PM_AO333X2_ASAP7_75T_L%3
x_PM_AO333X2_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_68_n N_A3_M13_g A3 N_A3_c_75_p VSS
+ PM_AO333X2_ASAP7_75T_L%A3
x_PM_AO333X2_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_81_n N_A2_M14_g N_A2_c_79_n A2 VSS
+ PM_AO333X2_ASAP7_75T_L%A2
x_PM_AO333X2_ASAP7_75T_L%A1 N_A1_M4_g N_A1_c_95_n N_A1_M15_g A1 VSS
+ PM_AO333X2_ASAP7_75T_L%A1
x_PM_AO333X2_ASAP7_75T_L%B3 N_B3_M5_g N_B3_c_110_n N_B3_M16_g N_B3_c_106_n B3
+ VSS PM_AO333X2_ASAP7_75T_L%B3
x_PM_AO333X2_ASAP7_75T_L%B2 N_B2_M6_g N_B2_c_122_n N_B2_M17_g B2 VSS
+ PM_AO333X2_ASAP7_75T_L%B2
x_PM_AO333X2_ASAP7_75T_L%B1 N_B1_M7_g N_B1_c_135_n N_B1_M18_g N_B1_c_132_n B1
+ VSS PM_AO333X2_ASAP7_75T_L%B1
x_PM_AO333X2_ASAP7_75T_L%C3 N_C3_M8_g N_C3_c_147_n N_C3_M19_g C3 VSS
+ PM_AO333X2_ASAP7_75T_L%C3
x_PM_AO333X2_ASAP7_75T_L%C2 N_C2_M9_g N_C2_c_160_n N_C2_M20_g N_C2_c_157_n C2
+ VSS PM_AO333X2_ASAP7_75T_L%C2
x_PM_AO333X2_ASAP7_75T_L%C1 N_C1_M10_g N_C1_c_174_n N_C1_M21_g C1 VSS
+ PM_AO333X2_ASAP7_75T_L%C1
x_PM_AO333X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_c_179_n N_Y_M12_d N_Y_M11_d
+ N_Y_c_192_p Y N_Y_c_181_n N_Y_c_191_n N_Y_c_183_n N_Y_c_185_n N_Y_c_186_n
+ N_Y_c_188_n VSS PM_AO333X2_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M2_g 2.13359e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_A3_M2_g 0.00268443f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_A3_M2_g 2.64276e-19 $X=0.198 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_4 N_3_c_4_p N_A3_c_68_n 0.00111166f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_5 N_3_c_5_p A3 0.00614289f $X=0.153 $Y=0.099 $X2=0.1875 $Y2=0.0925
cc_6 N_3_c_3_p A3 0.00125352f $X=0.198 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_7 N_3_M1_g N_A2_M3_g 2.13359e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_8 N_3_c_8_p N_A2_M3_g 3.38929e-19 $X=0.252 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_9 N_3_c_8_p N_A2_c_79_n 0.00123604f $X=0.252 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_10 N_3_c_10_p N_A1_M4_g 2.56935e-19 $X=0.306 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_11 N_3_c_11_p A1 0.0013295f $X=0.324 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_12 N_3_c_10_p A1 0.00123604f $X=0.306 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_13 N_3_c_13_p N_B3_M5_g 2.64276e-19 $X=0.36 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_14 N_3_c_11_p N_B3_c_106_n 0.0013295f $X=0.324 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_15 N_3_c_13_p N_B3_c_106_n 0.00124805f $X=0.36 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_16 N_3_c_16_p N_B2_M6_g 3.38929e-19 $X=0.414 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_17 N_3_c_16_p B2 0.00123064f $X=0.414 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_18 N_3_c_18_p N_B1_M7_g 2.56935e-19 $X=0.468 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_19 N_3_c_18_p N_B1_c_132_n 0.00123064f $X=0.468 $Y=0.036 $X2=0.1875
+ $Y2=0.0925
cc_20 N_3_c_20_p N_C3_M8_g 2.56935e-19 $X=0.522 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_21 N_3_c_20_p C3 0.00123064f $X=0.522 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_22 N_3_c_22_p N_C2_M9_g 3.38929e-19 $X=0.576 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_23 N_3_c_23_p N_C2_M9_g 2.38303e-19 $X=0.63 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_24 N_3_c_22_p N_C2_c_157_n 0.00123064f $X=0.576 $Y=0.036 $X2=0.1875
+ $Y2=0.0925
cc_25 N_3_c_25_p N_C1_M10_g 2.56935e-19 $X=0.63 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_26 N_3_c_23_p N_C1_M10_g 2.34993e-19 $X=0.63 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_27 N_3_c_27_p C1 0.0013295f $X=0.648 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_28 N_3_c_25_p C1 0.00123064f $X=0.63 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_29 N_3_c_29_p C1 0.00392202f $X=0.675 $Y=0.164 $X2=0.1875 $Y2=0.0925
cc_30 N_3_c_4_p N_Y_M1_d 4.01556e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_31 N_3_c_31_p N_Y_c_179_n 0.00112295f $X=0.162 $Y=0.036 $X2=0.189 $Y2=0.135
cc_32 N_3_c_4_p N_Y_M12_d 3.80218e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_33 N_3_c_4_p N_Y_c_181_n 4.17004e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_34 N_3_c_34_p N_Y_c_181_n 8.21717e-19 $X=0.117 $Y=0.135 $X2=0 $Y2=0
cc_35 N_3_M0_g N_Y_c_183_n 2.50197e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_3_c_34_p N_Y_c_183_n 0.00246923f $X=0.117 $Y=0.135 $X2=0 $Y2=0
cc_37 N_3_c_37_p N_Y_c_185_n 4.13141e-19 $X=0.122 $Y=0.135 $X2=0 $Y2=0
cc_38 N_3_M0_g N_Y_c_186_n 3.32206e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_3_c_34_p N_Y_c_186_n 4.13141e-19 $X=0.117 $Y=0.135 $X2=0 $Y2=0
cc_40 N_3_M0_g N_Y_c_188_n 2.87828e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_41 N_3_c_41_p N_Y_c_188_n 0.00159053f $X=0.153 $Y=0.07 $X2=0 $Y2=0
cc_42 N_3_c_5_p N_Y_c_188_n 0.00159053f $X=0.153 $Y=0.099 $X2=0 $Y2=0
cc_43 VSS N_3_c_11_p 0.00107252f $X=0.324 $Y=0.036 $X2=0.1875 $Y2=0.0925
cc_44 VSS N_3_c_23_p 3.07534e-19 $X=0.63 $Y=0.234 $X2=0 $Y2=0
cc_45 VSS N_3_c_45_p 0.00323404f $X=0.54 $Y=0.2025 $X2=0.1875 $Y2=0.0925
cc_46 VSS N_3_c_23_p 4.49076e-19 $X=0.63 $Y=0.234 $X2=0.1875 $Y2=0.0925
cc_47 VSS N_3_c_45_p 0.00355395f $X=0.54 $Y=0.2025 $X2=0 $Y2=0
cc_48 VSS N_3_c_48_p 0.00377613f $X=0.646 $Y=0.2025 $X2=0 $Y2=0
cc_49 VSS N_3_c_23_p 0.00250965f $X=0.63 $Y=0.234 $X2=0 $Y2=0
cc_50 VSS N_3_c_50_p 3.02632e-19 $X=0.396 $Y=0.036 $X2=0 $Y2=0
cc_51 VSS N_3_c_51_p 3.02632e-19 $X=0.45 $Y=0.036 $X2=0 $Y2=0
cc_52 VSS N_3_c_52_p 3.02632e-19 $X=0.504 $Y=0.036 $X2=0 $Y2=0
cc_53 VSS N_3_c_48_p 5.59317e-19 $X=0.646 $Y=0.2025 $X2=0 $Y2=0
cc_54 VSS N_3_c_54_p 5.85806e-19 $X=0.675 $Y=0.207 $X2=0 $Y2=0
cc_55 VSS N_3_c_55_p 3.02632e-19 $X=0.558 $Y=0.036 $X2=0 $Y2=0
cc_56 VSS N_3_c_45_p 0.00233206f $X=0.54 $Y=0.2025 $X2=0 $Y2=0
cc_57 VSS N_3_c_23_p 0.00880749f $X=0.63 $Y=0.234 $X2=0 $Y2=0
cc_58 VSS N_3_c_58_p 3.02632e-19 $X=0.612 $Y=0.036 $X2=0 $Y2=0
cc_59 VSS N_3_c_59_p 3.25855e-19 $X=0.234 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_60 VSS N_3_c_60_p 3.56327e-19 $X=0.288 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_61 VSS N_3_c_50_p 3.22747e-19 $X=0.396 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_62 VSS N_3_c_51_p 3.50993e-19 $X=0.45 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_63 VSS N_3_c_55_p 3.3687e-19 $X=0.558 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_64 VSS N_3_c_58_p 3.50993e-19 $X=0.612 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_65 N_A3_M2_g N_A2_M3_g 0.00328721f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_66 N_A3_c_68_n N_A2_c_81_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_67 A3 N_A2_c_79_n 0.00582603f $X=0.1875 $Y=0.0925 $X2=0.135 $Y2=0.0675
cc_68 N_A3_M2_g N_A1_M4_g 2.48122e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_69 N_A3_c_75_p N_Y_c_191_n 2.88614e-19 $X=0.189 $Y=0.135 $X2=0.307 $Y2=0.0675
cc_70 VSS N_A3_c_75_p 0.00114532f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_71 N_A2_M3_g N_A1_M4_g 0.00312021f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_72 N_A2_c_81_n N_A1_c_95_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_73 N_A2_c_79_n A1 0.00581998f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_74 N_A2_M3_g N_B3_M5_g 2.53865e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_75 VSS N_A2_c_79_n 0.00114532f $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_76 VSS N_A2_M3_g 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_77 VSS N_A2_c_79_n 0.00125352f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_78 N_A1_M4_g N_B3_M5_g 0.00353416f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_79 N_A1_c_95_n N_B3_c_110_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_80 A1 N_B3_c_106_n 0.00389755f $X=0.2975 $Y=0.1345 $X2=0.135 $Y2=0.0675
cc_81 N_A1_M4_g N_B2_M6_g 2.88628e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_82 VSS A1 8.74436e-19 $X=0.2975 $Y=0.1345 $X2=0.135 $Y2=0.0675
cc_83 VSS N_A1_M4_g 2.64276e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_84 VSS A1 0.00125352f $X=0.2975 $Y=0.1345 $X2=0 $Y2=0
cc_85 VSS A1 2.64861e-19 $X=0.2975 $Y=0.1345 $X2=0.646 $Y2=0.0675
cc_86 N_B3_M5_g N_B2_M6_g 0.00355599f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_87 N_B3_c_110_n N_B2_c_122_n 9.06722e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_88 N_B3_c_106_n B2 0.00483098f $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_89 N_B3_M5_g N_B1_M7_g 2.88628e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_90 VSS N_B3_M5_g 3.57119e-19 $X=0.351 $Y=0.0675 $X2=0.54 $Y2=0.2025
cc_91 VSS N_B3_c_106_n 5.37372e-19 $X=0.351 $Y=0.135 $X2=0.54 $Y2=0.2025
cc_92 N_B2_M6_g N_B1_M7_g 0.00353416f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_93 N_B2_c_122_n N_B1_c_135_n 9.07977e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_94 B2 N_B1_c_132_n 0.00483098f $X=0.4045 $Y=0.0845 $X2=0.135 $Y2=0.0675
cc_95 N_B2_M6_g N_C3_M8_g 2.53865e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_96 VSS N_B2_M6_g 2.08515e-19 $X=0.405 $Y=0.0675 $X2=0.523 $Y2=0.2025
cc_97 VSS N_B2_M6_g 2.76185e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_98 VSS B2 0.0012322f $X=0.4045 $Y=0.0845 $X2=0 $Y2=0
cc_99 N_B1_M7_g N_C3_M8_g 0.00317103f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_100 N_B1_c_135_n N_C3_c_147_n 9.07977e-19 $X=0.459 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_101 N_B1_c_132_n C3 0.0040634f $X=0.459 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_102 N_B1_M7_g N_C2_M9_g 2.53865e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_103 VSS N_B1_M7_g 3.51973e-19 $X=0.459 $Y=0.0675 $X2=0.557 $Y2=0.2025
cc_104 VSS N_B1_c_132_n 0.00121543f $X=0.459 $Y=0.135 $X2=0.557 $Y2=0.2025
cc_105 N_C3_M8_g N_C2_M9_g 0.00353416f $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_106 N_C3_c_147_n N_C2_c_160_n 9.07977e-19 $X=0.513 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_107 C3 N_C2_c_157_n 0.00483098f $X=0.5105 $Y=0.0835 $X2=0.135 $Y2=0.0675
cc_108 N_C3_M8_g N_C1_M10_g 2.88628e-19 $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_109 VSS N_C3_M8_g 3.62029e-19 $X=0.513 $Y=0.0675 $X2=0.646 $Y2=0.2025
cc_110 VSS C3 0.0012322f $X=0.5105 $Y=0.0835 $X2=0.646 $Y2=0.2025
cc_111 N_C2_M9_g N_C1_M10_g 0.00360681f $X=0.567 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_112 N_C2_c_160_n N_C1_c_174_n 9.55934e-19 $X=0.567 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_113 N_C2_c_157_n C1 0.00482806f $X=0.567 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_114 VSS N_C2_M9_g 2.68514e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_115 VSS N_C2_c_157_n 0.00121543f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_116 VSS N_C1_M10_g 2.83408e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_117 VSS C1 0.00147374f $X=0.6255 $Y=0.0815 $X2=0 $Y2=0
cc_118 VSS N_Y_c_192_p 2.23372e-19 $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_119 VSS N_Y_c_185_n 2.92971e-19 $X=0.108 $Y=0.234 $X2=0.646 $Y2=0.0675

* END of "./AO333x2_ASAP7_75t_L.pex.sp.AO333X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AO33x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:09:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AO33x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AO33x2_ASAP7_75t_L.pex.sp.pex"
* File: AO33x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:09:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AO33X2_ASAP7_75T_L%3 2 7 10 13 15 17 18 22 23 26 27 30 37 38 40 41 42
+ 44 47 49 51 52 53 54 55 57 59 60 61 62 72 73 74 76 81 VSS
c57 81 VSS 0.00433728f $X=0.513 $Y=0.164
c58 80 VSS 0.0011536f $X=0.513 $Y=0.07
c59 79 VSS 0.00114086f $X=0.513 $Y=0.189
c60 77 VSS 4.44014e-19 $X=0.477 $Y=0.198
c61 76 VSS 5.17397e-19 $X=0.468 $Y=0.198
c62 75 VSS 3.76924e-20 $X=0.45 $Y=0.198
c63 74 VSS 4.61151e-19 $X=0.449 $Y=0.198
c64 73 VSS 8.46035e-21 $X=0.414 $Y=0.198
c65 72 VSS 6.53455e-19 $X=0.396 $Y=0.198
c66 64 VSS 0.00364529f $X=0.504 $Y=0.198
c67 63 VSS 0.00338644f $X=0.486 $Y=0.036
c68 62 VSS 0.00142296f $X=0.468 $Y=0.036
c69 61 VSS 0.00344621f $X=0.45 $Y=0.036
c70 60 VSS 0.00142296f $X=0.414 $Y=0.036
c71 59 VSS 0.00320368f $X=0.396 $Y=0.036
c72 57 VSS 0.00146362f $X=0.36 $Y=0.036
c73 56 VSS 0.00258409f $X=0.342 $Y=0.036
c74 55 VSS 8.97023e-19 $X=0.315 $Y=0.036
c75 54 VSS 0.00142296f $X=0.306 $Y=0.036
c76 53 VSS 0.00360252f $X=0.288 $Y=0.036
c77 52 VSS 0.00142296f $X=0.252 $Y=0.036
c78 51 VSS 0.0034188f $X=0.234 $Y=0.036
c79 49 VSS 0.00146362f $X=0.198 $Y=0.036
c80 48 VSS 0.00294815f $X=0.18 $Y=0.036
c81 47 VSS 0.00218387f $X=0.324 $Y=0.036
c82 44 VSS 0.00270205f $X=0.162 $Y=0.036
c83 43 VSS 0.00579233f $X=0.504 $Y=0.036
c84 42 VSS 2.58269e-19 $X=0.153 $Y=0.081
c85 41 VSS 0.00127834f $X=0.153 $Y=0.07
c86 40 VSS 0.00121245f $X=0.153 $Y=0.126
c87 38 VSS 4.68643e-20 $X=0.122 $Y=0.135
c88 37 VSS 3.0544e-19 $X=0.117 $Y=0.135
c89 32 VSS 0.00151949f $X=0.144 $Y=0.135
c90 30 VSS 0.00307504f $X=0.484 $Y=0.216
c91 26 VSS 0.00272791f $X=0.378 $Y=0.216
c92 22 VSS 5.85232e-19 $X=0.395 $Y=0.216
c93 17 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c94 13 VSS 0.00533596f $X=0.135 $Y=0.1345
c95 10 VSS 0.06188f $X=0.135 $Y=0.0675
c96 2 VSS 0.0645473f $X=0.081 $Y=0.0675
r97 80 81 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.07 $X2=0.513 $Y2=0.164
r98 79 81 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.513 $Y2=0.164
r99 78 80 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.07
r100 76 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.198 $X2=0.477 $Y2=0.198
r101 75 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.198 $X2=0.468 $Y2=0.198
r102 74 75 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.449
+ $Y=0.198 $X2=0.45 $Y2=0.198
r103 73 74 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.449 $Y2=0.198
r104 72 73 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.414 $Y2=0.198
r105 70 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.198 $X2=0.477 $Y2=0.198
r106 66 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.198 $X2=0.396 $Y2=0.198
r107 64 79 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.198 $X2=0.513 $Y2=0.189
r108 64 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.198 $X2=0.486 $Y2=0.198
r109 62 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.486 $Y2=0.036
r110 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r111 60 61 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.45 $Y2=0.036
r112 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r113 58 59 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.361
+ $Y=0.036 $X2=0.396 $Y2=0.036
r114 57 58 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.361 $Y2=0.036
r115 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r116 54 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.315 $Y2=0.036
r117 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r118 52 53 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r119 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r120 50 51 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.199
+ $Y=0.036 $X2=0.234 $Y2=0.036
r121 49 50 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.199 $Y2=0.036
r122 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r123 46 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r124 46 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.315 $Y2=0.036
r125 46 47 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r126 44 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r127 43 78 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.036 $X2=0.513 $Y2=0.045
r128 43 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.486 $Y2=0.036
r129 41 42 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.07 $X2=0.153 $Y2=0.081
r130 40 42 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.126 $X2=0.153 $Y2=0.081
r131 39 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.153 $Y=0.045 $X2=0.162 $Y2=0.036
r132 39 41 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.045 $X2=0.153 $Y2=0.07
r133 37 38 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.135 $X2=0.122 $Y2=0.135
r134 34 37 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.117 $Y2=0.135
r135 32 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.144 $Y=0.135 $X2=0.153 $Y2=0.126
r136 32 38 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.122 $Y2=0.135
r137 30 70 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.198
+ $X2=0.486 $Y2=0.198
r138 27 30 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.216 $X2=0.484 $Y2=0.216
r139 26 66 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.198
+ $X2=0.378 $Y2=0.198
r140 23 26 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.216 $X2=0.378 $Y2=0.216
r141 22 26 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.216 $X2=0.378 $Y2=0.216
r142 21 47 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r143 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r144 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r145 13 15 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1345 $X2=0.135 $Y2=0.2025
r146 10 13 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1345
r147 5 13 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1345 $X2=0.135 $Y2=0.1345
r148 5 34 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r149 5 7 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1345 $X2=0.081 $Y2=0.2025
r150 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.1345
.ends

.subckt PM_AO33X2_ASAP7_75T_L%A3 2 5 7 10 14 16 VSS
c12 16 VSS 1.45426e-20 $X=0.189 $Y=0.14525
c13 14 VSS 0.00253613f $X=0.186 $Y=0.1465
c14 10 VSS 3.03777e-19 $X=0.189 $Y=0.135
c15 5 VSS 0.00115606f $X=0.189 $Y=0.135
c16 2 VSS 0.0592433f $X=0.189 $Y=0.0675
r17 15 16 0.0848765 $w=1.8e-08 $l=1.25e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.14525
r18 14 16 0.0848765 $w=1.8e-08 $l=1.25e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.1465 $X2=0.189 $Y2=0.14525
r19 10 15 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.144
r20 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r21 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AO33X2_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c13 10 VSS 0.00154873f $X=0.243 $Y=0.135
c14 5 VSS 0.00106612f $X=0.243 $Y=0.135
c15 2 VSS 0.059998f $X=0.243 $Y=0.0675
r16 10 14 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.19
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AO33X2_ASAP7_75T_L%A1 2 5 7 10 13 VSS
c15 13 VSS 0.00116352f $X=0.297 $Y=0.135
c16 10 VSS 3.80937e-19 $X=0.2995 $Y=0.116
c17 5 VSS 0.00110907f $X=0.297 $Y=0.135
c18 2 VSS 0.061059f $X=0.297 $Y=0.0675
r19 10 13 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.116 $X2=0.297 $Y2=0.135
r20 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r21 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AO33X2_ASAP7_75T_L%B1 2 5 7 10 VSS
c13 10 VSS 5.11375e-19 $X=0.3505 $Y=0.0795
c14 5 VSS 0.00107674f $X=0.351 $Y=0.135
c15 2 VSS 0.0623138f $X=0.351 $Y=0.0675
r16 10 13 3.76852 $w=1.8e-08 $l=5.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.0795 $X2=0.351 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.216
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AO33X2_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c12 10 VSS 4.78074e-19 $X=0.405 $Y=0.135
c13 5 VSS 0.00114557f $X=0.405 $Y=0.135
c14 2 VSS 0.0624468f $X=0.405 $Y=0.0675
r15 10 14 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.1465
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.216
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AO33X2_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c9 10 VSS 7.06488e-19 $X=0.459 $Y=0.135
c10 5 VSS 0.00170532f $X=0.459 $Y=0.135
c11 2 VSS 0.0661705f $X=0.459 $Y=0.0675
r12 10 14 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.1465
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.216
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AO33X2_ASAP7_75T_L%Y 1 2 5 6 7 10 14 15 16 19 25 28 35 VSS
c18 35 VSS 0.00756417f $X=0.108 $Y=0.054
c19 28 VSS 0.00187149f $X=0.0875 $Y=0.234
c20 27 VSS 0.00716014f $X=0.067 $Y=0.234
c21 25 VSS 0.00373005f $X=0.108 $Y=0.234
c22 23 VSS 0.00319564f $X=0.027 $Y=0.234
c23 22 VSS 6.90579e-19 $X=0.067 $Y=0.072
c24 21 VSS 0.0042436f $X=0.062 $Y=0.072
c25 20 VSS 0.00165989f $X=0.027 $Y=0.072
c26 19 VSS 3.75751e-19 $X=0.099 $Y=0.072
c27 18 VSS 7.00744e-19 $X=0.018 $Y=0.2125
c28 16 VSS 7.30811e-19 $X=0.018 $Y=0.144
c29 15 VSS 0.0023893f $X=0.018 $Y=0.126
c30 14 VSS 0.00322658f $X=0.019 $Y=0.1465
c31 12 VSS 5.68738e-19 $X=0.018 $Y=0.225
c32 10 VSS 0.00902026f $X=0.108 $Y=0.2025
c33 6 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c34 5 VSS 0.0105145f $X=0.108 $Y=0.0675
c35 1 VSS 5.945e-19 $X=0.125 $Y=0.0675
r36 33 35 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.063 $X2=0.108 $Y2=0.054
r37 27 28 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.067
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r38 25 28 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r39 23 27 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.067 $Y2=0.234
r40 21 22 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.062
+ $Y=0.072 $X2=0.067 $Y2=0.072
r41 20 21 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.072 $X2=0.062 $Y2=0.072
r42 19 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.099 $Y=0.072 $X2=0.108 $Y2=0.063
r43 19 22 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.072 $X2=0.067 $Y2=0.072
r44 17 18 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r45 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.144
r46 14 17 3.63272 $w=1.8e-08 $l=5.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1465 $X2=0.018 $Y2=0.2
r47 14 16 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1465 $X2=0.018 $Y2=0.144
r48 12 23 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r49 12 18 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r50 11 20 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.081 $X2=0.027 $Y2=0.072
r51 11 15 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.126
r52 10 25 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r53 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r54 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r55 5 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.054 $X2=0.108
+ $Y2=0.054
r56 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r57 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./AO33x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AO33x2_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 Y
* 
* Y	Y
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_12 N_A3_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_13 N_A2_M3_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_3_M4_d N_A1_M4_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_14 N_B1_M5_g N_3_M5_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_15 N_B2_M6_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 VSS N_B3_M7_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_Y_M8_d N_3_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M9 N_Y_M9_d N_3_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M10 noxref_11 N_A3_M10_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M11 VDD N_A2_M11_g noxref_11 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M12 noxref_11 N_A1_M12_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.189
M13 N_3_M13_d N_B1_M13_g noxref_11 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.341 $Y=0.189
M14 noxref_11 N_B2_M14_g N_3_M14_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.395 $Y=0.189
M15 N_3_M15_d N_B3_M15_g noxref_11 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.449 $Y=0.189
*
* 
* .include "AO33x2_ASAP7_75t_L.pex.sp.AO33X2_ASAP7_75T_L.pxi"
* BEGIN of "./AO33x2_ASAP7_75t_L.pex.sp.AO33X2_ASAP7_75T_L.pxi"
* File: AO33x2_ASAP7_75t_L.pex.sp.AO33X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:09:10 2017
* 
x_PM_AO33X2_ASAP7_75T_L%3 N_3_M0_g N_3_M8_g N_3_M1_g N_3_c_4_p N_3_M9_g N_3_M5_s
+ N_3_M4_d N_3_M14_s N_3_M13_d N_3_c_41_p N_3_M15_d N_3_c_45_p N_3_c_31_p
+ N_3_c_35_p N_3_c_29_p N_3_c_39_p N_3_c_5_p N_3_c_27_p N_3_c_11_p N_3_c_3_p
+ N_3_c_47_p N_3_c_8_p N_3_c_48_p N_3_c_10_p N_3_c_51_p N_3_c_14_p N_3_c_56_p
+ N_3_c_17_p N_3_c_57_p N_3_c_21_p N_3_c_13_p N_3_c_18_p N_3_c_46_p N_3_c_22_p
+ N_3_c_25_p VSS PM_AO33X2_ASAP7_75T_L%3
x_PM_AO33X2_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_61_n N_A3_M10_g N_A3_c_62_n A3
+ N_A3_c_68_p VSS PM_AO33X2_ASAP7_75T_L%A3
x_PM_AO33X2_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_74_n N_A2_M11_g N_A2_c_72_n A2 VSS
+ PM_AO33X2_ASAP7_75T_L%A2
x_PM_AO33X2_ASAP7_75T_L%A1 N_A1_M4_g N_A1_c_89_n N_A1_M12_g A1 N_A1_c_86_n VSS
+ PM_AO33X2_ASAP7_75T_L%A1
x_PM_AO33X2_ASAP7_75T_L%B1 N_B1_M5_g N_B1_c_103_n N_B1_M13_g B1 VSS
+ PM_AO33X2_ASAP7_75T_L%B1
x_PM_AO33X2_ASAP7_75T_L%B2 N_B2_M6_g N_B2_c_117_n N_B2_M14_g N_B2_c_113_n B2 VSS
+ PM_AO33X2_ASAP7_75T_L%B2
x_PM_AO33X2_ASAP7_75T_L%B3 N_B3_M7_g N_B3_c_130_n N_B3_M15_g N_B3_c_125_n B3 VSS
+ PM_AO33X2_ASAP7_75T_L%B3
x_PM_AO33X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_c_133_n N_Y_M9_d N_Y_M8_d
+ N_Y_c_148_p Y N_Y_c_135_n N_Y_c_136_n N_Y_c_138_n N_Y_c_141_n N_Y_c_142_n
+ N_Y_c_144_n VSS PM_AO33X2_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_A3_M2_g 0.00287079f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_A3_M2_g 2.64276e-19 $X=0.198 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_4 N_3_c_4_p N_A3_c_61_n 0.00148152f $X=0.135 $Y=0.1345 $X2=0.189 $Y2=0.135
cc_5 N_3_c_5_p N_A3_c_62_n 0.00611271f $X=0.153 $Y=0.081 $X2=0.189 $Y2=0.135
cc_6 N_3_c_3_p N_A3_c_62_n 0.00125352f $X=0.198 $Y=0.036 $X2=0.189 $Y2=0.135
cc_7 N_3_M1_g N_A2_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_8 N_3_c_8_p N_A2_M3_g 3.38929e-19 $X=0.252 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_9 N_3_c_8_p N_A2_c_72_n 0.00123604f $X=0.252 $Y=0.036 $X2=0.189 $Y2=0.135
cc_10 N_3_c_10_p N_A1_M4_g 2.56935e-19 $X=0.306 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_11 N_3_c_11_p A1 0.0013295f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.135
cc_12 N_3_c_10_p A1 0.00123604f $X=0.306 $Y=0.036 $X2=0.189 $Y2=0.135
cc_13 N_3_c_13_p N_A1_c_86_n 2.74755e-19 $X=0.396 $Y=0.198 $X2=0.189 $Y2=0.1465
cc_14 N_3_c_14_p N_B1_M5_g 2.64276e-19 $X=0.36 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_15 N_3_c_11_p B1 0.0013295f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.135
cc_16 N_3_c_14_p B1 0.00124805f $X=0.36 $Y=0.036 $X2=0.189 $Y2=0.135
cc_17 N_3_c_17_p N_B2_M6_g 3.38929e-19 $X=0.414 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_18 N_3_c_18_p N_B2_M6_g 2.76185e-19 $X=0.414 $Y=0.198 $X2=0.189 $Y2=0.0675
cc_19 N_3_c_17_p N_B2_c_113_n 0.00123064f $X=0.414 $Y=0.036 $X2=0.189 $Y2=0.135
cc_20 N_3_c_18_p N_B2_c_113_n 0.0012322f $X=0.414 $Y=0.198 $X2=0.189 $Y2=0.135
cc_21 N_3_c_21_p N_B3_M7_g 2.56935e-19 $X=0.468 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_22 N_3_c_22_p N_B3_M7_g 3.51973e-19 $X=0.468 $Y=0.198 $X2=0.189 $Y2=0.0675
cc_23 N_3_c_21_p N_B3_c_125_n 0.00123064f $X=0.468 $Y=0.036 $X2=0.189 $Y2=0.135
cc_24 N_3_c_22_p N_B3_c_125_n 0.00121543f $X=0.468 $Y=0.198 $X2=0.189 $Y2=0.135
cc_25 N_3_c_25_p N_B3_c_125_n 0.00392202f $X=0.513 $Y=0.164 $X2=0.189 $Y2=0.135
cc_26 N_3_c_4_p N_Y_M1_d 3.89919e-19 $X=0.135 $Y=0.1345 $X2=0.189 $Y2=0.0675
cc_27 N_3_c_27_p N_Y_c_133_n 0.0012315f $X=0.162 $Y=0.036 $X2=0.189 $Y2=0.135
cc_28 N_3_c_4_p N_Y_M9_d 3.83239e-19 $X=0.135 $Y=0.1345 $X2=0.189 $Y2=0.216
cc_29 N_3_c_29_p N_Y_c_135_n 2.91973e-19 $X=0.153 $Y=0.126 $X2=0.189 $Y2=0.144
cc_30 N_3_c_4_p N_Y_c_136_n 4.23217e-19 $X=0.135 $Y=0.1345 $X2=0.189 $Y2=0.14525
cc_31 N_3_c_31_p N_Y_c_136_n 8.31928e-19 $X=0.117 $Y=0.135 $X2=0.189 $Y2=0.14525
cc_32 N_3_M0_g N_Y_c_138_n 3.02973e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_33 N_3_c_31_p N_Y_c_138_n 0.0014224f $X=0.117 $Y=0.135 $X2=0 $Y2=0
cc_34 N_3_c_5_p N_Y_c_138_n 0.00110256f $X=0.153 $Y=0.081 $X2=0 $Y2=0
cc_35 N_3_c_35_p N_Y_c_141_n 4.13141e-19 $X=0.122 $Y=0.135 $X2=0 $Y2=0
cc_36 N_3_M0_g N_Y_c_142_n 3.32206e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_3_c_31_p N_Y_c_142_n 4.13141e-19 $X=0.117 $Y=0.135 $X2=0 $Y2=0
cc_38 N_3_M0_g N_Y_c_144_n 2.35764e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_3_c_39_p N_Y_c_144_n 0.00110256f $X=0.153 $Y=0.07 $X2=0 $Y2=0
cc_40 N_3_c_27_p N_Y_c_144_n 0.00110256f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_41 VSS N_3_c_41_p 0.00364136f $X=0.378 $Y=0.216 $X2=0.189 $Y2=0.135
cc_42 VSS N_3_c_11_p 0.00107252f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.135
cc_43 VSS N_3_c_13_p 3.5761e-19 $X=0.396 $Y=0.198 $X2=0.189 $Y2=0.135
cc_44 VSS N_3_c_41_p 0.0035539f $X=0.378 $Y=0.216 $X2=0.189 $Y2=0.144
cc_45 VSS N_3_c_45_p 0.00339392f $X=0.484 $Y=0.216 $X2=0.189 $Y2=0.144
cc_46 VSS N_3_c_46_p 0.00233206f $X=0.449 $Y=0.198 $X2=0.189 $Y2=0.144
cc_47 VSS N_3_c_47_p 2.20337e-19 $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_48 VSS N_3_c_48_p 2.20337e-19 $X=0.288 $Y=0.036 $X2=0 $Y2=0
cc_49 VSS N_3_c_45_p 2.9027e-19 $X=0.484 $Y=0.216 $X2=0 $Y2=0
cc_50 VSS N_3_c_18_p 0.00378945f $X=0.414 $Y=0.198 $X2=0 $Y2=0
cc_51 VSS N_3_c_51_p 2.20337e-19 $X=0.315 $Y=0.036 $X2=0 $Y2=0
cc_52 VSS N_3_c_41_p 0.00250965f $X=0.378 $Y=0.216 $X2=0 $Y2=0
cc_53 VSS N_3_c_13_p 0.00378945f $X=0.396 $Y=0.198 $X2=0 $Y2=0
cc_54 VSS N_3_c_47_p 3.56327e-19 $X=0.234 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_55 VSS N_3_c_48_p 3.56327e-19 $X=0.288 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_56 VSS N_3_c_56_p 3.48201e-19 $X=0.396 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_57 VSS N_3_c_57_p 3.48201e-19 $X=0.45 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_58 N_A3_M2_g N_A2_M3_g 0.00347357f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_59 N_A3_c_61_n N_A2_c_74_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.1345
cc_60 N_A3_c_62_n N_A2_c_72_n 0.00581377f $X=0.189 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_61 N_A3_M2_g N_A1_M4_g 2.69148e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_62 N_A3_c_68_p Y 2.86883e-19 $X=0.189 $Y=0.14525 $X2=0.135 $Y2=0.2025
cc_63 VSS A3 0.00114532f $X=0.186 $Y=0.1465 $X2=0.081 $Y2=0.1345
cc_64 N_A2_M3_g N_A1_M4_g 0.00330657f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_65 N_A2_c_74_n N_A1_c_89_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.1345
cc_66 N_A2_c_72_n A1 0.00581998f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_67 N_A2_M3_g N_B1_M5_g 2.74891e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_68 VSS N_A2_c_72_n 0.00114532f $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.1345
cc_69 VSS N_A2_M3_g 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0.378 $Y2=0.216
cc_70 VSS N_A2_c_72_n 0.00125352f $X=0.243 $Y=0.135 $X2=0.378 $Y2=0.216
cc_71 N_A1_M4_g N_B1_M5_g 0.00372052f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_72 N_A1_c_89_n N_B1_c_103_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081
+ $Y2=0.1345
cc_73 A1 B1 0.00389755f $X=0.2995 $Y=0.116 $X2=0.135 $Y2=0.0675
cc_74 N_A1_M4_g N_B2_M6_g 3.09654e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_75 VSS A1 9.89065e-19 $X=0.2995 $Y=0.116 $X2=0.135 $Y2=0.0675
cc_76 VSS N_A1_M4_g 2.64276e-19 $X=0.297 $Y=0.0675 $X2=0.378 $Y2=0.216
cc_77 VSS N_A1_c_86_n 0.00125352f $X=0.297 $Y=0.135 $X2=0.378 $Y2=0.216
cc_78 N_B1_M5_g N_B2_M6_g 0.00374235f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_79 N_B1_c_103_n N_B2_c_117_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.1345
cc_80 B1 N_B2_c_113_n 0.00483372f $X=0.3505 $Y=0.0795 $X2=0.135 $Y2=0.0675
cc_81 N_B1_M5_g N_B3_M7_g 3.09654e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_82 VSS N_B1_M5_g 3.57119e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_83 VSS B1 5.37372e-19 $X=0.3505 $Y=0.0795 $X2=0 $Y2=0
cc_84 N_B2_M6_g N_B3_M7_g 0.00372052f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_85 N_B2_c_117_n N_B3_c_130_n 9.33263e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.1345
cc_86 N_B2_c_113_n N_B3_c_125_n 0.0048308f $X=0.405 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_87 VSS N_B2_M6_g 2.28374e-19 $X=0.405 $Y=0.0675 $X2=0.484 $Y2=0.216
cc_88 VSS N_Y_c_148_p 2.23372e-19 $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.1345
cc_89 VSS N_Y_c_141_n 2.92683e-19 $X=0.108 $Y=0.234 $X2=0.361 $Y2=0.216

* END of "./AO33x2_ASAP7_75t_L.pex.sp.AO33X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI211x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:09:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI211x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI211x1_ASAP7_75t_L.pex.sp.pex"
* File: AOI211x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:09:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI211X1_ASAP7_75T_L%A2 2 5 8 11 13 19 21 24 27 29 VSS
c17 29 VSS 0.00716305f $X=0.018 $Y=0.135
c18 27 VSS 7.1121e-21 $X=0.1 $Y=0.135
c19 26 VSS 0.00388635f $X=0.091 $Y=0.135
c20 24 VSS 9.81575e-20 $X=0.109 $Y=0.135
c21 19 VSS 0.00709438f $X=0.018 $Y=0.144
c22 11 VSS 0.00532396f $X=0.135 $Y=0.135
c23 8 VSS 0.0623423f $X=0.135 $Y=0.0675
c24 2 VSS 0.0674994f $X=0.081 $Y=0.135
r25 26 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.091
+ $Y=0.135 $X2=0.1 $Y2=0.135
r26 24 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.135 $X2=0.1 $Y2=0.135
r27 24 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.109 $Y=0.135 $X2=0.109
+ $Y2=0.135
r28 22 29 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r29 22 26 4.34568 $w=1.8e-08 $l=6.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.091 $Y2=0.135
r30 19 29 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r31 19 21 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r32 11 25 23.6364 $w=2.2e-08 $l=2.6e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.109 $Y2=0.135
r33 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r34 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r35 2 25 25.4545 $w=2.2e-08 $l=2.8e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.109 $Y2=0.135
r36 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
.ends

.subckt PM_AOI211X1_ASAP7_75T_L%A1 2 7 10 13 18 25 30 VSS
c20 30 VSS 3.38062e-21 $X=0.198 $Y=0.135
c21 28 VSS 3.01861e-19 $X=0.215 $Y=0.135
c22 25 VSS 0.00281941f $X=0.189 $Y=0.135
c23 18 VSS 0.00355513f $X=0.192 $Y=0.119
c24 10 VSS 0.0725763f $X=0.243 $Y=0.135
c25 2 VSS 0.0627171f $X=0.189 $Y=0.0675
r26 30 31 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.135 $X2=0.2065 $Y2=0.135
r27 28 31 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.215
+ $Y=0.135 $X2=0.2065 $Y2=0.135
r28 28 29 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.215 $Y=0.135 $X2=0.215
+ $Y2=0.135
r29 25 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.198 $Y2=0.135
r30 16 25 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.135
r31 16 18 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.119
r32 10 29 25.4545 $w=2.2e-08 $l=2.8e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.215 $Y2=0.135
r33 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r34 5 29 23.6364 $w=2.2e-08 $l=2.6e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.215 $Y2=0.135
r35 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r36 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI211X1_ASAP7_75T_L%B 2 5 8 11 13 18 20 VSS
c20 23 VSS 6.94455e-20 $X=0.405 $Y=0.1305
c21 20 VSS 7.29745e-19 $X=0.405 $Y=0.135
c22 18 VSS 0.00326036f $X=0.405 $Y=0.113
c23 11 VSS 0.00749434f $X=0.459 $Y=0.135
c24 8 VSS 0.063706f $X=0.459 $Y=0.0675
c25 2 VSS 0.0673022f $X=0.405 $Y=0.135
r26 22 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.126 $X2=0.405 $Y2=0.1305
r27 20 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.1305
r28 18 22 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.113 $X2=0.405 $Y2=0.126
r29 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r30 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r31 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r32 2 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r33 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
.ends

.subckt PM_AOI211X1_ASAP7_75T_L%C 2 7 10 13 18 21 VSS
c24 21 VSS 6.65148e-19 $X=0.513 $Y=0.144
c25 18 VSS 0.00313242f $X=0.516 $Y=0.122
c26 10 VSS 0.0739416f $X=0.567 $Y=0.135
c27 2 VSS 0.0629624f $X=0.513 $Y=0.0675
r28 23 24 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.54 $Y=0.135 $X2=0.54
+ $Y2=0.135
r29 21 23 1.32 $w=2.5e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.144 $X2=0.54 $Y2=0.144
r30 16 21 0.266695 $w=2.5e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.126 $X2=0.513 $Y2=0.144
r31 16 18 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.126 $X2=0.513 $Y2=0.122
r32 10 24 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.567
+ $Y=0.135 $X2=0.54 $Y2=0.135
r33 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r34 5 24 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.54 $Y2=0.135
r35 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r36 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AOI211X1_ASAP7_75T_L%Y 1 6 7 11 12 15 19 23 24 25 26 27 28 29 30 31
+ 32 33 34 35 38 44 48 50 52 53 54 VSS
c45 56 VSS 4.55454e-19 $X=0.621 $Y=0.18
c46 55 VSS 2.54842e-19 $X=0.621 $Y=0.171
c47 54 VSS 0.00101339f $X=0.621 $Y=0.164
c48 53 VSS 7.59359e-19 $X=0.621 $Y=0.144
c49 52 VSS 0.00237814f $X=0.621 $Y=0.126
c50 50 VSS 1.23835e-19 $X=0.621 $Y=0.0655
c51 49 VSS 0.00104959f $X=0.621 $Y=0.063
c52 48 VSS 7.43007e-19 $X=0.624 $Y=0.068
c53 46 VSS 4.30151e-19 $X=0.621 $Y=0.189
c54 44 VSS 3.76365e-19 $X=0.608 $Y=0.198
c55 43 VSS 6.71593e-20 $X=0.554 $Y=0.198
c56 38 VSS 2.16721e-19 $X=0.54 $Y=0.198
c57 36 VSS 0.00216197f $X=0.612 $Y=0.198
c58 35 VSS 0.00274314f $X=0.583 $Y=0.036
c59 34 VSS 0.00118989f $X=0.554 $Y=0.036
c60 33 VSS 0.00587023f $X=0.55 $Y=0.036
c61 32 VSS 0.00524487f $X=0.504 $Y=0.036
c62 31 VSS 0.0011926f $X=0.449 $Y=0.036
c63 30 VSS 0.00625661f $X=0.442 $Y=0.036
c64 29 VSS 0.0129118f $X=0.396 $Y=0.036
c65 28 VSS 0.00577461f $X=0.288 $Y=0.036
c66 27 VSS 0.00253628f $X=0.229 $Y=0.036
c67 26 VSS 0.0049651f $X=0.22 $Y=0.036
c68 25 VSS 0.00543357f $X=0.18 $Y=0.036
c69 24 VSS 0.0030221f $X=0.123 $Y=0.036
c70 23 VSS 0.0100448f $X=0.486 $Y=0.036
c71 19 VSS 0.00428719f $X=0.108 $Y=0.036
c72 16 VSS 0.00642245f $X=0.612 $Y=0.036
c73 15 VSS 0.00453444f $X=0.54 $Y=0.2025
c74 11 VSS 5.97305e-19 $X=0.557 $Y=0.2025
c75 6 VSS 6.15054e-19 $X=0.503 $Y=0.0675
c76 1 VSS 4.46186e-19 $X=0.125 $Y=0.0675
r77 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.171 $X2=0.621 $Y2=0.18
r78 54 55 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.164 $X2=0.621 $Y2=0.171
r79 53 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.144 $X2=0.621 $Y2=0.164
r80 52 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.126 $X2=0.621 $Y2=0.144
r81 51 52 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.081 $X2=0.621 $Y2=0.126
r82 49 50 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.063 $X2=0.621 $Y2=0.0655
r83 48 51 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.068 $X2=0.621 $Y2=0.081
r84 48 50 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.068 $X2=0.621 $Y2=0.0655
r85 46 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.189 $X2=0.621 $Y2=0.18
r86 45 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.063
r87 43 44 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.554
+ $Y=0.198 $X2=0.608 $Y2=0.198
r88 38 43 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.198 $X2=0.554 $Y2=0.198
r89 36 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.198 $X2=0.621 $Y2=0.189
r90 36 44 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.198 $X2=0.608 $Y2=0.198
r91 34 35 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.554
+ $Y=0.036 $X2=0.583 $Y2=0.036
r92 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.55
+ $Y=0.036 $X2=0.554 $Y2=0.036
r93 32 33 3.12346 $w=1.8e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.55 $Y2=0.036
r94 30 31 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.442
+ $Y=0.036 $X2=0.449 $Y2=0.036
r95 29 30 3.12346 $w=1.8e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.442 $Y2=0.036
r96 28 29 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.396 $Y2=0.036
r97 27 28 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.229
+ $Y=0.036 $X2=0.288 $Y2=0.036
r98 26 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.22
+ $Y=0.036 $X2=0.229 $Y2=0.036
r99 25 26 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.22 $Y2=0.036
r100 24 25 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.123
+ $Y=0.036 $X2=0.18 $Y2=0.036
r101 22 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.504 $Y2=0.036
r102 22 31 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.449 $Y2=0.036
r103 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036
+ $X2=0.486 $Y2=0.036
r104 18 24 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.123 $Y2=0.036
r105 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r106 16 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r107 16 35 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.583 $Y2=0.036
r108 15 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.198 $X2=0.54
+ $Y2=0.198
r109 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r110 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r111 10 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.486 $Y=0.0675 $X2=0.486 $Y2=0.036
r112 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.486 $Y2=0.0675
r113 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.0675 $X2=0.486 $Y2=0.0675
r114 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r115 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.11 $Y2=0.0675
.ends


* END of "./AOI211x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI211x1_ASAP7_75t_L  VSS VDD A2 A1 B C Y
* 
* Y	Y
* C	C
* B	B
* A1	A1
* A2	A2
M0 noxref_10 N_A2_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M1 VSS N_A1_M1_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M2 N_Y_M2_d N_B_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M3 VSS N_C_M3_g N_Y_M3_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M4 noxref_7 N_A2_M4_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 noxref_7 N_A2_M5_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 noxref_7 N_A1_M6_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M7 noxref_7 N_A1_M7_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M8 noxref_7 N_B_M8_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M9 noxref_7 N_B_M9_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M10 N_Y_M10_d N_C_M10_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M11 N_Y_M11_d N_C_M11_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
*
* 
* .include "AOI211x1_ASAP7_75t_L.pex.sp.AOI211X1_ASAP7_75T_L.pxi"
* BEGIN of "./AOI211x1_ASAP7_75t_L.pex.sp.AOI211X1_ASAP7_75T_L.pxi"
* File: AOI211x1_ASAP7_75t_L.pex.sp.AOI211X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:09:33 2017
* 
x_PM_AOI211X1_ASAP7_75T_L%A2 N_A2_c_1_p N_A2_M4_g N_A2_M0_g N_A2_c_4_p N_A2_M5_g
+ N_A2_c_6_p A2 N_A2_c_7_p N_A2_c_10_p N_A2_c_5_p VSS PM_AOI211X1_ASAP7_75T_L%A2
x_PM_AOI211X1_ASAP7_75T_L%A1 N_A1_M1_g N_A1_M6_g N_A1_c_20_n N_A1_M7_g A1
+ N_A1_c_23_n N_A1_c_24_n VSS PM_AOI211X1_ASAP7_75T_L%A1
x_PM_AOI211X1_ASAP7_75T_L%B N_B_c_39_p N_B_M8_g N_B_M2_g N_B_c_42_p N_B_M9_g B
+ N_B_c_44_p VSS PM_AOI211X1_ASAP7_75T_L%B
x_PM_AOI211X1_ASAP7_75T_L%C N_C_M3_g N_C_M10_g N_C_c_60_n N_C_M11_g C N_C_c_63_n
+ VSS PM_AOI211X1_ASAP7_75T_L%C
x_PM_AOI211X1_ASAP7_75T_L%Y N_Y_M0_s N_Y_M3_s N_Y_M2_d N_Y_M11_d N_Y_M10_d
+ N_Y_c_118_n N_Y_c_82_n N_Y_c_98_n N_Y_c_83_n N_Y_c_87_n N_Y_c_89_n N_Y_c_91_n
+ N_Y_c_92_n N_Y_c_115_n N_Y_c_93_n N_Y_c_95_n N_Y_c_96_n N_Y_c_99_n N_Y_c_101_n
+ N_Y_c_102_n N_Y_c_103_n N_Y_c_106_n Y N_Y_c_107_n N_Y_c_108_n N_Y_c_110_n
+ N_Y_c_111_n VSS PM_AOI211X1_ASAP7_75T_L%Y
cc_1 N_A2_c_1_p N_A1_M1_g 2.69148e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_2 N_A2_M0_g N_A1_M1_g 0.00323392f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A2_M0_g N_A1_c_20_n 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_4 N_A2_c_4_p N_A1_c_20_n 0.00126537f $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_5 N_A2_c_5_p A1 4.69586e-19 $X=0.018 $Y=0.135 $X2=0.192 $Y2=0.119
cc_6 N_A2_c_6_p N_A1_c_23_n 3.05337e-19 $X=0.018 $Y=0.144 $X2=0.189 $Y2=0.135
cc_7 N_A2_c_7_p N_A1_c_24_n 3.59908e-19 $X=0.109 $Y=0.135 $X2=0.198 $Y2=0.135
cc_8 VSS N_A2_c_4_p 3.80307e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_9 VSS N_A2_c_4_p 3.61857e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_10 VSS N_A2_c_10_p 3.56949e-19 $X=0.1 $Y=0.135 $X2=0 $Y2=0
cc_11 VSS N_A2_M0_g 4.58656e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_12 N_A2_c_5_p N_Y_c_82_n 0.00123601f $X=0.018 $Y=0.135 $X2=0 $Y2=0
cc_13 N_A2_c_1_p N_Y_c_83_n 5.44741e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_14 N_A2_c_4_p N_Y_c_83_n 3.40112e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_15 N_A2_c_10_p N_Y_c_83_n 3.69009e-19 $X=0.1 $Y=0.135 $X2=0 $Y2=0
cc_16 N_A2_c_5_p N_Y_c_83_n 3.16757e-19 $X=0.018 $Y=0.135 $X2=0 $Y2=0
cc_17 N_A2_M0_g N_Y_c_87_n 4.58656e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_18 A1 B 2.10129e-19 $X=0.192 $Y=0.119 $X2=0 $Y2=0
cc_19 VSS N_A1_c_20_n 3.80618e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_20 VSS N_A1_c_23_n 0.0020361f $X=0.189 $Y=0.135 $X2=0.135 $Y2=0.135
cc_21 VSS N_A1_c_20_n 4.58656e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_22 VSS N_A1_M1_g 2.34993e-19 $X=0.189 $Y=0.0675 $X2=0.091 $Y2=0.135
cc_23 VSS N_A1_c_23_n 0.00421074f $X=0.189 $Y=0.135 $X2=0.091 $Y2=0.135
cc_24 VSS N_A1_c_20_n 2.80703e-19 $X=0.243 $Y=0.135 $X2=0.1 $Y2=0.135
cc_25 VSS N_A1_c_23_n 2.57943e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_26 A1 N_Y_c_82_n 8.24105e-19 $X=0.192 $Y=0.119 $X2=0.018 $Y2=0.144
cc_27 N_A1_M1_g N_Y_c_89_n 2.34993e-19 $X=0.189 $Y=0.0675 $X2=0.091 $Y2=0.135
cc_28 A1 N_Y_c_89_n 0.00398267f $X=0.192 $Y=0.119 $X2=0.091 $Y2=0.135
cc_29 N_A1_c_20_n N_Y_c_91_n 2.62066e-19 $X=0.243 $Y=0.135 $X2=0.1 $Y2=0.135
cc_30 N_A1_c_20_n N_Y_c_92_n 4.58656e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 N_B_c_39_p N_C_M3_g 2.74891e-19 $X=0.405 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_32 N_B_M2_g N_C_M3_g 0.00359705f $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_33 N_B_M2_g N_C_c_60_n 2.74891e-19 $X=0.459 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_34 N_B_c_42_p N_C_c_60_n 0.0013547f $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.135
cc_35 B C 7.4949e-19 $X=0.405 $Y=0.113 $X2=0.192 $Y2=0.119
cc_36 N_B_c_44_p N_C_c_63_n 8.47457e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_37 VSS N_B_c_42_p 3.78279e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_38 VSS N_B_c_42_p 8.00061e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_39 VSS N_B_c_44_p 0.00133904f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_40 VSS N_B_c_39_p 2.52885e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_41 VSS N_B_c_44_p 0.00452229f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_42 VSS N_B_c_44_p 3.13188e-19 $X=0.405 $Y=0.135 $X2=0.189 $Y2=0.135
cc_43 VSS N_B_c_39_p 2.38303e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_44 VSS N_B_M2_g 4.24257e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_45 VSS N_B_c_42_p 2.04785e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_46 N_B_c_39_p N_Y_c_93_n 2.34993e-19 $X=0.405 $Y=0.135 $X2=0.198 $Y2=0.135
cc_47 B N_Y_c_93_n 0.0044179f $X=0.405 $Y=0.113 $X2=0.198 $Y2=0.135
cc_48 N_B_c_42_p N_Y_c_95_n 3.10711e-19 $X=0.459 $Y=0.135 $X2=0.2065 $Y2=0.135
cc_49 N_B_M2_g N_Y_c_96_n 4.52923e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_50 VSS N_C_c_60_n 2.64781e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_51 VSS N_C_M3_g 2.87679e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_52 VSS N_C_c_63_n 4.40991e-19 $X=0.513 $Y=0.144 $X2=0 $Y2=0
cc_53 N_C_c_60_n N_Y_M11_d 3.80538e-19 $X=0.567 $Y=0.135 $X2=0.459 $Y2=0.135
cc_54 C N_Y_c_98_n 0.00155697f $X=0.516 $Y=0.122 $X2=0.405 $Y2=0.1305
cc_55 N_C_M3_g N_Y_c_99_n 2.31683e-19 $X=0.513 $Y=0.0675 $X2=0.459 $Y2=0.135
cc_56 C N_Y_c_99_n 0.00445939f $X=0.516 $Y=0.122 $X2=0.459 $Y2=0.135
cc_57 N_C_c_60_n N_Y_c_101_n 2.42614e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_58 N_C_c_60_n N_Y_c_102_n 4.59758e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_59 N_C_M3_g N_Y_c_103_n 2.09481e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_60 N_C_c_60_n N_Y_c_103_n 5.86791e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_61 N_C_c_63_n N_Y_c_103_n 7.76964e-19 $X=0.513 $Y=0.144 $X2=0 $Y2=0
cc_62 N_C_c_60_n N_Y_c_106_n 3.95625e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_63 C N_Y_c_107_n 4.26481e-19 $X=0.516 $Y=0.122 $X2=0 $Y2=0
cc_64 N_C_c_60_n N_Y_c_108_n 3.86913e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_65 C N_Y_c_108_n 6.35237e-19 $X=0.516 $Y=0.122 $X2=0 $Y2=0
cc_66 N_C_c_63_n N_Y_c_110_n 3.91894e-19 $X=0.513 $Y=0.144 $X2=0 $Y2=0
cc_67 N_C_c_63_n N_Y_c_111_n 3.6017e-19 $X=0.513 $Y=0.144 $X2=0 $Y2=0
cc_68 VSS N_Y_c_82_n 9.50123e-19 $X=0.108 $Y=0.2025 $X2=0.018 $Y2=0.144
cc_69 VSS N_Y_c_83_n 4.01707e-19 $X=0.18 $Y=0.234 $X2=0.109 $Y2=0.135
cc_70 VSS N_Y_c_91_n 4.01707e-19 $X=0.288 $Y=0.234 $X2=0.1 $Y2=0.135
cc_71 VSS N_Y_c_115_n 7.4287e-19 $X=0.306 $Y=0.198 $X2=0.018 $Y2=0.135
cc_72 VSS N_Y_c_95_n 7.4287e-19 $X=0.396 $Y=0.198 $X2=0 $Y2=0
cc_73 VSS N_Y_c_103_n 3.08477e-19 $X=0.432 $Y=0.198 $X2=0 $Y2=0
cc_74 VSS N_Y_c_118_n 0.00326537f $X=0.486 $Y=0.2025 $X2=0 $Y2=0
cc_75 VSS N_Y_c_118_n 0.00371671f $X=0.592 $Y=0.2025 $X2=0 $Y2=0
cc_76 VSS N_Y_c_118_n 0.00249183f $X=0.594 $Y=0.234 $X2=0 $Y2=0
cc_77 VSS N_Y_c_98_n 0.00107252f $X=0.486 $Y=0.2025 $X2=0.405 $Y2=0.1305
cc_78 VSS N_Y_c_103_n 4.79394e-19 $X=0.486 $Y=0.2025 $X2=0 $Y2=0
cc_79 VSS N_Y_c_103_n 0.00769046f $X=0.594 $Y=0.234 $X2=0 $Y2=0
cc_80 VSS N_Y_c_106_n 0.00285209f $X=0.592 $Y=0.2025 $X2=0 $Y2=0
cc_81 VSS N_Y_c_111_n 3.46411e-19 $X=0.592 $Y=0.2025 $X2=0 $Y2=0
cc_82 VSS N_Y_c_87_n 4.6368e-19 $X=0.18 $Y=0.036 $X2=0.081 $Y2=0.135

* END of "./AOI211x1_ASAP7_75t_L.pex.sp.AOI211X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI211xp5_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:09:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI211xp5_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI211xp5_ASAP7_75t_L.pex.sp.pex"
* File: AOI211xp5_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:09:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI211XP5_ASAP7_75T_L%A2 2 5 7 13 14 20 23 25 VSS
c12 25 VSS 0.00462465f $X=0.027 $Y=0.135
c13 23 VSS 4.81186e-19 $X=0.0605 $Y=0.135
c14 22 VSS 5.77998e-19 $X=0.04 $Y=0.135
c15 20 VSS 2.24273e-19 $X=0.081 $Y=0.135
c16 15 VSS 4.88551e-19 $X=0.027 $Y=0.1755
c17 14 VSS 0.00101957f $X=0.027 $Y=0.164
c18 13 VSS 0.00212468f $X=0.023 $Y=0.187
c19 5 VSS 0.00258107f $X=0.081 $Y=0.135
c20 2 VSS 0.0662757f $X=0.081 $Y=0.054
r21 22 23 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.135 $X2=0.0605 $Y2=0.135
r22 20 23 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0605 $Y2=0.135
r23 18 25 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.135 $X2=0.027 $Y2=0.135
r24 18 22 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.135 $X2=0.04 $Y2=0.135
r25 14 15 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.164 $X2=0.027 $Y2=0.1755
r26 13 15 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.187 $X2=0.027 $Y2=0.1755
r27 11 25 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.144 $X2=0.027 $Y2=0.135
r28 11 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.144 $X2=0.027 $Y2=0.164
r29 5 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r30 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r31 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI211XP5_ASAP7_75T_L%A1 2 5 7 10 13 16 VSS
c14 16 VSS 2.89025e-20 $X=0.135 $Y=0.1305
c15 13 VSS 3.31287e-19 $X=0.135 $Y=0.135
c16 10 VSS 0.00106027f $X=0.134 $Y=0.109
c17 5 VSS 0.00117984f $X=0.135 $Y=0.135
c18 2 VSS 0.0601206f $X=0.135 $Y=0.054
r19 15 16 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.1305
r20 13 16 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.1305
r21 10 15 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.109 $X2=0.135 $Y2=0.126
r22 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r23 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r24 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI211XP5_ASAP7_75T_L%B 2 5 7 10 14 VSS
c12 10 VSS 9.85944e-19 $X=0.189 $Y=0.135
c13 5 VSS 0.00116143f $X=0.189 $Y=0.135
c14 2 VSS 0.0590835f $X=0.189 $Y=0.054
r15 10 14 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.148
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI211XP5_ASAP7_75T_L%C 2 5 7 10 VSS
c10 10 VSS 9.75038e-19 $X=0.241 $Y=0.123
c11 5 VSS 0.00170784f $X=0.243 $Y=0.135
c12 2 VSS 0.0618315f $X=0.243 $Y=0.054
r13 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.123 $X2=0.243 $Y2=0.135
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI211XP5_ASAP7_75T_L%Y 1 4 6 7 10 11 12 15 24 27 29 31 37 38 39 41
+ 42 43 48 50 VSS
c26 50 VSS 0.00431076f $X=0.297 $Y=0.164
c27 49 VSS 0.00131846f $X=0.297 $Y=0.07
c28 48 VSS 0.00131846f $X=0.299 $Y=0.172
c29 44 VSS 0.00236172f $X=0.27 $Y=0.198
c30 43 VSS 5.17397e-19 $X=0.252 $Y=0.198
c31 42 VSS 0.00175846f $X=0.234 $Y=0.198
c32 41 VSS 5.17397e-19 $X=0.198 $Y=0.198
c33 40 VSS 2.28963e-19 $X=0.18 $Y=0.198
c34 39 VSS 4.67884e-19 $X=0.176 $Y=0.198
c35 38 VSS 8.46035e-21 $X=0.144 $Y=0.198
c36 37 VSS 7.17059e-19 $X=0.126 $Y=0.198
c37 32 VSS 0.00390806f $X=0.288 $Y=0.198
c38 31 VSS 0.00146362f $X=0.252 $Y=0.036
c39 30 VSS 0.00346254f $X=0.234 $Y=0.036
c40 29 VSS 0.00146362f $X=0.198 $Y=0.036
c41 28 VSS 0.00577782f $X=0.18 $Y=0.036
c42 27 VSS 0.00146362f $X=0.144 $Y=0.036
c43 26 VSS 0.00257933f $X=0.126 $Y=0.036
c44 25 VSS 9.06382e-19 $X=0.099 $Y=0.036
c45 24 VSS 0.00532554f $X=0.09 $Y=0.036
c46 16 VSS 0.00884695f $X=0.288 $Y=0.036
c47 15 VSS 0.00210856f $X=0.108 $Y=0.2025
c48 11 VSS 6.64001e-19 $X=0.125 $Y=0.2025
c49 10 VSS 0.00790803f $X=0.216 $Y=0.054
c50 6 VSS 5.3314e-19 $X=0.233 $Y=0.054
c51 4 VSS 0.00348545f $X=0.056 $Y=0.054
c52 1 VSS 2.6657e-19 $X=0.071 $Y=0.054
r53 49 50 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.07 $X2=0.297 $Y2=0.164
r54 48 50 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.172 $X2=0.297 $Y2=0.164
r55 46 48 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.172
r56 45 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.07
r57 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.27 $Y2=0.198
r58 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.252 $Y2=0.198
r59 41 42 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.198 $X2=0.234 $Y2=0.198
r60 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.198 $X2=0.198 $Y2=0.198
r61 39 40 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.198 $X2=0.18 $Y2=0.198
r62 38 39 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.198 $X2=0.176 $Y2=0.198
r63 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.198 $X2=0.144 $Y2=0.198
r64 34 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.198 $X2=0.126 $Y2=0.198
r65 32 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.198 $X2=0.297 $Y2=0.189
r66 32 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.27 $Y2=0.198
r67 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r68 28 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r69 27 28 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.18 $Y2=0.036
r70 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r71 25 26 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.036 $X2=0.126 $Y2=0.036
r72 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.099 $Y2=0.036
r73 22 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.234 $Y2=0.036
r74 22 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.198 $Y2=0.036
r75 18 24 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.09 $Y2=0.036
r76 16 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r77 16 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.252 $Y2=0.036
r78 15 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.198 $X2=0.108
+ $Y2=0.198
r79 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r80 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r81 10 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r82 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.054 $X2=0.216 $Y2=0.054
r83 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.054 $X2=0.216 $Y2=0.054
r84 4 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r85 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.054 $X2=0.056 $Y2=0.054
.ends


* END of "./AOI211xp5_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI211xp5_ASAP7_75t_L  VSS VDD A2 A1 B C Y
* 
* Y	Y
* C	C
* B	B
* A1	A1
* A2	A2
M0 noxref_9 N_A2_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 VSS N_A1_M1_g noxref_9 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_B_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 VSS N_C_M3_g N_Y_M3_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_A2_M4_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 noxref_7 N_A1_M5_g N_Y_M5_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 noxref_10 N_B_M6_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M7 VDD N_C_M7_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
*
* 
* .include "AOI211xp5_ASAP7_75t_L.pex.sp.AOI211XP5_ASAP7_75T_L.pxi"
* BEGIN of "./AOI211xp5_ASAP7_75t_L.pex.sp.AOI211XP5_ASAP7_75T_L.pxi"
* File: AOI211xp5_ASAP7_75t_L.pex.sp.AOI211XP5_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:09:56 2017
* 
x_PM_AOI211XP5_ASAP7_75T_L%A2 N_A2_M0_g N_A2_c_2_p N_A2_M4_g A2 N_A2_c_4_p
+ N_A2_c_5_p N_A2_c_9_p N_A2_c_3_p VSS PM_AOI211XP5_ASAP7_75T_L%A2
x_PM_AOI211XP5_ASAP7_75T_L%A1 N_A1_M1_g N_A1_c_14_n N_A1_M5_g A1 N_A1_c_16_n
+ N_A1_c_17_n VSS PM_AOI211XP5_ASAP7_75T_L%A1
x_PM_AOI211XP5_ASAP7_75T_L%B N_B_M2_g N_B_c_29_n N_B_M6_g N_B_c_30_n B VSS
+ PM_AOI211XP5_ASAP7_75T_L%B
x_PM_AOI211XP5_ASAP7_75T_L%C N_C_M3_g N_C_c_41_n N_C_M7_g C VSS
+ PM_AOI211XP5_ASAP7_75T_L%C
x_PM_AOI211XP5_ASAP7_75T_L%Y N_Y_M0_s N_Y_c_49_n N_Y_M3_s N_Y_M2_d N_Y_c_56_n
+ N_Y_M5_s N_Y_M4_d N_Y_c_68_n N_Y_c_50_n N_Y_c_52_n N_Y_c_57_n N_Y_c_62_n
+ N_Y_c_72_n N_Y_c_54_n N_Y_c_73_n N_Y_c_59_n N_Y_c_74_p N_Y_c_64_n Y N_Y_c_66_n
+ VSS PM_AOI211XP5_ASAP7_75T_L%Y
cc_1 N_A2_M0_g N_A1_M1_g 0.00364065f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A2_c_2_p N_A1_c_14_n 9.83624e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A2_c_3_p A1 0.00108189f $X=0.027 $Y=0.135 $X2=0.134 $Y2=0.109
cc_4 N_A2_c_4_p N_A1_c_16_n 4.17105e-19 $X=0.027 $Y=0.164 $X2=0.135 $Y2=0.135
cc_5 N_A2_c_5_p N_A1_c_17_n 6.03818e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.1305
cc_6 N_A2_M0_g N_B_M2_g 2.6588e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_7 VSS N_A2_c_4_p 0.00163879f $X=0.027 $Y=0.164 $X2=0.135 $Y2=0.135
cc_8 VSS N_A2_M0_g 4.01862e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_9 VSS N_A2_c_9_p 9.66105e-19 $X=0.0605 $Y=0.135 $X2=0 $Y2=0
cc_10 N_A2_c_3_p N_Y_c_49_n 3.85925e-19 $X=0.027 $Y=0.135 $X2=0.135 $Y2=0.135
cc_11 N_A2_M0_g N_Y_c_50_n 4.01862e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_12 N_A2_c_9_p N_Y_c_50_n 9.13307e-19 $X=0.0605 $Y=0.135 $X2=0 $Y2=0
cc_13 N_A1_M1_g N_B_M2_g 0.0032267f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_14 N_A1_c_14_n N_B_c_29_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 A1 N_B_c_30_n 0.0045518f $X=0.134 $Y=0.109 $X2=0 $Y2=0
cc_16 N_A1_M1_g N_C_M3_g 2.60137e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_17 VSS N_A1_M1_g 2.38303e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_18 N_A1_M1_g N_Y_c_52_n 2.64276e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_19 A1 N_Y_c_52_n 0.00124805f $X=0.134 $Y=0.109 $X2=0 $Y2=0
cc_20 N_A1_M1_g N_Y_c_54_n 2.76185e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_21 N_A1_c_16_n N_Y_c_54_n 0.0012322f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_22 N_B_M2_g N_C_M3_g 0.0033937f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_23 N_B_c_29_n N_C_c_41_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_B_c_30_n C 0.0046131f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_25 N_B_c_30_n N_Y_c_56_n 3.31541e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_26 N_B_M2_g N_Y_c_57_n 2.64276e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_27 N_B_c_30_n N_Y_c_57_n 0.00124805f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_28 N_B_M2_g N_Y_c_59_n 3.51973e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_29 N_B_c_30_n N_Y_c_59_n 0.00121543f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_30 C N_Y_c_56_n 3.31541e-19 $X=0.241 $Y=0.123 $X2=0.134 $Y2=0.109
cc_31 N_C_M3_g N_Y_c_62_n 2.64276e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_32 C N_Y_c_62_n 0.00124805f $X=0.241 $Y=0.123 $X2=0 $Y2=0
cc_33 N_C_M3_g N_Y_c_64_n 3.51973e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_34 C N_Y_c_64_n 0.00121543f $X=0.241 $Y=0.123 $X2=0 $Y2=0
cc_35 C N_Y_c_66_n 0.00441847f $X=0.241 $Y=0.123 $X2=0 $Y2=0
cc_36 VSS N_Y_c_49_n 8.7738e-19 $X=0.056 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_37 VSS N_Y_c_68_n 0.0036868f $X=0.056 $Y=0.2025 $X2=0.027 $Y2=0.1755
cc_38 VSS N_Y_c_68_n 0.00359726f $X=0.162 $Y=0.2025 $X2=0.027 $Y2=0.1755
cc_39 VSS N_Y_c_68_n 0.00189275f $X=0.162 $Y=0.234 $X2=0.027 $Y2=0.1755
cc_40 VSS N_Y_c_68_n 6.35113e-19 $X=0.099 $Y=0.234 $X2=0.027 $Y2=0.1755
cc_41 VSS N_Y_c_72_n 0.00666759f $X=0.162 $Y=0.234 $X2=0 $Y2=0
cc_42 VSS N_Y_c_73_n 0.00262229f $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_43 VSS N_Y_c_74_p 4.30621e-19 $X=0.234 $Y=0.198 $X2=0.081 $Y2=0.054

* END of "./AOI211xp5_ASAP7_75t_L.pex.sp.AOI211XP5_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI21x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:10:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI21x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI21x1_ASAP7_75t_L.pex.sp.pex"
* File: AOI21x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:10:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI21X1_ASAP7_75T_L%B 2 5 7 10 13 15 22 28 29 30 31 32 33 34 35 36 39
+ 43 VSS
c36 43 VSS 1.30627e-19 $X=0.351 $Y=0.171
c37 39 VSS 2.04795e-19 $X=0.351 $Y=0.134
c38 36 VSS 1.62028e-19 $X=0.3375 $Y=0.198
c39 35 VSS 2.77255e-19 $X=0.333 $Y=0.198
c40 34 VSS 7.99121e-21 $X=0.306 $Y=0.198
c41 33 VSS 0.00327176f $X=0.288 $Y=0.198
c42 32 VSS 2.08366e-19 $X=0.256 $Y=0.198
c43 31 VSS 1.73836e-19 $X=0.227 $Y=0.198
c44 30 VSS 0.0016554f $X=0.19 $Y=0.198
c45 29 VSS 0.00126552f $X=0.163 $Y=0.198
c46 28 VSS 4.27363e-19 $X=0.126 $Y=0.198
c47 27 VSS 5.57344e-19 $X=0.099 $Y=0.198
c48 26 VSS 8.76255e-19 $X=0.09 $Y=0.198
c49 25 VSS 0.00103635f $X=0.342 $Y=0.198
c50 22 VSS 7.77592e-19 $X=0.0835 $Y=0.1355
c51 13 VSS 0.00239017f $X=0.351 $Y=0.135
c52 10 VSS 0.0654656f $X=0.351 $Y=0.054
c53 5 VSS 0.00243208f $X=0.081 $Y=0.135
c54 2 VSS 0.0651238f $X=0.081 $Y=0.054
r55 42 43 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.151 $X2=0.351 $Y2=0.171
r56 39 42 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.134 $X2=0.351 $Y2=0.151
r57 37 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.171
r58 35 36 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.198 $X2=0.3375 $Y2=0.198
r59 34 35 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.198 $X2=0.333 $Y2=0.198
r60 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.306 $Y2=0.198
r61 32 33 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.198 $X2=0.288 $Y2=0.198
r62 31 32 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.227
+ $Y=0.198 $X2=0.256 $Y2=0.198
r63 30 31 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.19
+ $Y=0.198 $X2=0.227 $Y2=0.198
r64 29 30 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.163
+ $Y=0.198 $X2=0.19 $Y2=0.198
r65 28 29 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.198 $X2=0.163 $Y2=0.198
r66 27 28 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.198 $X2=0.126 $Y2=0.198
r67 26 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.198 $X2=0.099 $Y2=0.198
r68 25 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.198 $X2=0.351 $Y2=0.189
r69 25 36 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.3375 $Y2=0.198
r70 23 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.171 $X2=0.081 $Y2=0.18
r71 22 23 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.134 $X2=0.081 $Y2=0.171
r72 17 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.189 $X2=0.09 $Y2=0.198
r73 17 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.189 $X2=0.081 $Y2=0.18
r74 13 39 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.134 $X2=0.351
+ $Y2=0.134
r75 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r76 10 13 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.054 $X2=0.351 $Y2=0.135
r77 5 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.134 $X2=0.081
+ $Y2=0.134
r78 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r79 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI21X1_ASAP7_75T_L%A1 2 5 7 10 13 15 23 24 25 26 27 28 29 30 33 36
+ 37 38 VSS
c37 38 VSS 2.64813e-20 $X=0.297 $Y=0.1295
c38 37 VSS 1.16016e-19 $X=0.297 $Y=0.125
c39 36 VSS 1.88379e-19 $X=0.297 $Y=0.116
c40 35 VSS 3.51388e-19 $X=0.297 $Y=0.099
c41 33 VSS 4.98993e-20 $X=0.297 $Y=0.134
c42 30 VSS 9.36428e-19 $X=0.256 $Y=0.072
c43 29 VSS 0.00235496f $X=0.227 $Y=0.072
c44 28 VSS 6.28049e-19 $X=0.19 $Y=0.072
c45 27 VSS 1.08538e-19 $X=0.163 $Y=0.072
c46 26 VSS 1.13858e-19 $X=0.144 $Y=0.072
c47 25 VSS 3.61504e-19 $X=0.288 $Y=0.072
c48 24 VSS 0.00161747f $X=0.1345 $Y=0.1355
c49 23 VSS 5.19271e-20 $X=0.135 $Y=0.1165
c50 22 VSS 3.51388e-19 $X=0.135 $Y=0.099
c51 13 VSS 0.00167162f $X=0.297 $Y=0.135
c52 10 VSS 0.0606486f $X=0.297 $Y=0.0675
c53 5 VSS 0.00154002f $X=0.135 $Y=0.135
c54 2 VSS 0.0604776f $X=0.135 $Y=0.0675
r55 37 38 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.125 $X2=0.297 $Y2=0.1295
r56 36 37 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.116 $X2=0.297 $Y2=0.125
r57 35 36 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.099 $X2=0.297 $Y2=0.116
r58 33 38 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.134 $X2=0.297 $Y2=0.1295
r59 31 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.081 $X2=0.297 $Y2=0.099
r60 29 30 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.227
+ $Y=0.072 $X2=0.256 $Y2=0.072
r61 28 29 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.19
+ $Y=0.072 $X2=0.227 $Y2=0.072
r62 27 28 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.163
+ $Y=0.072 $X2=0.19 $Y2=0.072
r63 26 27 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.163 $Y2=0.072
r64 25 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.072 $X2=0.297 $Y2=0.081
r65 25 30 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.256 $Y2=0.072
r66 23 24 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.1165 $X2=0.135 $Y2=0.134
r67 22 23 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.099 $X2=0.135 $Y2=0.1165
r68 17 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.081 $X2=0.144 $Y2=0.072
r69 17 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.081 $X2=0.135 $Y2=0.099
r70 13 33 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.134 $X2=0.297
+ $Y2=0.134
r71 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r72 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r73 5 24 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.134 $X2=0.135
+ $Y2=0.134
r74 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r75 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI21X1_ASAP7_75T_L%A2 2 7 10 13 15 18 VSS
c29 18 VSS 0.00293381f $X=0.2085 $Y=0.1355
c30 13 VSS 0.00737317f $X=0.243 $Y=0.135
c31 10 VSS 0.0624282f $X=0.243 $Y=0.0675
c32 2 VSS 0.0626776f $X=0.189 $Y=0.0675
r33 18 20 0.797927 $w=4.825e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2085 $Y=0.135 $X2=0.24 $Y2=0.135
r34 13 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.24 $Y=0.134 $X2=0.24
+ $Y2=0.134
r35 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r36 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r37 5 13 46.3636 $w=2.2e-08 $l=5.1e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.24 $Y2=0.135
r38 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r39 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI21X1_ASAP7_75T_L%Y 2 3 6 8 9 12 19 22 24 27 32 44 50 52 58 59 64
+ 74 VSS
c25 74 VSS 0.00340693f $X=0.396 $Y=0.234
c26 73 VSS 0.00277971f $X=0.405 $Y=0.234
c27 67 VSS 0.00102136f $X=0.045 $Y=0.234
c28 66 VSS 0.00328948f $X=0.036 $Y=0.234
c29 64 VSS 0.00235662f $X=0.054 $Y=0.234
c30 60 VSS 2.98008e-19 $X=0.405 $Y=0.216
c31 59 VSS 0.00387072f $X=0.405 $Y=0.207
c32 58 VSS 0.0026043f $X=0.405 $Y=0.116
c33 57 VSS 0.00108941f $X=0.405 $Y=0.063
c34 56 VSS 7.30208e-19 $X=0.405 $Y=0.225
c35 54 VSS 0.00197751f $X=0.3825 $Y=0.036
c36 53 VSS 0.00144534f $X=0.369 $Y=0.036
c37 52 VSS 0.00146498f $X=0.36 $Y=0.036
c38 51 VSS 0.00374035f $X=0.342 $Y=0.036
c39 50 VSS 0.0175638f $X=0.306 $Y=0.036
c40 49 VSS 0.00273151f $X=0.126 $Y=0.036
c41 45 VSS 9.76757e-19 $X=0.099 $Y=0.036
c42 44 VSS 0.00142432f $X=0.09 $Y=0.036
c43 43 VSS 0.00150542f $X=0.072 $Y=0.036
c44 42 VSS 0.00373221f $X=0.063 $Y=0.036
c45 38 VSS 0.00340653f $X=0.036 $Y=0.036
c46 37 VSS 0.00521081f $X=0.396 $Y=0.036
c47 36 VSS 2.98008e-19 $X=0.027 $Y=0.216
c48 34 VSS 3.99179e-19 $X=0.027 $Y=0.07
c49 33 VSS 0.00108941f $X=0.027 $Y=0.063
c50 32 VSS 0.00592912f $X=0.025 $Y=0.111
c51 30 VSS 2.81452e-19 $X=0.027 $Y=0.225
c52 27 VSS 0.00425628f $X=0.376 $Y=0.2025
c53 22 VSS 0.00385394f $X=0.056 $Y=0.2025
c54 19 VSS 4.01171e-19 $X=0.071 $Y=0.2025
c55 12 VSS 0.0066737f $X=0.313 $Y=0.028
c56 6 VSS 0.00670586f $X=0.097 $Y=0.028
r57 74 75 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.4005 $Y2=0.234
r58 73 75 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.234 $X2=0.4005 $Y2=0.234
r59 70 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r60 66 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.045 $Y2=0.234
r61 64 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.045 $Y2=0.234
r62 61 66 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.036 $Y2=0.234
r63 59 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.207 $X2=0.405 $Y2=0.216
r64 58 59 6.17901 $w=1.8e-08 $l=9.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.116 $X2=0.405 $Y2=0.207
r65 57 58 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.063 $X2=0.405 $Y2=0.116
r66 56 73 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.234
r67 56 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.216
r68 55 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.063
r69 53 54 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.369
+ $Y=0.036 $X2=0.3825 $Y2=0.036
r70 52 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.369 $Y2=0.036
r71 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r72 49 50 12.2222 $w=1.8e-08 $l=1.8e-07 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.306 $Y2=0.036
r73 47 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r74 47 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.306 $Y2=0.036
r75 44 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.099 $Y2=0.036
r76 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r77 42 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.036 $X2=0.072 $Y2=0.036
r78 40 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r79 40 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.099 $Y2=0.036
r80 38 42 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.063 $Y2=0.036
r81 37 55 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r82 37 54 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.3825 $Y2=0.036
r83 35 36 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.207 $X2=0.027 $Y2=0.216
r84 33 34 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.063 $X2=0.027 $Y2=0.07
r85 32 35 6.51852 $w=1.8e-08 $l=9.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.111 $X2=0.027 $Y2=0.207
r86 32 34 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.111 $X2=0.027 $Y2=0.07
r87 30 61 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.234
r88 30 36 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.216
r89 29 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r90 29 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.063
r91 27 70 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r92 24 27 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.376 $Y2=0.2025
r93 22 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r94 19 22 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r95 12 47 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r96 9 12 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0455 $X2=0.324 $Y2=0.0455
r97 8 12 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0455 $X2=0.324 $Y2=0.0455
r98 6 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r99 3 6 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0455 $X2=0.108 $Y2=0.0455
r100 2 6 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0455 $X2=0.108 $Y2=0.0455
.ends


* END of "./AOI21x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI21x1_ASAP7_75t_L  VSS VDD B A1 A2 Y
* 
* Y	Y
* A2	A2
* A1	A1
* B	B
M0 N_Y_M0_d N_B_M0_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A1_M1_g noxref_8 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_8 N_A2_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_9 N_A2_M3_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_A1_M4_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 N_Y_M5_d N_B_M5_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341 $Y=0.027
M6 noxref_6 N_B_M6_g N_Y_M6_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 VDD N_A1_M7_g noxref_6 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 noxref_6 N_A2_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 noxref_6 N_A2_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 VDD N_A1_M10_g noxref_6 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 noxref_6 N_B_M11_g N_Y_M11_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "AOI21x1_ASAP7_75t_L.pex.sp.AOI21X1_ASAP7_75T_L.pxi"
* BEGIN of "./AOI21x1_ASAP7_75t_L.pex.sp.AOI21X1_ASAP7_75T_L.pxi"
* File: AOI21x1_ASAP7_75t_L.pex.sp.AOI21X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:10:18 2017
* 
x_PM_AOI21X1_ASAP7_75T_L%B N_B_M0_g N_B_c_3_p N_B_M6_g N_B_M5_g N_B_c_6_p
+ N_B_M11_g B N_B_c_21_p N_B_c_2_p N_B_c_9_p N_B_c_17_p N_B_c_16_p N_B_c_10_p
+ N_B_c_5_p N_B_c_24_p N_B_c_25_p N_B_c_12_p N_B_c_19_p VSS
+ PM_AOI21X1_ASAP7_75T_L%B
x_PM_AOI21X1_ASAP7_75T_L%A1 N_A1_M1_g N_A1_c_39_n N_A1_M7_g N_A1_M4_g
+ N_A1_c_42_n N_A1_M10_g N_A1_c_57_p A1 N_A1_c_68_p N_A1_c_44_n N_A1_c_45_n
+ N_A1_c_46_n N_A1_c_59_p N_A1_c_54_p N_A1_c_47_n N_A1_c_62_p N_A1_c_48_n
+ N_A1_c_63_p VSS PM_AOI21X1_ASAP7_75T_L%A1
x_PM_AOI21X1_ASAP7_75T_L%A2 N_A2_M2_g N_A2_M8_g N_A2_M3_g N_A2_c_87_n N_A2_M9_g
+ A2 VSS PM_AOI21X1_ASAP7_75T_L%A2
x_PM_AOI21X1_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_c_103_n N_Y_M5_d N_Y_M4_d
+ N_Y_c_113_n N_Y_M6_s N_Y_c_104_n N_Y_M11_s N_Y_c_105_n Y N_Y_c_107_n
+ N_Y_c_114_n N_Y_c_109_n N_Y_c_117_n N_Y_c_111_n N_Y_c_124_n N_Y_c_125_n VSS
+ PM_AOI21X1_ASAP7_75T_L%Y
cc_1 N_B_M0_g N_A1_M1_g 0.00354623f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.0675
cc_2 N_B_c_2_p N_A1_M1_g 2.52885e-19 $X=0.163 $Y=0.198 $X2=0.135 $Y2=0.0675
cc_3 N_B_c_3_p N_A1_c_39_n 9.56181e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_B_M5_g N_A1_M4_g 0.00354623f $X=0.351 $Y=0.054 $X2=0.297 $Y2=0.0675
cc_5 N_B_c_5_p N_A1_M4_g 3.05028e-19 $X=0.306 $Y=0.198 $X2=0.297 $Y2=0.0675
cc_6 N_B_c_6_p N_A1_c_42_n 9.56181e-19 $X=0.351 $Y=0.135 $X2=0.297 $Y2=0.135
cc_7 N_B_c_2_p A1 0.00373908f $X=0.163 $Y=0.198 $X2=0.1345 $Y2=0.1355
cc_8 B N_A1_c_44_n 0.00391061f $X=0.0835 $Y=0.1355 $X2=0.144 $Y2=0.072
cc_9 N_B_c_9_p N_A1_c_45_n 2.44969e-19 $X=0.19 $Y=0.198 $X2=0.163 $Y2=0.072
cc_10 N_B_c_10_p N_A1_c_46_n 2.44969e-19 $X=0.288 $Y=0.198 $X2=0.19 $Y2=0.072
cc_11 N_B_c_5_p N_A1_c_47_n 8.29113e-19 $X=0.306 $Y=0.198 $X2=0.297 $Y2=0.134
cc_12 N_B_c_12_p N_A1_c_48_n 0.00146838f $X=0.351 $Y=0.134 $X2=0.297 $Y2=0.125
cc_13 N_B_M0_g N_A2_M2_g 2.63406e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.0675
cc_14 N_B_c_9_p N_A2_M2_g 2.19803e-19 $X=0.19 $Y=0.198 $X2=0.135 $Y2=0.0675
cc_15 N_B_M5_g N_A2_M3_g 2.63406e-19 $X=0.351 $Y=0.054 $X2=0.297 $Y2=0.0675
cc_16 N_B_c_16_p N_A2_M3_g 3.48794e-19 $X=0.256 $Y=0.198 $X2=0.297 $Y2=0.0675
cc_17 N_B_c_17_p A2 0.00368224f $X=0.227 $Y=0.198 $X2=0 $Y2=0
cc_18 N_B_c_16_p A2 9.10799e-19 $X=0.256 $Y=0.198 $X2=0 $Y2=0
cc_19 N_B_c_19_p A2 2.41734e-19 $X=0.351 $Y=0.171 $X2=0 $Y2=0
cc_20 VSS B 5.87812e-19 $X=0.0835 $Y=0.1355 $X2=0.135 $Y2=0.135
cc_21 VSS N_B_c_21_p 0.0016619f $X=0.126 $Y=0.198 $X2=0.135 $Y2=0.135
cc_22 VSS N_B_c_17_p 0.00191933f $X=0.227 $Y=0.198 $X2=0.297 $Y2=0.0675
cc_23 VSS N_B_c_16_p 4.19603e-19 $X=0.256 $Y=0.198 $X2=0.297 $Y2=0.0675
cc_24 VSS N_B_c_24_p 0.00164678f $X=0.333 $Y=0.198 $X2=0.297 $Y2=0.2025
cc_25 VSS N_B_c_25_p 2.08682e-19 $X=0.3375 $Y=0.198 $X2=0.297 $Y2=0.2025
cc_26 VSS N_B_c_19_p 6.39016e-19 $X=0.351 $Y=0.171 $X2=0.297 $Y2=0.2025
cc_27 VSS N_B_c_21_p 0.0195441f $X=0.126 $Y=0.198 $X2=0.1345 $Y2=0.1355
cc_28 B N_Y_c_103_n 0.00127618f $X=0.0835 $Y=0.1355 $X2=0.135 $Y2=0.2025
cc_29 B N_Y_c_104_n 0.00135317f $X=0.0835 $Y=0.1355 $X2=0.135 $Y2=0.099
cc_30 N_B_c_19_p N_Y_c_105_n 0.00135988f $X=0.351 $Y=0.171 $X2=0.163 $Y2=0.072
cc_31 B Y 0.00566958f $X=0.0835 $Y=0.1355 $X2=0.297 $Y2=0.134
cc_32 N_B_M0_g N_Y_c_107_n 2.56935e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_33 B N_Y_c_107_n 0.00123678f $X=0.0835 $Y=0.1355 $X2=0 $Y2=0
cc_34 N_B_M5_g N_Y_c_109_n 3.7308e-19 $X=0.351 $Y=0.054 $X2=0 $Y2=0
cc_35 N_B_c_12_p N_Y_c_109_n 4.52873e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_36 N_B_c_12_p N_Y_c_111_n 0.00369681f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_37 N_A1_M1_g N_A2_M2_g 0.0031831f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_38 N_A1_M4_g N_A2_M2_g 2.34385e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_39 N_A1_c_46_n N_A2_M2_g 2.19803e-19 $X=0.19 $Y=0.072 $X2=0.081 $Y2=0.054
cc_40 N_A1_M1_g N_A2_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.351 $Y2=0.054
cc_41 N_A1_M4_g N_A2_M3_g 0.0031831f $X=0.297 $Y=0.0675 $X2=0.351 $Y2=0.054
cc_42 N_A1_c_54_p N_A2_M3_g 3.45411e-19 $X=0.256 $Y=0.072 $X2=0.351 $Y2=0.054
cc_43 N_A1_c_39_n N_A2_c_87_n 0.0010272f $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.135
cc_44 N_A1_c_42_n N_A2_c_87_n 0.00123834f $X=0.297 $Y=0.135 $X2=0.351 $Y2=0.135
cc_45 N_A1_c_57_p A2 0.00195033f $X=0.135 $Y=0.1165 $X2=0.081 $Y2=0.134
cc_46 A1 A2 0.00126974f $X=0.1345 $Y=0.1355 $X2=0.081 $Y2=0.134
cc_47 N_A1_c_59_p A2 0.00368242f $X=0.227 $Y=0.072 $X2=0.081 $Y2=0.134
cc_48 N_A1_c_54_p A2 9.58063e-19 $X=0.256 $Y=0.072 $X2=0.081 $Y2=0.134
cc_49 N_A1_c_47_n A2 2.10898e-19 $X=0.297 $Y=0.134 $X2=0.081 $Y2=0.134
cc_50 N_A1_c_62_p A2 7.41627e-19 $X=0.297 $Y=0.116 $X2=0.081 $Y2=0.134
cc_51 N_A1_c_63_p A2 8.45393e-19 $X=0.297 $Y=0.1295 $X2=0.081 $Y2=0.134
cc_52 VSS A1 2.75878e-19 $X=0.1345 $Y=0.1355 $X2=0.081 $Y2=0.135
cc_53 VSS N_A1_M1_g 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.18
cc_54 VSS N_A1_M4_g 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.18
cc_55 N_A1_c_44_n N_Y_c_103_n 0.00162967f $X=0.144 $Y=0.072 $X2=0.081 $Y2=0.2025
cc_56 N_A1_c_68_p N_Y_c_113_n 0.00180885f $X=0.288 $Y=0.072 $X2=0.351 $Y2=0.135
cc_57 N_A1_M1_g N_Y_c_114_n 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_A1_M4_g N_Y_c_114_n 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_59 N_A1_c_44_n N_Y_c_114_n 0.016421f $X=0.144 $Y=0.072 $X2=0 $Y2=0
cc_60 N_A1_c_68_p N_Y_c_117_n 6.11332e-19 $X=0.288 $Y=0.072 $X2=0 $Y2=0
cc_61 VSS N_A1_c_68_p 2.44151e-19 $X=0.288 $Y=0.072 $X2=0.081 $Y2=0.054
cc_62 VSS N_A2_c_87_n 3.51308e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_63 VSS N_A2_c_87_n 7.78051e-19 $X=0.243 $Y=0.135 $X2=0.351 $Y2=0.054
cc_64 VSS A2 0.00161796f $X=0.2085 $Y=0.1355 $X2=0.351 $Y2=0.054
cc_65 VSS N_A2_M2_g 2.64781e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.18
cc_66 VSS N_A2_M3_g 2.64781e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.18
cc_67 N_A2_M2_g N_Y_c_114_n 2.64781e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_68 N_A2_M3_g N_Y_c_114_n 2.60867e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_69 VSS N_Y_c_103_n 0.00122706f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.2025
cc_70 VSS N_Y_c_113_n 0.00122706f $X=0.324 $Y=0.2025 $X2=0.351 $Y2=0.135
cc_71 VSS N_Y_c_104_n 0.00379431f $X=0.108 $Y=0.2025 $X2=0.0835 $Y2=0.1355
cc_72 VSS N_Y_c_105_n 0.00363401f $X=0.324 $Y=0.2025 $X2=0.099 $Y2=0.198
cc_73 VSS N_Y_c_124_n 6.57673e-19 $X=0.324 $Y=0.234 $X2=0 $Y2=0
cc_74 VSS N_Y_c_125_n 6.57673e-19 $X=0.324 $Y=0.234 $X2=0 $Y2=0
cc_75 VSS N_Y_c_114_n 2.33741e-19 $X=0.306 $Y=0.036 $X2=0.081 $Y2=0.054
cc_76 VSS N_Y_c_114_n 2.33741e-19 $X=0.306 $Y=0.036 $X2=0.081 $Y2=0.054

* END of "./AOI21x1_ASAP7_75t_L.pex.sp.AOI21X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI21xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:10:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI21xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI21xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI21xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:10:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI21XP33_ASAP7_75T_L%A2 2 5 7 17 19 20 25 VSS
c12 25 VSS 0.0167214f $X=0.0215 $Y=0.1355
c13 20 VSS 5.48708e-19 $X=0.068 $Y=0.134
c14 19 VSS 7.80909e-19 $X=0.055 $Y=0.134
c15 17 VSS 7.04765e-19 $X=0.081 $Y=0.134
c16 5 VSS 0.00333772f $X=0.081 $Y=0.135
c17 2 VSS 0.0653048f $X=0.081 $Y=0.054
r18 19 20 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.055
+ $Y=0.134 $X2=0.068 $Y2=0.134
r19 17 20 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.134 $X2=0.068 $Y2=0.134
r20 15 25 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.134 $X2=0.027 $Y2=0.134
r21 15 19 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.134 $X2=0.055 $Y2=0.134
r22 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.134 $X2=0.081
+ $Y2=0.134
r23 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r24 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI21XP33_ASAP7_75T_L%A1 2 5 7 16 VSS
c13 16 VSS 0.00422246f $X=0.1355 $Y=0.1355
c14 5 VSS 0.00163652f $X=0.135 $Y=0.135
c15 2 VSS 0.0612549f $X=0.135 $Y=0.054
r16 5 16 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.134 $X2=0.135
+ $Y2=0.134
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI21XP33_ASAP7_75T_L%B 2 5 7 10 VSS
c10 10 VSS 0.00169226f $X=0.1865 $Y=0.1355
c11 5 VSS 0.0023144f $X=0.189 $Y=0.135
c12 2 VSS 0.0649588f $X=0.189 $Y=0.054
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.134 $X2=0.189
+ $Y2=0.134
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI21XP33_ASAP7_75T_L%Y 1 2 5 6 9 13 20 25 35 VSS
c14 35 VSS 0.00379235f $X=0.234 $Y=0.234
c15 34 VSS 0.00278493f $X=0.243 $Y=0.234
c16 29 VSS 3.05844e-19 $X=0.243 $Y=0.207
c17 27 VSS 3.96661e-19 $X=0.243 $Y=0.07
c18 26 VSS 0.00104909f $X=0.243 $Y=0.063
c19 25 VSS 0.00588822f $X=0.245 $Y=0.111
c20 23 VSS 0.00102822f $X=0.243 $Y=0.225
c21 21 VSS 3.86697e-19 $X=0.202 $Y=0.036
c22 20 VSS 0.00142432f $X=0.198 $Y=0.036
c23 19 VSS 9.92285e-19 $X=0.18 $Y=0.036
c24 18 VSS 0.0017508f $X=0.171 $Y=0.036
c25 13 VSS 0.00486475f $X=0.162 $Y=0.036
c26 11 VSS 0.00889285f $X=0.234 $Y=0.036
c27 9 VSS 0.00365932f $X=0.214 $Y=0.216
c28 5 VSS 0.00620776f $X=0.162 $Y=0.054
c29 1 VSS 5.3314e-19 $X=0.179 $Y=0.054
r30 35 36 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.2385 $Y2=0.234
r31 34 36 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.234 $X2=0.2385 $Y2=0.234
r32 31 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.234 $Y2=0.234
r33 28 29 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.2 $X2=0.243 $Y2=0.207
r34 26 27 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.063 $X2=0.243 $Y2=0.07
r35 25 28 6.04321 $w=1.8e-08 $l=8.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.111 $X2=0.243 $Y2=0.2
r36 25 27 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.111 $X2=0.243 $Y2=0.07
r37 23 34 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.234
r38 23 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.207
r39 22 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.063
r40 20 21 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.202 $Y2=0.036
r41 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r42 18 19 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.036 $X2=0.18 $Y2=0.036
r43 13 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.171 $Y2=0.036
r44 11 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r45 11 21 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.202 $Y2=0.036
r46 9 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r47 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.216 $X2=0.214 $Y2=0.216
r48 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r49 2 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.054 $X2=0.162 $Y2=0.054
r50 1 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.054 $X2=0.162 $Y2=0.054
.ends


* END of "./AOI21xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI21xp33_ASAP7_75t_L  VSS VDD A2 A1 B Y
* 
* Y	Y
* B	B
* A1	A1
* A2	A2
M0 noxref_8 N_A2_M0_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_Y_M1_d N_A1_M1_g noxref_8 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 VSS N_B_M2_g N_Y_M2_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 VDD N_A2_M3_g noxref_6 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M4 noxref_6 N_A1_M4_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M5 N_Y_M5_d N_B_M5_g noxref_6 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
*
* 
* .include "AOI21xp33_ASAP7_75t_L.pex.sp.AOI21XP33_ASAP7_75T_L.pxi"
* BEGIN of "./AOI21xp33_ASAP7_75t_L.pex.sp.AOI21XP33_ASAP7_75T_L.pxi"
* File: AOI21xp33_ASAP7_75t_L.pex.sp.AOI21XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:10:41 2017
* 
x_PM_AOI21XP33_ASAP7_75T_L%A2 N_A2_M0_g N_A2_c_2_p N_A2_M3_g N_A2_c_3_p
+ N_A2_c_8_p N_A2_c_11_p A2 VSS PM_AOI21XP33_ASAP7_75T_L%A2
x_PM_AOI21XP33_ASAP7_75T_L%A1 N_A1_M1_g N_A1_c_14_n N_A1_M4_g A1 VSS
+ PM_AOI21XP33_ASAP7_75T_L%A1
x_PM_AOI21XP33_ASAP7_75T_L%B N_B_M2_g N_B_c_28_n N_B_M5_g B VSS
+ PM_AOI21XP33_ASAP7_75T_L%B
x_PM_AOI21XP33_ASAP7_75T_L%Y N_Y_M2_s N_Y_M1_d N_Y_c_37_n N_Y_M5_d N_Y_c_41_n
+ N_Y_c_36_n N_Y_c_42_n Y N_Y_c_47_n VSS PM_AOI21XP33_ASAP7_75T_L%Y
cc_1 N_A2_M0_g N_A1_M1_g 0.0031831f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A2_c_2_p N_A1_c_14_n 0.00126427f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A2_c_3_p A1 8.75147e-19 $X=0.081 $Y=0.134 $X2=0.1355 $Y2=0.1355
cc_4 A2 A1 0.00246643f $X=0.0215 $Y=0.1355 $X2=0.1355 $Y2=0.1355
cc_5 N_A2_M0_g N_B_M2_g 2.63406e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_6 VSS A2 2.0764e-19 $X=0.0215 $Y=0.1355 $X2=0.135 $Y2=0.054
cc_7 VSS A2 0.00208864f $X=0.0215 $Y=0.1355 $X2=0.135 $Y2=0.135
cc_8 VSS N_A2_c_8_p 3.7965e-19 $X=0.055 $Y=0.134 $X2=0 $Y2=0
cc_9 VSS A2 0.00170831f $X=0.0215 $Y=0.1355 $X2=0 $Y2=0
cc_10 VSS N_A2_M0_g 4.29887e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_11 VSS N_A2_c_11_p 3.7965e-19 $X=0.068 $Y=0.134 $X2=0 $Y2=0
cc_12 A2 N_Y_c_36_n 5.4399e-19 $X=0.0215 $Y=0.1355 $X2=0.135 $Y2=0.134
cc_13 N_A1_M1_g N_B_M2_g 0.00354623f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_14 N_A1_c_14_n N_B_c_28_n 9.56181e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 A1 B 0.0058998f $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_16 VSS A1 5.77254e-19 $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_17 VSS N_A1_M1_g 2.38303e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_18 VSS A1 0.00377208f $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_19 A1 N_Y_c_37_n 6.66766e-19 $X=0.1355 $Y=0.1355 $X2=0.081 $Y2=0.135
cc_20 N_A1_M1_g N_Y_c_36_n 2.34993e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_21 A1 N_Y_c_36_n 0.00399257f $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_22 VSS B 3.31541e-19 $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_23 B N_Y_c_37_n 3.31541e-19 $X=0.1865 $Y=0.1355 $X2=0.081 $Y2=0.135
cc_24 B N_Y_c_41_n 3.31541e-19 $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_25 N_B_M2_g N_Y_c_42_n 2.56935e-19 $X=0.189 $Y=0.054 $X2=0.068 $Y2=0.134
cc_26 B N_Y_c_42_n 0.00123604f $X=0.1865 $Y=0.1355 $X2=0.068 $Y2=0.134
cc_27 B Y 0.00595614f $X=0.1865 $Y=0.1355 $X2=0.0215 $Y2=0.1355
cc_28 VSS N_Y_c_37_n 6.85003e-19 $X=0.162 $Y=0.216 $X2=0.081 $Y2=0.135
cc_29 VSS N_Y_c_41_n 0.00293888f $X=0.162 $Y=0.216 $X2=0 $Y2=0
cc_30 VSS N_Y_c_47_n 2.53478e-19 $X=0.162 $Y=0.216 $X2=0 $Y2=0
cc_31 VSS N_Y_c_47_n 9.02777e-19 $X=0.162 $Y=0.234 $X2=0 $Y2=0
cc_32 VSS N_Y_c_36_n 2.84666e-19 $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.054

* END of "./AOI21xp33_ASAP7_75t_L.pex.sp.AOI21XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI21xp5_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:11:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI21xp5_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI21xp5_ASAP7_75t_L.pex.sp.pex"
* File: AOI21xp5_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:11:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI21XP5_ASAP7_75T_L%A2 2 5 7 17 19 20 25 VSS
c13 25 VSS 0.018141f $X=0.0215 $Y=0.1355
c14 20 VSS 1.57648e-20 $X=0.053 $Y=0.134
c15 19 VSS 0.00113569f $X=0.052 $Y=0.134
c16 17 VSS 0.001369f $X=0.081 $Y=0.134
c17 5 VSS 0.00343311f $X=0.081 $Y=0.135
c18 2 VSS 0.0653048f $X=0.081 $Y=0.0675
r19 19 20 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.052
+ $Y=0.134 $X2=0.053 $Y2=0.134
r20 17 20 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.134 $X2=0.053 $Y2=0.134
r21 15 25 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.134 $X2=0.018 $Y2=0.134
r22 15 19 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.134 $X2=0.052 $Y2=0.134
r23 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.134 $X2=0.081
+ $Y2=0.134
r24 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r25 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI21XP5_ASAP7_75T_L%A1 2 5 7 16 VSS
c13 16 VSS 0.00491414f $X=0.1355 $Y=0.1355
c14 5 VSS 0.0017472f $X=0.135 $Y=0.135
c15 2 VSS 0.0612549f $X=0.135 $Y=0.0675
r16 5 16 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.134 $X2=0.135
+ $Y2=0.134
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI21XP5_ASAP7_75T_L%B 2 5 7 10 VSS
c10 10 VSS 0.00138458f $X=0.1865 $Y=0.1355
c11 5 VSS 0.00239523f $X=0.189 $Y=0.135
c12 2 VSS 0.0649588f $X=0.189 $Y=0.054
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.134 $X2=0.189
+ $Y2=0.134
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI21XP5_ASAP7_75T_L%Y 2 3 6 10 13 17 24 29 39 VSS
c14 39 VSS 0.00375612f $X=0.234 $Y=0.234
c15 38 VSS 0.00278493f $X=0.243 $Y=0.234
c16 33 VSS 3.05844e-19 $X=0.243 $Y=0.207
c17 31 VSS 3.96661e-19 $X=0.243 $Y=0.07
c18 30 VSS 0.00108941f $X=0.243 $Y=0.063
c19 29 VSS 0.00566596f $X=0.245 $Y=0.111
c20 27 VSS 0.00102822f $X=0.243 $Y=0.225
c21 25 VSS 3.86697e-19 $X=0.202 $Y=0.036
c22 24 VSS 0.00142432f $X=0.198 $Y=0.036
c23 23 VSS 9.16023e-19 $X=0.18 $Y=0.036
c24 22 VSS 0.00178735f $X=0.171 $Y=0.036
c25 17 VSS 0.00474529f $X=0.162 $Y=0.036
c26 15 VSS 0.008388f $X=0.234 $Y=0.036
c27 13 VSS 0.00420068f $X=0.214 $Y=0.2025
c28 6 VSS 0.00684356f $X=0.151 $Y=0.028
r29 39 40 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.2385 $Y2=0.234
r30 38 40 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.234 $X2=0.2385 $Y2=0.234
r31 35 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.234 $Y2=0.234
r32 32 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.2 $X2=0.243 $Y2=0.207
r33 30 31 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.063 $X2=0.243 $Y2=0.07
r34 29 32 6.04321 $w=1.8e-08 $l=8.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.111 $X2=0.243 $Y2=0.2
r35 29 31 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.111 $X2=0.243 $Y2=0.07
r36 27 38 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.234
r37 27 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.207
r38 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.063
r39 24 25 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.202 $Y2=0.036
r40 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r41 22 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.036 $X2=0.18 $Y2=0.036
r42 17 22 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.171 $Y2=0.036
r43 15 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r44 15 25 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.202 $Y2=0.036
r45 13 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r46 10 13 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.214 $Y2=0.2025
r47 6 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r48 3 6 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.0455 $X2=0.162 $Y2=0.0455
r49 2 6 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0455 $X2=0.162 $Y2=0.0455
.ends


* END of "./AOI21xp5_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI21xp5_ASAP7_75t_L  VSS VDD A2 A1 B Y
* 
* Y	Y
* B	B
* A1	A1
* A2	A2
M0 noxref_8 N_A2_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_Y_M1_d N_A1_M1_g noxref_8 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_B_M2_g N_Y_M2_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 VDD N_A2_M3_g noxref_6 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M4 noxref_6 N_A1_M4_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M5 N_Y_M5_d N_B_M5_g noxref_6 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
*
* 
* .include "AOI21xp5_ASAP7_75t_L.pex.sp.AOI21XP5_ASAP7_75T_L.pxi"
* BEGIN of "./AOI21xp5_ASAP7_75t_L.pex.sp.AOI21XP5_ASAP7_75T_L.pxi"
* File: AOI21xp5_ASAP7_75t_L.pex.sp.AOI21XP5_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:11:03 2017
* 
x_PM_AOI21XP5_ASAP7_75T_L%A2 N_A2_M0_g N_A2_c_2_p N_A2_M3_g N_A2_c_3_p
+ N_A2_c_8_p N_A2_c_9_p A2 VSS PM_AOI21XP5_ASAP7_75T_L%A2
x_PM_AOI21XP5_ASAP7_75T_L%A1 N_A1_M1_g N_A1_c_15_n N_A1_M4_g A1 VSS
+ PM_AOI21XP5_ASAP7_75T_L%A1
x_PM_AOI21XP5_ASAP7_75T_L%B N_B_M2_g N_B_c_29_n N_B_M5_g B VSS
+ PM_AOI21XP5_ASAP7_75T_L%B
x_PM_AOI21XP5_ASAP7_75T_L%Y N_Y_M2_s N_Y_M1_d N_Y_c_38_n N_Y_M5_d N_Y_c_42_n
+ N_Y_c_37_n N_Y_c_43_n Y N_Y_c_48_n VSS PM_AOI21XP5_ASAP7_75T_L%Y
cc_1 N_A2_M0_g N_A1_M1_g 0.0031831f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A2_c_2_p N_A1_c_15_n 0.00126818f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A2_c_3_p A1 8.76965e-19 $X=0.081 $Y=0.134 $X2=0.1355 $Y2=0.1355
cc_4 A2 A1 0.00162822f $X=0.0215 $Y=0.1355 $X2=0.1355 $Y2=0.1355
cc_5 N_A2_M0_g N_B_M2_g 2.63406e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 VSS A2 2.23359e-19 $X=0.0215 $Y=0.1355 $X2=0.135 $Y2=0.0675
cc_7 VSS A2 0.00234739f $X=0.0215 $Y=0.1355 $X2=0.135 $Y2=0.135
cc_8 VSS N_A2_c_8_p 2.61145e-19 $X=0.052 $Y=0.134 $X2=0.135 $Y2=0.134
cc_9 VSS N_A2_c_9_p 2.61145e-19 $X=0.053 $Y=0.134 $X2=0.135 $Y2=0.134
cc_10 VSS A2 0.00147537f $X=0.0215 $Y=0.1355 $X2=0.135 $Y2=0.134
cc_11 VSS N_A2_M0_g 4.29887e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_12 VSS N_A2_c_3_p 2.61145e-19 $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_13 A2 N_Y_c_37_n 5.25878e-19 $X=0.0215 $Y=0.1355 $X2=0 $Y2=0
cc_14 N_A1_M1_g N_B_M2_g 0.00354623f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_15 N_A1_c_15_n N_B_c_29_n 9.56181e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_16 A1 B 0.00491377f $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_17 VSS A1 0.00137761f $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_18 VSS N_A1_M1_g 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 VSS A1 0.00375081f $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_20 A1 N_Y_c_38_n 0.00161209f $X=0.1355 $Y=0.1355 $X2=0.081 $Y2=0.2025
cc_21 N_A1_M1_g N_Y_c_37_n 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.134
cc_22 A1 N_Y_c_37_n 0.00399256f $X=0.1355 $Y=0.1355 $X2=0.081 $Y2=0.134
cc_23 VSS B 0.00114532f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_24 B N_Y_c_38_n 0.00127618f $X=0.1865 $Y=0.1355 $X2=0.081 $Y2=0.2025
cc_25 B N_Y_c_42_n 0.00114532f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_26 N_B_M2_g N_Y_c_43_n 2.56935e-19 $X=0.189 $Y=0.054 $X2=0.018 $Y2=0.134
cc_27 B N_Y_c_43_n 0.00123604f $X=0.1865 $Y=0.1355 $X2=0.018 $Y2=0.134
cc_28 B Y 0.00542605f $X=0.1865 $Y=0.1355 $X2=0 $Y2=0
cc_29 VSS N_Y_c_38_n 0.00107253f $X=0.162 $Y=0.2025 $X2=0.081 $Y2=0.2025
cc_30 VSS N_Y_c_42_n 0.0040698f $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_31 VSS N_Y_c_48_n 2.53478e-19 $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_32 VSS N_Y_c_48_n 9.02777e-19 $X=0.162 $Y=0.234 $X2=0 $Y2=0
cc_33 VSS N_Y_c_37_n 2.78119e-19 $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.0675

* END of "./AOI21xp5_ASAP7_75t_L.pex.sp.AOI21XP5_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI221x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:11:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI221x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI221x1_ASAP7_75t_L.pex.sp.pex"
* File: AOI221x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:11:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI221X1_ASAP7_75T_L%A2 2 7 10 13 19 21 VSS
c14 21 VSS 8.38057e-19 $X=0.135 $Y=0.135
c15 19 VSS 0.0118282f $X=0.1035 $Y=0.1365
c16 10 VSS 0.0676656f $X=0.135 $Y=0.1345
c17 2 VSS 0.063392f $X=0.081 $Y=0.0675
r18 19 21 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.1035
+ $Y=0.135 $X2=0.135 $Y2=0.135
r19 10 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r20 10 13 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1345 $X2=0.135 $Y2=0.2025
r21 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1345 $X2=0.135 $Y2=0.1345
r22 5 7 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1345 $X2=0.081 $Y2=0.2025
r23 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.1345
.ends

.subckt PM_AOI221X1_ASAP7_75T_L%A1 2 5 8 11 13 18 22 25 VSS
c22 25 VSS 1.97014e-19 $X=0.189 $Y=0.1305
c23 22 VSS 0.00223404f $X=0.189 $Y=0.135
c24 18 VSS 0.00570545f $X=0.187 $Y=0.081
c25 11 VSS 0.00617017f $X=0.243 $Y=0.1345
c26 8 VSS 0.0617105f $X=0.243 $Y=0.0675
c27 2 VSS 0.0593999f $X=0.189 $Y=0.1345
r28 24 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.1305
r29 22 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.1305
r30 18 24 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.081 $X2=0.189 $Y2=0.126
r31 11 13 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1345 $X2=0.243 $Y2=0.2025
r32 8 11 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.1345
r33 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.1345 $X2=0.243 $Y2=0.1345
r34 2 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r35 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1345 $X2=0.189 $Y2=0.2025
.ends

.subckt PM_AOI221X1_ASAP7_75T_L%B1 2 7 10 13 18 20 23 VSS
c30 23 VSS 1.82154e-19 $X=0.297 $Y=0.1305
c31 20 VSS 0.00125985f $X=0.297 $Y=0.135
c32 18 VSS 9.80015e-19 $X=0.2955 $Y=0.1165
c33 10 VSS 0.0643808f $X=0.351 $Y=0.1345
c34 2 VSS 0.0606561f $X=0.297 $Y=0.0675
r35 22 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.1305
r36 20 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.1305
r37 18 22 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1165 $X2=0.297 $Y2=0.126
r38 10 13 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.1345 $X2=0.351 $Y2=0.2025
r39 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.1345 $X2=0.351 $Y2=0.1345
r40 5 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r41 5 7 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.1345 $X2=0.297 $Y2=0.2025
r42 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.1345
.ends

.subckt PM_AOI221X1_ASAP7_75T_L%B2 2 5 8 11 13 20 26 28 VSS
c27 26 VSS 0.00231068f $X=0.468 $Y=0.135
c28 20 VSS 5.28708e-19 $X=0.431 $Y=0.135
c29 11 VSS 0.0043293f $X=0.459 $Y=0.1345
c30 8 VSS 0.0636211f $X=0.459 $Y=0.0675
c31 2 VSS 0.0618739f $X=0.405 $Y=0.1345
r32 26 28 0.83878 $w=2.55e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.135 $X2=0.468 $Y2=0.1525
r33 20 21 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.135 $X2=0.4405 $Y2=0.135
r34 17 20 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.431 $Y2=0.135
r35 15 26 0.278257 $w=2.55e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.135 $X2=0.468 $Y2=0.135
r36 15 21 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.135 $X2=0.4405 $Y2=0.135
r37 11 13 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.1345 $X2=0.459 $Y2=0.2025
r38 8 11 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.1345
r39 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.1345 $X2=0.459 $Y2=0.1345
r40 2 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r41 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.1345 $X2=0.405 $Y2=0.2025
.ends

.subckt PM_AOI221X1_ASAP7_75T_L%C 2 7 10 13 20 22 25 33 VSS
c23 33 VSS 0.0029575f $X=0.567 $Y=0.135
c24 25 VSS 0.00110768f $X=0.621 $Y=0.135
c25 22 VSS 5.84898e-19 $X=0.567 $Y=0.171
c26 21 VSS 4.35275e-19 $X=0.567 $Y=0.153
c27 20 VSS 0.00122901f $X=0.571 $Y=0.1885
c28 10 VSS 0.0723308f $X=0.675 $Y=0.1345
c29 2 VSS 0.0654137f $X=0.621 $Y=0.054
r30 23 33 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.135 $X2=0.567 $Y2=0.135
r31 23 25 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.135 $X2=0.621 $Y2=0.135
r32 21 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.153 $X2=0.567 $Y2=0.171
r33 20 22 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.1885 $X2=0.567 $Y2=0.171
r34 17 33 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.144 $X2=0.567 $Y2=0.135
r35 17 21 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.144 $X2=0.567 $Y2=0.153
r36 10 13 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.1345 $X2=0.675 $Y2=0.2025
r37 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621
+ $Y=0.1345 $X2=0.675 $Y2=0.1345
r38 5 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r39 5 7 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.1345 $X2=0.621 $Y2=0.2025
r40 2 5 301.593 $w=2e-08 $l=8.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.054 $X2=0.621 $Y2=0.1345
.ends

.subckt PM_AOI221X1_ASAP7_75T_L%Y 1 2 5 6 9 11 12 15 18 26 27 28 29 30 31 34 35
+ 36 37 40 45 50 52 54 VSS
c44 54 VSS 0.00131807f $X=0.729 $Y=0.1665
c45 52 VSS 0.00266121f $X=0.729 $Y=0.126
c46 51 VSS 0.00104959f $X=0.729 $Y=0.081
c47 50 VSS 7.73365e-19 $X=0.7305 $Y=0.1335
c48 48 VSS 0.00115971f $X=0.729 $Y=0.189
c49 46 VSS 1.40401e-19 $X=0.718 $Y=0.198
c50 45 VSS 5.10798e-19 $X=0.716 $Y=0.198
c51 40 VSS 1.07894e-19 $X=0.648 $Y=0.198
c52 38 VSS 0.00199737f $X=0.72 $Y=0.198
c53 37 VSS 0.00523334f $X=0.678 $Y=0.054
c54 36 VSS 0.00230531f $X=0.636 $Y=0.054
c55 35 VSS 6.11608e-19 $X=0.585 $Y=0.054
c56 34 VSS 0.00220631f $X=0.576 $Y=0.054
c57 33 VSS 0.00355372f $X=0.539 $Y=0.054
c58 32 VSS 0.00285603f $X=0.5 $Y=0.054
c59 31 VSS 0.00241564f $X=0.487 $Y=0.054
c60 30 VSS 0.00153912f $X=0.468 $Y=0.054
c61 29 VSS 0.0020516f $X=0.431 $Y=0.054
c62 28 VSS 0.00395673f $X=0.391 $Y=0.054
c63 27 VSS 0.00156238f $X=0.325 $Y=0.054
c64 26 VSS 8.77986e-19 $X=0.288 $Y=0.054
c65 18 VSS 0.00122401f $X=0.27 $Y=0.054
c66 16 VSS 0.00554217f $X=0.72 $Y=0.054
c67 15 VSS 0.00374804f $X=0.648 $Y=0.2025
c68 11 VSS 5.71486e-19 $X=0.665 $Y=0.2025
c69 9 VSS 0.00439245f $X=0.596 $Y=0.054
c70 6 VSS 3.29654e-19 $X=0.611 $Y=0.054
c71 5 VSS 7.50005e-19 $X=0.27 $Y=0.0675
c72 1 VSS 7.79082e-19 $X=0.287 $Y=0.0675
r73 53 54 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.144 $X2=0.729 $Y2=0.1665
r74 51 52 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.081 $X2=0.729 $Y2=0.126
r75 50 53 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.1335 $X2=0.729 $Y2=0.144
r76 50 52 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.1335 $X2=0.729 $Y2=0.126
r77 48 54 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.189 $X2=0.729 $Y2=0.1665
r78 47 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.063 $X2=0.729 $Y2=0.081
r79 45 46 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.716
+ $Y=0.198 $X2=0.718 $Y2=0.198
r80 40 45 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.198 $X2=0.716 $Y2=0.198
r81 38 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.198 $X2=0.729 $Y2=0.189
r82 38 46 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.198 $X2=0.718 $Y2=0.198
r83 36 37 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.636
+ $Y=0.054 $X2=0.678 $Y2=0.054
r84 34 35 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.054 $X2=0.585 $Y2=0.054
r85 33 34 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.539
+ $Y=0.054 $X2=0.576 $Y2=0.054
r86 32 33 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5
+ $Y=0.054 $X2=0.539 $Y2=0.054
r87 31 32 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.487
+ $Y=0.054 $X2=0.5 $Y2=0.054
r88 30 31 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.054 $X2=0.487 $Y2=0.054
r89 29 30 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.054 $X2=0.468 $Y2=0.054
r90 28 29 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.391
+ $Y=0.054 $X2=0.431 $Y2=0.054
r91 27 28 4.48148 $w=1.8e-08 $l=6.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.325
+ $Y=0.054 $X2=0.391 $Y2=0.054
r92 26 27 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.054 $X2=0.325 $Y2=0.054
r93 24 36 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.054 $X2=0.636 $Y2=0.054
r94 24 35 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.054 $X2=0.585 $Y2=0.054
r95 18 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.054 $X2=0.288 $Y2=0.054
r96 16 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.054 $X2=0.729 $Y2=0.063
r97 16 37 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.054 $X2=0.678 $Y2=0.054
r98 15 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.198 $X2=0.648
+ $Y2=0.198
r99 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.648 $Y2=0.2025
r100 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.648 $Y2=0.2025
r101 9 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.054 $X2=0.594
+ $Y2=0.054
r102 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.054 $X2=0.596 $Y2=0.054
r103 5 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.054 $X2=0.27
+ $Y2=0.054
r104 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r105 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends


* END of "./AOI221x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI221x1_ASAP7_75t_L  VSS VDD A2 A1 B1 B2 C Y
* 
* Y	Y
* C	C
* B2	B2
* B1	B1
* A1	A1
* A2	A2
M0 noxref_11 N_A2_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_Y_M1_d N_A1_M1_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M2 noxref_12 N_B1_M2_g N_Y_M2_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 VSS N_B2_M3_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M4 VSS N_C_M4_g N_Y_M4_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.611 $Y=0.027
M5 VDD N_A2_M5_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M6 VDD N_A2_M6_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 VDD N_A1_M7_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M8 VDD N_A1_M8_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M9 noxref_9 N_B1_M9_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M10 noxref_9 N_B1_M10_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M11 noxref_9 N_B2_M11_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M12 noxref_9 N_B2_M12_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M13 N_Y_M13_d N_C_M13_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M14 N_Y_M14_d N_C_M14_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
*
* 
* .include "AOI221x1_ASAP7_75t_L.pex.sp.AOI221X1_ASAP7_75T_L.pxi"
* BEGIN of "./AOI221x1_ASAP7_75t_L.pex.sp.AOI221X1_ASAP7_75T_L.pxi"
* File: AOI221x1_ASAP7_75t_L.pex.sp.AOI221X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:11:25 2017
* 
x_PM_AOI221X1_ASAP7_75T_L%A2 N_A2_M0_g N_A2_M5_g N_A2_c_2_p N_A2_M6_g A2
+ N_A2_c_7_p VSS PM_AOI221X1_ASAP7_75T_L%A2
x_PM_AOI221X1_ASAP7_75T_L%A1 N_A1_c_15_n N_A1_M7_g N_A1_M1_g N_A1_c_18_n
+ N_A1_M8_g A1 N_A1_c_20_n N_A1_c_21_n VSS PM_AOI221X1_ASAP7_75T_L%A1
x_PM_AOI221X1_ASAP7_75T_L%B1 N_B1_M2_g N_B1_M9_g N_B1_c_39_n N_B1_M10_g B1
+ N_B1_c_41_n N_B1_c_46_p VSS PM_AOI221X1_ASAP7_75T_L%B1
x_PM_AOI221X1_ASAP7_75T_L%B2 N_B2_c_67_n N_B2_M11_g N_B2_M3_g N_B2_c_70_n
+ N_B2_M12_g N_B2_c_71_n N_B2_c_72_n B2 VSS PM_AOI221X1_ASAP7_75T_L%B2
x_PM_AOI221X1_ASAP7_75T_L%C N_C_M4_g N_C_M13_g N_C_c_101_p N_C_M14_g C
+ N_C_c_94_n N_C_c_100_p N_C_c_95_n VSS PM_AOI221X1_ASAP7_75T_L%C
x_PM_AOI221X1_ASAP7_75T_L%Y N_Y_M2_s N_Y_M1_d N_Y_c_118_n N_Y_M4_s N_Y_c_143_n
+ N_Y_M14_d N_Y_M13_d N_Y_c_129_n N_Y_c_117_n N_Y_c_119_n N_Y_c_120_n
+ N_Y_c_122_n N_Y_c_123_n N_Y_c_125_n N_Y_c_127_n N_Y_c_130_n N_Y_c_131_n
+ N_Y_c_132_n N_Y_c_135_n N_Y_c_136_n N_Y_c_138_n Y N_Y_c_140_n N_Y_c_151_n VSS
+ PM_AOI221X1_ASAP7_75T_L%Y
cc_1 N_A2_M0_g N_A1_c_15_n 2.48122e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.1345
cc_2 N_A2_c_2_p N_A1_c_15_n 0.00335986f $X=0.135 $Y=0.1345 $X2=0.189 $Y2=0.1345
cc_3 N_A2_c_2_p N_A1_M1_g 2.53865e-19 $X=0.135 $Y=0.1345 $X2=0.243 $Y2=0.0675
cc_4 N_A2_c_2_p N_A1_c_18_n 0.00121867f $X=0.135 $Y=0.1345 $X2=0.243 $Y2=0.1345
cc_5 A2 A1 0.00134782f $X=0.1035 $Y=0.1365 $X2=0.187 $Y2=0.081
cc_6 A2 N_A1_c_20_n 4.36364e-19 $X=0.1035 $Y=0.1365 $X2=0.189 $Y2=0.135
cc_7 N_A2_c_7_p N_A1_c_21_n 8.75147e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.1305
cc_8 VSS A2 0.00124033f $X=0.1035 $Y=0.1365 $X2=0.189 $Y2=0.2025
cc_9 VSS N_A2_M0_g 3.37932e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_10 VSS A2 0.0037268f $X=0.1035 $Y=0.1365 $X2=0 $Y2=0
cc_11 VSS N_A2_c_2_p 6.72287e-19 $X=0.135 $Y=0.1345 $X2=0 $Y2=0
cc_12 VSS N_A2_c_7_p 0.0016731f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_13 VSS A2 0.00272629f $X=0.1035 $Y=0.1365 $X2=0 $Y2=0
cc_14 VSS N_A2_c_2_p 0.00283759f $X=0.135 $Y=0.1345 $X2=0.243 $Y2=0.1345
cc_15 N_A1_c_15_n N_B1_M2_g 2.53865e-19 $X=0.189 $Y=0.1345 $X2=0.081 $Y2=0.0675
cc_16 N_A1_M1_g N_B1_M2_g 0.00353416f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 N_A1_M1_g N_B1_c_39_n 2.88628e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.1345
cc_18 N_A1_c_18_n N_B1_c_39_n 0.00136604f $X=0.243 $Y=0.1345 $X2=0.135
+ $Y2=0.1345
cc_19 N_A1_c_20_n N_B1_c_41_n 5.64422e-19 $X=0.189 $Y=0.135 $X2=0.135 $Y2=0.135
cc_20 VSS N_A1_c_20_n 3.18961e-19 $X=0.189 $Y=0.135 $X2=0.135 $Y2=0.1345
cc_21 VSS N_A1_c_15_n 3.42691e-19 $X=0.189 $Y=0.1345 $X2=0 $Y2=0
cc_22 VSS N_A1_c_20_n 0.00376061f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_23 VSS N_A1_M1_g 4.8541e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_24 VSS N_A1_c_18_n 7.80906e-19 $X=0.243 $Y=0.1345 $X2=0 $Y2=0
cc_25 A1 N_Y_c_117_n 3.8748e-19 $X=0.187 $Y=0.081 $X2=0.1035 $Y2=0.135
cc_26 VSS A1 5.62512e-19 $X=0.187 $Y=0.081 $X2=0.081 $Y2=0.2025
cc_27 VSS N_A1_c_15_n 0.00180933f $X=0.189 $Y=0.1345 $X2=0 $Y2=0
cc_28 VSS N_A1_c_18_n 0.00123462f $X=0.243 $Y=0.1345 $X2=0 $Y2=0
cc_29 VSS A1 0.00538014f $X=0.187 $Y=0.081 $X2=0 $Y2=0
cc_30 N_B1_M2_g N_B2_c_67_n 2.94371e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.1345
cc_31 N_B1_c_39_n N_B2_c_67_n 0.00360681f $X=0.351 $Y=0.1345 $X2=0.189
+ $Y2=0.1345
cc_32 N_B1_c_39_n N_B2_M3_g 2.88628e-19 $X=0.351 $Y=0.1345 $X2=0.243 $Y2=0.0675
cc_33 N_B1_c_39_n N_B2_c_70_n 0.00129516f $X=0.351 $Y=0.1345 $X2=0.243
+ $Y2=0.1345
cc_34 N_B1_c_46_p N_B2_c_71_n 3.36034e-19 $X=0.297 $Y=0.1305 $X2=0 $Y2=0
cc_35 B1 N_B2_c_72_n 4.25612e-19 $X=0.2955 $Y=0.1165 $X2=0 $Y2=0
cc_36 N_B1_c_41_n N_B2_c_72_n 2.36455e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_37 VSS N_B1_c_41_n 9.17001e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_38 VSS N_B1_M2_g 3.37932e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_39 VSS N_B1_c_41_n 0.00373387f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_40 VSS N_B1_c_39_n 8.10164e-19 $X=0.351 $Y=0.1345 $X2=0 $Y2=0
cc_41 VSS N_B1_c_39_n 2.10893e-19 $X=0.351 $Y=0.1345 $X2=0 $Y2=0
cc_42 VSS N_B1_c_39_n 3.77106e-19 $X=0.351 $Y=0.1345 $X2=0.189 $Y2=0.1345
cc_43 VSS N_B1_c_39_n 7.79752e-19 $X=0.351 $Y=0.1345 $X2=0.189 $Y2=0.2025
cc_44 VSS N_B1_c_41_n 3.21662e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_45 VSS N_B1_c_39_n 2.64905e-19 $X=0.351 $Y=0.1345 $X2=0 $Y2=0
cc_46 B1 N_Y_c_118_n 9.43494e-19 $X=0.2955 $Y=0.1165 $X2=0.189 $Y2=0.2025
cc_47 N_B1_c_41_n N_Y_c_119_n 3.25138e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_48 N_B1_M2_g N_Y_c_120_n 2.94721e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_49 B1 N_Y_c_120_n 0.00376017f $X=0.2955 $Y=0.1165 $X2=0 $Y2=0
cc_50 N_B1_c_39_n N_Y_c_122_n 7.88415e-19 $X=0.351 $Y=0.1345 $X2=0 $Y2=0
cc_51 VSS N_B1_c_39_n 0.00284027f $X=0.351 $Y=0.1345 $X2=0.189 $Y2=0.1345
cc_52 VSS N_B1_c_39_n 0.00322695f $X=0.351 $Y=0.1345 $X2=0.189 $Y2=0.1345
cc_53 VSS B1 0.00215266f $X=0.2955 $Y=0.1165 $X2=0.189 $Y2=0.1345
cc_54 VSS N_B1_c_39_n 2.13371e-19 $X=0.351 $Y=0.1345 $X2=0.243 $Y2=0.0675
cc_55 N_B2_c_72_n N_C_c_94_n 4.27572e-19 $X=0.468 $Y=0.135 $X2=0.297 $Y2=0.126
cc_56 N_B2_c_72_n N_C_c_95_n 0.00118005f $X=0.468 $Y=0.135 $X2=0 $Y2=0
cc_57 VSS N_B2_c_72_n 9.62431e-19 $X=0.468 $Y=0.135 $X2=0 $Y2=0
cc_58 VSS N_B2_M3_g 2.5328e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_59 VSS N_B2_c_72_n 0.00373387f $X=0.468 $Y=0.135 $X2=0 $Y2=0
cc_60 VSS N_B2_c_67_n 3.32571e-19 $X=0.405 $Y=0.1345 $X2=0 $Y2=0
cc_61 VSS N_B2_c_70_n 2.44334e-19 $X=0.459 $Y=0.1345 $X2=0 $Y2=0
cc_62 VSS N_B2_c_71_n 0.00166652f $X=0.431 $Y=0.135 $X2=0 $Y2=0
cc_63 VSS N_B2_c_70_n 3.77535e-19 $X=0.459 $Y=0.1345 $X2=0.297 $Y2=0.2025
cc_64 VSS N_B2_c_72_n 3.21662e-19 $X=0.468 $Y=0.135 $X2=0.351 $Y2=0.1345
cc_65 VSS N_B2_c_67_n 2.64905e-19 $X=0.405 $Y=0.1345 $X2=0 $Y2=0
cc_66 VSS N_B2_M3_g 2.38414e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_67 N_B2_c_67_n N_Y_c_123_n 3.63954e-19 $X=0.405 $Y=0.1345 $X2=0 $Y2=0
cc_68 N_B2_c_71_n N_Y_c_123_n 6.46728e-19 $X=0.431 $Y=0.135 $X2=0 $Y2=0
cc_69 N_B2_M3_g N_Y_c_125_n 2.90628e-19 $X=0.459 $Y=0.0675 $X2=0.297 $Y2=0.1345
cc_70 N_B2_c_72_n N_Y_c_125_n 0.00373901f $X=0.468 $Y=0.135 $X2=0.297 $Y2=0.1345
cc_71 N_B2_c_72_n N_Y_c_127_n 3.3127e-19 $X=0.468 $Y=0.135 $X2=0 $Y2=0
cc_72 VSS N_B2_c_67_n 0.00284008f $X=0.405 $Y=0.1345 $X2=0.297 $Y2=0.0675
cc_73 VSS N_B2_c_72_n 0.00207431f $X=0.468 $Y=0.135 $X2=0.297 $Y2=0.0675
cc_74 VSS N_B2_c_70_n 2.1361e-19 $X=0.459 $Y=0.1345 $X2=0.351 $Y2=0.1345
cc_75 VSS N_C_c_94_n 3.59874e-19 $X=0.567 $Y=0.171 $X2=0 $Y2=0
cc_76 VSS C 9.35091e-19 $X=0.571 $Y=0.1885 $X2=0 $Y2=0
cc_77 VSS N_C_c_94_n 0.00148695f $X=0.567 $Y=0.171 $X2=0 $Y2=0
cc_78 VSS C 0.00372728f $X=0.571 $Y=0.1885 $X2=0 $Y2=0
cc_79 VSS N_C_c_100_p 0.00105872f $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_80 VSS N_C_c_101_p 2.21858e-19 $X=0.675 $Y=0.1345 $X2=0 $Y2=0
cc_81 VSS N_C_M4_g 4.29408e-19 $X=0.621 $Y=0.054 $X2=0 $Y2=0
cc_82 N_C_c_101_p N_Y_M14_d 3.77145e-19 $X=0.675 $Y=0.1345 $X2=0.459 $Y2=0.1345
cc_83 N_C_c_101_p N_Y_c_129_n 8.94806e-19 $X=0.675 $Y=0.1345 $X2=0.45 $Y2=0.135
cc_84 N_C_c_95_n N_Y_c_130_n 0.0037574f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_85 N_C_c_100_p N_Y_c_131_n 7.12585e-19 $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_86 N_C_M4_g N_Y_c_132_n 4.1691e-19 $X=0.621 $Y=0.054 $X2=0 $Y2=0
cc_87 N_C_c_101_p N_Y_c_132_n 9.19156e-19 $X=0.675 $Y=0.1345 $X2=0 $Y2=0
cc_88 N_C_c_100_p N_Y_c_132_n 7.12585e-19 $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_89 N_C_c_101_p N_Y_c_135_n 3.11627e-19 $X=0.675 $Y=0.1345 $X2=0 $Y2=0
cc_90 N_C_c_101_p N_Y_c_136_n 7.49672e-19 $X=0.675 $Y=0.1345 $X2=0 $Y2=0
cc_91 C N_Y_c_136_n 3.66377e-19 $X=0.571 $Y=0.1885 $X2=0 $Y2=0
cc_92 N_C_c_101_p N_Y_c_138_n 3.97853e-19 $X=0.675 $Y=0.1345 $X2=0 $Y2=0
cc_93 N_C_c_100_p Y 2.33843e-19 $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_94 N_C_c_101_p N_Y_c_140_n 5.00201e-19 $X=0.675 $Y=0.1345 $X2=0 $Y2=0
cc_95 N_C_c_95_n N_Y_c_140_n 5.26187e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_96 VSS N_Y_c_118_n 0.00117451f $X=0.27 $Y=0.2025 $X2=0.081 $Y2=0.1345
cc_97 VSS N_Y_c_143_n 8.7738e-19 $X=0.596 $Y=0.2025 $X2=0.351 $Y2=0.1345
cc_98 VSS N_Y_c_129_n 0.00374846f $X=0.596 $Y=0.2025 $X2=0 $Y2=0
cc_99 VSS N_Y_c_129_n 0.00368895f $X=0.7 $Y=0.2025 $X2=0 $Y2=0
cc_100 VSS N_Y_c_129_n 0.0025501f $X=0.668 $Y=0.234 $X2=0 $Y2=0
cc_101 VSS N_Y_c_136_n 3.96143e-19 $X=0.596 $Y=0.2025 $X2=0 $Y2=0
cc_102 VSS N_Y_c_136_n 0.00353151f $X=0.702 $Y=0.234 $X2=0 $Y2=0
cc_103 VSS N_Y_c_136_n 0.00353151f $X=0.668 $Y=0.234 $X2=0 $Y2=0
cc_104 VSS N_Y_c_138_n 0.00281841f $X=0.7 $Y=0.2025 $X2=0 $Y2=0
cc_105 VSS N_Y_c_151_n 3.50898e-19 $X=0.7 $Y=0.2025 $X2=0 $Y2=0
cc_106 VSS N_Y_c_118_n 0.0039137f $X=0.27 $Y=0.0675 $X2=0.243 $Y2=0.1345
cc_107 VSS N_Y_c_117_n 4.2769e-19 $X=0.27 $Y=0.054 $X2=0.243 $Y2=0.1345
cc_108 VSS N_Y_c_122_n 0.00211877f $X=0.391 $Y=0.054 $X2=0.189 $Y2=0.1345
cc_109 VSS N_Y_c_118_n 0.00316448f $X=0.27 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_110 VSS N_Y_c_120_n 0.00107451f $X=0.325 $Y=0.054 $X2=0.243 $Y2=0.0675
cc_111 VSS N_Y_c_122_n 0.00159956f $X=0.391 $Y=0.054 $X2=0.243 $Y2=0.0675
cc_112 VSS N_Y_c_123_n 2.87556e-19 $X=0.431 $Y=0.054 $X2=0.243 $Y2=0.1345
cc_113 VSS N_Y_c_123_n 0.00133661f $X=0.431 $Y=0.054 $X2=0.243 $Y2=0.2025
cc_114 VSS N_Y_c_125_n 0.00106132f $X=0.468 $Y=0.054 $X2=0.243 $Y2=0.2025

* END of "./AOI221x1_ASAP7_75t_L.pex.sp.AOI221X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI221xp5_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:11:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI221xp5_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI221xp5_ASAP7_75t_L.pex.sp.pex"
* File: AOI221xp5_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:11:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI221XP5_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c11 10 VSS 6.95749e-19 $X=0.081 $Y=0.135
c12 5 VSS 0.00170784f $X=0.081 $Y=0.135
c13 2 VSS 0.0655264f $X=0.081 $Y=0.054
r14 10 14 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.148
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI221XP5_ASAP7_75T_L%B2 2 5 7 10 VSS
c11 10 VSS 0.00105185f $X=0.134 $Y=0.109
c12 5 VSS 0.00113686f $X=0.135 $Y=0.135
c13 2 VSS 0.0607092f $X=0.135 $Y=0.054
r14 10 13 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.109 $X2=0.135 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI221XP5_ASAP7_75T_L%C 2 5 7 10 VSS
c11 10 VSS 0.00138457f $X=0.188 $Y=0.123
c12 5 VSS 0.00120113f $X=0.189 $Y=0.135
c13 2 VSS 0.0599046f $X=0.189 $Y=0.054
r14 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.123 $X2=0.189 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI221XP5_ASAP7_75T_L%A1 2 5 7 10 VSS
c10 10 VSS 0.00122183f $X=0.24 $Y=0.09
c11 5 VSS 0.00124202f $X=0.243 $Y=0.135
c12 2 VSS 0.0597675f $X=0.243 $Y=0.054
r13 10 13 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.09 $X2=0.243 $Y2=0.135
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI221XP5_ASAP7_75T_L%A2 2 5 7 10 VSS
c8 10 VSS 0.00516661f $X=0.295 $Y=0.123
c9 5 VSS 0.00230503f $X=0.297 $Y=0.135
c10 2 VSS 0.0631596f $X=0.297 $Y=0.054
r11 10 15 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.123 $X2=0.297 $Y2=0.135
r12 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r14 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AOI221XP5_ASAP7_75T_L%Y 1 4 6 7 10 11 12 15 19 21 27 30 33 36 42 45
+ 46 VSS
c25 47 VSS 1.45514e-19 $X=0.099 $Y=0.198
c26 46 VSS 8.46035e-21 $X=0.09 $Y=0.198
c27 45 VSS 3.46932e-19 $X=0.072 $Y=0.198
c28 44 VSS 2.30435e-19 $X=0.04 $Y=0.198
c29 42 VSS 3.3737e-19 $X=0.108 $Y=0.198
c30 40 VSS 0.0019286f $X=0.036 $Y=0.198
c31 38 VSS 9.42062e-19 $X=0.2085 $Y=0.036
c32 37 VSS 2.39163e-19 $X=0.201 $Y=0.036
c33 36 VSS 0.00146362f $X=0.198 $Y=0.036
c34 35 VSS 3.78291e-19 $X=0.18 $Y=0.036
c35 34 VSS 0.00558992f $X=0.176 $Y=0.036
c36 33 VSS 0.00142296f $X=0.144 $Y=0.036
c37 32 VSS 3.47945e-19 $X=0.126 $Y=0.036
c38 31 VSS 0.00315399f $X=0.123 $Y=0.036
c39 30 VSS 0.00146362f $X=0.09 $Y=0.036
c40 29 VSS 0.00368249f $X=0.072 $Y=0.036
c41 27 VSS 0.00283822f $X=0.216 $Y=0.036
c42 22 VSS 0.00336615f $X=0.036 $Y=0.036
c43 21 VSS 0.00423691f $X=0.027 $Y=0.164
c44 20 VSS 0.00112176f $X=0.027 $Y=0.07
c45 19 VSS 0.00112176f $X=0.025 $Y=0.172
c46 15 VSS 0.00233317f $X=0.108 $Y=0.2025
c47 11 VSS 5.68239e-19 $X=0.125 $Y=0.2025
c48 10 VSS 0.00606778f $X=0.216 $Y=0.054
c49 6 VSS 5.5175e-19 $X=0.233 $Y=0.054
c50 4 VSS 0.00319205f $X=0.056 $Y=0.054
c51 1 VSS 2.6657e-19 $X=0.071 $Y=0.054
r52 46 47 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.198 $X2=0.099 $Y2=0.198
r53 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.198 $X2=0.09 $Y2=0.198
r54 44 45 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.198 $X2=0.072 $Y2=0.198
r55 42 47 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.198 $X2=0.099 $Y2=0.198
r56 40 44 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.198 $X2=0.04 $Y2=0.198
r57 37 38 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.201
+ $Y=0.036 $X2=0.2085 $Y2=0.036
r58 36 37 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.201 $Y2=0.036
r59 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r60 34 35 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.036 $X2=0.18 $Y2=0.036
r61 33 34 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.176 $Y2=0.036
r62 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r63 31 32 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.123
+ $Y=0.036 $X2=0.126 $Y2=0.036
r64 30 31 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.123 $Y2=0.036
r65 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r66 27 38 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.2085 $Y2=0.036
r67 24 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.072 $Y2=0.036
r68 22 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.054 $Y2=0.036
r69 20 21 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.164
r70 19 21 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.172 $X2=0.027 $Y2=0.164
r71 17 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.189 $X2=0.036 $Y2=0.198
r72 17 19 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.027 $Y2=0.172
r73 16 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r74 16 20 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r75 15 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.198 $X2=0.108
+ $Y2=0.198
r76 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r77 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r78 10 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r79 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.054 $X2=0.216 $Y2=0.054
r80 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.054 $X2=0.216 $Y2=0.054
r81 4 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r82 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.054 $X2=0.056 $Y2=0.054
.ends


* END of "./AOI221xp5_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI221xp5_ASAP7_75t_L  VSS VDD B1 B2 C A1 A2 Y
* 
* Y	Y
* A2	A2
* A1	A1
* C	C
* B2	B2
* B1	B1
M0 noxref_11 N_B1_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 VSS N_B2_M1_g noxref_11 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_C_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 noxref_12 N_A1_M3_g N_Y_M3_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 VSS N_A2_M4_g noxref_12 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.027
M5 N_Y_M5_d N_B1_M5_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M6 noxref_9 N_B2_M6_g N_Y_M6_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 noxref_10 N_C_M7_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M8 VDD N_A1_M8_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M9 noxref_10 N_A2_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
*
* 
* .include "AOI221xp5_ASAP7_75t_L.pex.sp.AOI221XP5_ASAP7_75T_L.pxi"
* BEGIN of "./AOI221xp5_ASAP7_75t_L.pex.sp.AOI221XP5_ASAP7_75T_L.pxi"
* File: AOI221xp5_ASAP7_75t_L.pex.sp.AOI221XP5_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:11:48 2017
* 
x_PM_AOI221XP5_ASAP7_75T_L%B1 N_B1_M0_g N_B1_c_2_p N_B1_M5_g N_B1_c_3_p B1 VSS
+ PM_AOI221XP5_ASAP7_75T_L%B1
x_PM_AOI221XP5_ASAP7_75T_L%B2 N_B2_M1_g N_B2_c_13_n N_B2_M6_g B2 VSS
+ PM_AOI221XP5_ASAP7_75T_L%B2
x_PM_AOI221XP5_ASAP7_75T_L%C N_C_M2_g N_C_c_25_n N_C_M7_g C VSS
+ PM_AOI221XP5_ASAP7_75T_L%C
x_PM_AOI221XP5_ASAP7_75T_L%A1 N_A1_M3_g N_A1_c_36_n N_A1_M8_g A1 VSS
+ PM_AOI221XP5_ASAP7_75T_L%A1
x_PM_AOI221XP5_ASAP7_75T_L%A2 N_A2_M4_g N_A2_c_46_n N_A2_M9_g A2 VSS
+ PM_AOI221XP5_ASAP7_75T_L%A2
x_PM_AOI221XP5_ASAP7_75T_L%Y N_Y_M0_s N_Y_c_52_n N_Y_M3_s N_Y_M2_d N_Y_c_60_n
+ N_Y_M6_s N_Y_M5_d N_Y_c_68_p Y N_Y_c_53_n N_Y_c_65_n N_Y_c_54_n N_Y_c_58_n
+ N_Y_c_61_n N_Y_c_72_p N_Y_c_66_p N_Y_c_56_n VSS PM_AOI221XP5_ASAP7_75T_L%Y
cc_1 N_B1_M0_g N_B2_M1_g 0.00364065f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_B1_c_2_p N_B2_c_13_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_B1_c_3_p B2 0.00484691f $X=0.081 $Y=0.135 $X2=0.134 $Y2=0.109
cc_4 N_B1_M0_g N_C_M2_g 2.6588e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 N_B1_c_3_p N_Y_c_52_n 3.87865e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_6 N_B1_c_3_p N_Y_c_53_n 0.00441847f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_7 N_B1_M0_g N_Y_c_54_n 2.64276e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_8 N_B1_c_3_p N_Y_c_54_n 0.00124805f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_B1_M0_g N_Y_c_56_n 2.68514e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_10 N_B1_c_3_p N_Y_c_56_n 0.00121543f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 VSS N_B1_M0_g 2.38303e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_12 N_B2_M1_g N_C_M2_g 0.0032267f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_13 N_B2_c_13_n N_C_c_25_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 B2 C 0.00456406f $X=0.134 $Y=0.109 $X2=0.081 $Y2=0.135
cc_15 N_B2_M1_g N_A1_M3_g 2.60137e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_16 N_B2_M1_g N_Y_c_58_n 2.56935e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_17 B2 N_Y_c_58_n 0.00123064f $X=0.134 $Y=0.109 $X2=0 $Y2=0
cc_18 VSS N_B2_M1_g 3.47199e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_19 VSS B2 5.30079e-19 $X=0.134 $Y=0.109 $X2=0 $Y2=0
cc_20 N_C_M2_g N_A1_M3_g 0.00346636f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_21 N_C_c_25_n N_A1_c_36_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 C A1 0.00456406f $X=0.188 $Y=0.123 $X2=0.081 $Y2=0.135
cc_23 N_C_M2_g N_A2_M4_g 2.54394e-19 $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_24 C N_Y_c_60_n 3.31541e-19 $X=0.188 $Y=0.123 $X2=0.081 $Y2=0.135
cc_25 N_C_M2_g N_Y_c_61_n 2.64276e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_26 C N_Y_c_61_n 0.00124805f $X=0.188 $Y=0.123 $X2=0 $Y2=0
cc_27 N_A1_M3_g N_A2_M4_g 0.00310323f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_28 N_A1_c_36_n N_A2_c_46_n 9.33263e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_29 A1 A2 0.00467338f $X=0.24 $Y=0.09 $X2=0.134 $Y2=0.109
cc_30 A1 N_Y_c_60_n 3.87865e-19 $X=0.24 $Y=0.09 $X2=0.134 $Y2=0.109
cc_31 VSS N_A1_M3_g 3.51973e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_32 VSS A1 0.00121543f $X=0.24 $Y=0.09 $X2=0 $Y2=0
cc_33 A2 N_Y_c_60_n 3.94305e-19 $X=0.295 $Y=0.123 $X2=0.188 $Y2=0.123
cc_34 A2 N_Y_c_65_n 4.37254e-19 $X=0.295 $Y=0.123 $X2=0 $Y2=0
cc_35 VSS N_A2_M4_g 3.51973e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_36 VSS A2 0.00122076f $X=0.295 $Y=0.123 $X2=0 $Y2=0
cc_37 VSS N_Y_c_66_p 2.47657e-19 $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.054
cc_38 VSS N_Y_c_52_n 9.98826e-19 $X=0.056 $Y=0.054 $X2=0.081 $Y2=0.135
cc_39 VSS N_Y_c_68_p 0.00371671f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_40 VSS N_Y_c_53_n 3.97918e-19 $X=0.027 $Y=0.164 $X2=0.081 $Y2=0.135
cc_41 VSS N_Y_c_66_p 0.00260156f $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.135
cc_42 VSS N_Y_c_68_p 0.00333582f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_43 VSS N_Y_c_72_p 4.54465e-19 $X=0.108 $Y=0.198 $X2=0.081 $Y2=0.135
cc_44 VSS N_Y_c_68_p 0.00250965f $X=0.108 $Y=0.2025 $X2=0 $Y2=0
cc_45 VSS N_Y_c_66_p 0.00714937f $X=0.072 $Y=0.198 $X2=0 $Y2=0
cc_46 VSS N_Y_c_60_n 9.98826e-19 $X=0.216 $Y=0.054 $X2=0.081 $Y2=0.135
cc_47 VSS N_Y_c_72_p 2.95791e-19 $X=0.108 $Y=0.198 $X2=0 $Y2=0

* END of "./AOI221xp5_ASAP7_75t_L.pex.sp.AOI221XP5_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI222xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:12:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI222xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI222xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI222xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:12:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI222XP33_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c11 10 VSS 6.95749e-19 $X=0.081 $Y=0.135
c12 5 VSS 0.00170784f $X=0.081 $Y=0.135
c13 2 VSS 0.066866f $X=0.081 $Y=0.054
r14 10 14 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.147
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI222XP33_ASAP7_75T_L%A2 2 5 7 10 VSS
c11 10 VSS 0.00105185f $X=0.135 $Y=0.106
c12 5 VSS 0.00113686f $X=0.135 $Y=0.135
c13 2 VSS 0.0624109f $X=0.135 $Y=0.054
r14 10 13 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.106 $X2=0.135 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI222XP33_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c11 10 VSS 0.00105185f $X=0.189 $Y=0.135
c12 5 VSS 0.00113407f $X=0.189 $Y=0.135
c13 2 VSS 0.0624109f $X=0.189 $Y=0.054
r14 10 14 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.151
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI222XP33_ASAP7_75T_L%B1 2 5 7 10 VSS
c11 10 VSS 0.00104792f $X=0.243 $Y=0.098
c12 5 VSS 0.00220625f $X=0.243 $Y=0.135
c13 2 VSS 0.0662287f $X=0.243 $Y=0.054
r14 10 13 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.098 $X2=0.243 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI222XP33_ASAP7_75T_L%C1 2 5 7 10 13 VSS
c11 13 VSS 0.00159102f $X=0.405 $Y=0.135
c12 10 VSS 0.00148639f $X=0.405 $Y=0.094
c13 5 VSS 0.00236647f $X=0.405 $Y=0.135
c14 2 VSS 0.0641039f $X=0.405 $Y=0.054
r15 10 13 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.094 $X2=0.405 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.054 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AOI222XP33_ASAP7_75T_L%C2 2 5 7 10 16 VSS
c8 10 VSS 0.00699786f $X=0.459 $Y=0.135
c9 5 VSS 0.00237052f $X=0.459 $Y=0.135
c10 2 VSS 0.0632655f $X=0.459 $Y=0.054
r11 10 16 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.147
r12 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r14 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.054 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AOI222XP33_ASAP7_75T_L%Y 1 4 6 9 11 14 16 17 20 24 26 37 40 42 44 45
+ 47 49 50 55 58 59 VSS
c32 60 VSS 1.45514e-19 $X=0.099 $Y=0.198
c33 59 VSS 8.46035e-21 $X=0.09 $Y=0.198
c34 58 VSS 3.46932e-19 $X=0.072 $Y=0.198
c35 57 VSS 2.30435e-19 $X=0.04 $Y=0.198
c36 55 VSS 3.25827e-19 $X=0.108 $Y=0.198
c37 53 VSS 0.00192809f $X=0.036 $Y=0.198
c38 50 VSS 9.85989e-19 $X=0.369 $Y=0.036
c39 49 VSS 0.0127368f $X=0.36 $Y=0.036
c40 47 VSS 0.00373091f $X=0.378 $Y=0.036
c41 45 VSS 0.00146362f $X=0.252 $Y=0.036
c42 44 VSS 0.00321019f $X=0.234 $Y=0.036
c43 43 VSS 4.57265e-19 $X=0.202 $Y=0.036
c44 42 VSS 0.00142296f $X=0.198 $Y=0.036
c45 41 VSS 0.00626341f $X=0.18 $Y=0.036
c46 40 VSS 0.00142296f $X=0.144 $Y=0.036
c47 39 VSS 4.57265e-19 $X=0.126 $Y=0.036
c48 38 VSS 0.00305683f $X=0.122 $Y=0.036
c49 37 VSS 0.00146362f $X=0.09 $Y=0.036
c50 36 VSS 0.0036669f $X=0.072 $Y=0.036
c51 29 VSS 0.00339961f $X=0.036 $Y=0.036
c52 28 VSS 5.10117e-19 $X=0.027 $Y=0.1765
c53 26 VSS 0.00171868f $X=0.027 $Y=0.1085
c54 25 VSS 0.00112176f $X=0.027 $Y=0.07
c55 24 VSS 0.00249834f $X=0.02 $Y=0.147
c56 22 VSS 6.07272e-19 $X=0.027 $Y=0.189
c57 20 VSS 0.0023085f $X=0.108 $Y=0.2025
c58 16 VSS 5.76042e-19 $X=0.125 $Y=0.2025
c59 14 VSS 0.0041606f $X=0.38 $Y=0.054
c60 11 VSS 2.6657e-19 $X=0.395 $Y=0.054
c61 9 VSS 0.00352765f $X=0.268 $Y=0.054
c62 4 VSS 0.00319205f $X=0.056 $Y=0.054
c63 1 VSS 2.6657e-19 $X=0.071 $Y=0.054
r64 59 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.198 $X2=0.099 $Y2=0.198
r65 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.198 $X2=0.09 $Y2=0.198
r66 57 58 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.198 $X2=0.072 $Y2=0.198
r67 55 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.198 $X2=0.099 $Y2=0.198
r68 53 57 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.198 $X2=0.04 $Y2=0.198
r69 49 50 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.369 $Y2=0.036
r70 47 50 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.369 $Y2=0.036
r71 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r72 43 44 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.036 $X2=0.234 $Y2=0.036
r73 42 43 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.202 $Y2=0.036
r74 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r75 40 41 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.18 $Y2=0.036
r76 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r77 38 39 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.122
+ $Y=0.036 $X2=0.126 $Y2=0.036
r78 37 38 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.122 $Y2=0.036
r79 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r80 34 49 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.36 $Y2=0.036
r81 34 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.252 $Y2=0.036
r82 31 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.072 $Y2=0.036
r83 29 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.054 $Y2=0.036
r84 27 28 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.164 $X2=0.027 $Y2=0.1765
r85 25 26 2.6142 $w=1.8e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.1085
r86 24 27 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.147 $X2=0.027 $Y2=0.164
r87 24 26 2.6142 $w=1.8e-08 $l=3.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.147 $X2=0.027 $Y2=0.1085
r88 22 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.189 $X2=0.036 $Y2=0.198
r89 22 28 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.027 $Y2=0.1765
r90 21 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r91 21 25 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r92 20 55 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.198 $X2=0.108
+ $Y2=0.198
r93 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r94 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r95 14 47 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r96 11 14 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.054 $X2=0.38 $Y2=0.054
r97 9 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r98 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.054 $X2=0.268 $Y2=0.054
r99 4 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r100 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
.ends


* END of "./AOI222xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI222xp33_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 C1 C2 Y
* 
* Y	Y
* C2	C2
* C1	C1
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 noxref_12 N_A1_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 VSS N_A2_M1_g noxref_12 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 noxref_13 N_B2_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.027
M3 N_Y_M3_d N_B1_M3_g noxref_13 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 noxref_14 N_C1_M4_g N_Y_M4_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.395
+ $Y=0.027
M5 VSS N_C2_M5_g noxref_14 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.449
+ $Y=0.027
M6 N_Y_M6_d N_A1_M6_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 noxref_10 N_A2_M7_g N_Y_M7_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 noxref_11 N_B2_M8_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 noxref_10 N_B1_M9_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 noxref_11 N_C1_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M11 VDD N_C2_M11_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "AOI222xp33_ASAP7_75t_L.pex.sp.AOI222XP33_ASAP7_75T_L.pxi"
* BEGIN of "./AOI222xp33_ASAP7_75t_L.pex.sp.AOI222XP33_ASAP7_75T_L.pxi"
* File: AOI222xp33_ASAP7_75t_L.pex.sp.AOI222XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:12:10 2017
* 
x_PM_AOI222XP33_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M6_g N_A1_c_3_p A1 VSS
+ PM_AOI222XP33_ASAP7_75T_L%A1
x_PM_AOI222XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_13_n N_A2_M7_g A2 VSS
+ PM_AOI222XP33_ASAP7_75T_L%A2
x_PM_AOI222XP33_ASAP7_75T_L%B2 N_B2_M2_g N_B2_c_25_n N_B2_M8_g N_B2_c_26_n B2
+ VSS PM_AOI222XP33_ASAP7_75T_L%B2
x_PM_AOI222XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_36_n N_B1_M9_g B1 VSS
+ PM_AOI222XP33_ASAP7_75T_L%B1
x_PM_AOI222XP33_ASAP7_75T_L%C1 N_C1_M4_g N_C1_c_47_p N_C1_M10_g C1 N_C1_c_53_p
+ VSS PM_AOI222XP33_ASAP7_75T_L%C1
x_PM_AOI222XP33_ASAP7_75T_L%C2 N_C2_M5_g N_C2_c_57_n N_C2_M11_g N_C2_c_58_n C2
+ VSS PM_AOI222XP33_ASAP7_75T_L%C2
x_PM_AOI222XP33_ASAP7_75T_L%Y N_Y_M0_s N_Y_c_64_n N_Y_M3_d N_Y_c_74_n N_Y_M4_s
+ N_Y_c_77_n N_Y_M7_s N_Y_M6_d N_Y_c_84_p Y N_Y_c_65_n N_Y_c_66_n N_Y_c_70_n
+ N_Y_c_72_n N_Y_c_92_p N_Y_c_75_n N_Y_c_78_n N_Y_c_94_p N_Y_c_95_p N_Y_c_88_p
+ N_Y_c_82_p N_Y_c_68_n VSS PM_AOI222XP33_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00372052f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A1_c_2_p N_A2_c_13_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p A2 0.00484691f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.106
cc_4 N_A1_M0_g N_B2_M2_g 2.74891e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 N_A1_c_3_p N_Y_c_64_n 3.87865e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_6 N_A1_c_3_p N_Y_c_65_n 0.00440851f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_7 N_A1_M0_g N_Y_c_66_n 2.64276e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_8 N_A1_c_3_p N_Y_c_66_n 0.00124805f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_A1_M0_g N_Y_c_68_n 2.68514e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_10 N_A1_c_3_p N_Y_c_68_n 0.00121543f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 VSS N_A1_M0_g 2.38303e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_12 N_A2_M1_g N_B2_M2_g 0.00335739f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_13 N_A2_c_13_n N_B2_c_25_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 A2 N_B2_c_26_n 0.00456406f $X=0.135 $Y=0.106 $X2=0.081 $Y2=0.135
cc_15 N_A2_M1_g N_B1_M3_g 2.74891e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_16 N_A2_M1_g N_Y_c_70_n 2.56935e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_17 A2 N_Y_c_70_n 0.00123064f $X=0.135 $Y=0.106 $X2=0 $Y2=0
cc_18 VSS N_A2_M1_g 3.47199e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_19 VSS A2 5.30079e-19 $X=0.135 $Y=0.106 $X2=0 $Y2=0
cc_20 N_B2_M2_g N_B1_M3_g 0.00372052f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_21 N_B2_c_25_n N_B1_c_36_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 N_B2_c_26_n B1 0.00484691f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 N_B2_M2_g N_Y_c_72_n 2.56935e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_24 N_B2_c_26_n N_Y_c_72_n 0.00123064f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_25 VSS N_B2_M2_g 3.57119e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_26 VSS N_B2_c_26_n 5.37372e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_27 B1 C1 7.84009e-19 $X=0.243 $Y=0.098 $X2=0.135 $Y2=0.106
cc_28 B1 N_Y_c_74_n 4.42987e-19 $X=0.243 $Y=0.098 $X2=0.135 $Y2=0.106
cc_29 N_B1_M3_g N_Y_c_75_n 2.64276e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_30 B1 N_Y_c_75_n 0.00124805f $X=0.243 $Y=0.098 $X2=0 $Y2=0
cc_31 VSS N_B1_M3_g 2.08515e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_32 VSS N_B1_M3_g 2.76185e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_33 VSS B1 0.0012322f $X=0.243 $Y=0.098 $X2=0 $Y2=0
cc_34 N_C1_M4_g N_C2_M5_g 0.00347357f $X=0.405 $Y=0.054 $X2=0.243 $Y2=0.054
cc_35 N_C1_c_47_p N_C2_c_57_n 9.79748e-19 $X=0.405 $Y=0.135 $X2=0.243 $Y2=0.135
cc_36 C1 N_C2_c_58_n 0.00565736f $X=0.405 $Y=0.094 $X2=0.243 $Y2=0.098
cc_37 C1 N_Y_c_77_n 4.42987e-19 $X=0.405 $Y=0.094 $X2=0.243 $Y2=0.135
cc_38 N_C1_M4_g N_Y_c_78_n 2.7362e-19 $X=0.405 $Y=0.054 $X2=0 $Y2=0
cc_39 C1 N_Y_c_78_n 2.0892e-19 $X=0.405 $Y=0.094 $X2=0 $Y2=0
cc_40 VSS C1 0.0011319f $X=0.405 $Y=0.094 $X2=0.243 $Y2=0.098
cc_41 VSS N_C1_c_53_p 4.64783e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_42 VSS N_C1_M4_g 2.56935e-19 $X=0.405 $Y=0.054 $X2=0 $Y2=0
cc_43 VSS N_C1_c_53_p 0.00125352f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_44 N_C2_c_58_n N_Y_c_77_n 3.94305e-19 $X=0.459 $Y=0.135 $X2=0.405 $Y2=0.135
cc_45 N_C2_c_58_n N_Y_c_78_n 4.94602e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_46 VSS N_C2_c_58_n 0.00114532f $X=0.459 $Y=0.135 $X2=0.405 $Y2=0.094
cc_47 VSS N_C2_M5_g 2.7596e-19 $X=0.459 $Y=0.054 $X2=0 $Y2=0
cc_48 VSS N_C2_c_58_n 0.00125674f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_49 VSS N_Y_c_82_p 2.47657e-19 $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.054
cc_50 VSS N_Y_c_64_n 9.98826e-19 $X=0.056 $Y=0.054 $X2=0.081 $Y2=0.135
cc_51 VSS N_Y_c_84_p 0.00371671f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_52 VSS Y 4.01247e-19 $X=0.02 $Y=0.147 $X2=0.081 $Y2=0.135
cc_53 VSS N_Y_c_82_p 0.00260156f $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.135
cc_54 VSS N_Y_c_84_p 0.0033367f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_55 VSS N_Y_c_88_p 4.49388e-19 $X=0.108 $Y=0.198 $X2=0.081 $Y2=0.135
cc_56 VSS N_Y_c_74_n 9.98826e-19 $X=0.268 $Y=0.054 $X2=0.081 $Y2=0.147
cc_57 VSS N_Y_c_84_p 0.00250965f $X=0.108 $Y=0.2025 $X2=0 $Y2=0
cc_58 VSS N_Y_c_82_p 0.00705695f $X=0.072 $Y=0.198 $X2=0 $Y2=0
cc_59 VSS N_Y_c_92_p 8.06874e-19 $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_60 VSS N_Y_c_88_p 2.89103e-19 $X=0.108 $Y=0.198 $X2=0 $Y2=0
cc_61 VSS N_Y_c_94_p 8.06874e-19 $X=0.36 $Y=0.036 $X2=0 $Y2=0
cc_62 VSS N_Y_c_95_p 2.13649e-19 $X=0.369 $Y=0.036 $X2=0 $Y2=0

* END of "./AOI222xp33_ASAP7_75t_L.pex.sp.AOI222XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI22x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:12:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI22x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI22x1_ASAP7_75t_L.pex.sp.pex"
* File: AOI22x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:12:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI22X1_ASAP7_75T_L%B2 2 5 7 10 13 15 20 22 24 26 27 28 29 30 34 36
+ 37 VSS
c34 37 VSS 6.90135e-20 $X=0.243 $Y=0.117
c35 36 VSS 3.51388e-19 $X=0.243 $Y=0.099
c36 34 VSS 1.78839e-19 $X=0.243 $Y=0.135
c37 31 VSS 5.67196e-19 $X=0.216 $Y=0.072
c38 30 VSS 0.00158425f $X=0.198 $Y=0.072
c39 29 VSS 0.00207482f $X=0.161 $Y=0.072
c40 28 VSS 1.5733e-19 $X=0.109 $Y=0.072
c41 27 VSS 4.68273e-20 $X=0.09 $Y=0.072
c42 26 VSS 1.94766e-19 $X=0.234 $Y=0.072
c43 24 VSS 0.00169746f $X=0.081 $Y=0.135
c44 22 VSS 3.54309e-19 $X=0.081 $Y=0.117
c45 21 VSS 3.51388e-19 $X=0.081 $Y=0.099
c46 20 VSS 0.00166207f $X=0.081 $Y=0.118
c47 13 VSS 9.94291e-19 $X=0.243 $Y=0.135
c48 10 VSS 0.0597239f $X=0.243 $Y=0.0675
c49 5 VSS 0.00251885f $X=0.081 $Y=0.135
c50 2 VSS 0.0641711f $X=0.081 $Y=0.0675
r51 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.099 $X2=0.243 $Y2=0.117
r52 34 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.117
r53 32 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.099
r54 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.072 $X2=0.216 $Y2=0.072
r55 29 30 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.161
+ $Y=0.072 $X2=0.198 $Y2=0.072
r56 28 29 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.072 $X2=0.161 $Y2=0.072
r57 27 28 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.109 $Y2=0.072
r58 26 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.072 $X2=0.243 $Y2=0.081
r59 26 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.216 $Y2=0.072
r60 21 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.099 $X2=0.081 $Y2=0.117
r61 20 24 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.118 $X2=0.081 $Y2=0.135
r62 20 22 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.118 $X2=0.081 $Y2=0.117
r63 17 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.081 $X2=0.09 $Y2=0.072
r64 17 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.081 $X2=0.081 $Y2=0.099
r65 13 34 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r66 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r67 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r68 5 24 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r69 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r70 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI22X1_ASAP7_75T_L%B1 2 7 10 13 15 20 25 VSS
c25 25 VSS 0.00123481f $X=0.183 $Y=0.108
c26 20 VSS 0.00303344f $X=0.189 $Y=0.135
c27 13 VSS 0.00532127f $X=0.189 $Y=0.135
c28 10 VSS 0.0613446f $X=0.189 $Y=0.0675
c29 2 VSS 0.0619872f $X=0.135 $Y=0.0675
r30 17 25 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.11225 $X2=0.183 $Y2=0.11225
r31 17 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.117 $X2=0.189 $Y2=0.135
r32 13 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r33 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r34 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r35 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r36 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r37 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI22X1_ASAP7_75T_L%A2 2 5 7 10 13 15 19 21 24 26 27 29 30 31 35 38
+ VSS
c39 38 VSS 2.00449e-19 $X=0.459 $Y=0.117
c40 37 VSS 3.51388e-19 $X=0.459 $Y=0.099
c41 35 VSS 7.84621e-19 $X=0.459 $Y=0.135
c42 31 VSS 0.00192557f $X=0.431 $Y=0.072
c43 30 VSS 0.00158425f $X=0.379 $Y=0.072
c44 29 VSS 3.27558e-19 $X=0.342 $Y=0.072
c45 28 VSS 2.02211e-20 $X=0.309 $Y=0.072
c46 27 VSS 4.67409e-20 $X=0.306 $Y=0.072
c47 26 VSS 1.49134e-19 $X=0.45 $Y=0.072
c48 24 VSS 6.90135e-20 $X=0.297 $Y=0.117
c49 21 VSS 1.26672e-19 $X=0.297 $Y=0.135
c50 19 VSS 3.51388e-19 $X=0.296 $Y=0.087
c51 13 VSS 0.00128572f $X=0.459 $Y=0.135
c52 10 VSS 0.065901f $X=0.459 $Y=0.0675
c53 5 VSS 0.00150858f $X=0.297 $Y=0.135
c54 2 VSS 0.0607585f $X=0.297 $Y=0.0675
r55 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.099 $X2=0.459 $Y2=0.117
r56 35 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.117
r57 32 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.099
r58 30 31 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.072 $X2=0.431 $Y2=0.072
r59 29 30 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.072 $X2=0.379 $Y2=0.072
r60 28 29 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.309
+ $Y=0.072 $X2=0.342 $Y2=0.072
r61 27 28 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.072 $X2=0.309 $Y2=0.072
r62 26 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.072 $X2=0.459 $Y2=0.081
r63 26 31 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.072 $X2=0.431 $Y2=0.072
r64 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.099 $X2=0.297 $Y2=0.117
r65 21 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.117
r66 19 23 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.087 $X2=0.297 $Y2=0.099
r67 17 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.297 $Y=0.081 $X2=0.306 $Y2=0.072
r68 17 19 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.081 $X2=0.297 $Y2=0.087
r69 13 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r70 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r71 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r72 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r73 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r74 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AOI22X1_ASAP7_75T_L%A1 2 7 10 13 15 18 20 28 VSS
c28 20 VSS 0.00143833f $X=0.351 $Y=0.135
c29 18 VSS 4.67848e-19 $X=0.351 $Y=0.153
c30 13 VSS 0.00513876f $X=0.405 $Y=0.135
c31 10 VSS 0.0637114f $X=0.405 $Y=0.0675
c32 2 VSS 0.0625799f $X=0.351 $Y=0.0675
r33 22 23 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.152 $X2=0.351 $Y2=0.1525
r34 20 22 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.152
r35 18 28 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1575 $X2=0.359 $Y2=0.1575
r36 18 23 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.153 $X2=0.351 $Y2=0.1525
r37 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r38 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
r39 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r40 5 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r41 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r42 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AOI22X1_ASAP7_75T_L%Y 1 6 7 11 16 17 20 21 22 25 29 35 37 40 42 51 52
+ 53 55 56 60 62 VSS
c46 64 VSS 4.55454e-19 $X=0.513 $Y=0.18
c47 62 VSS 9.85346e-19 $X=0.513 $Y=0.0885
c48 61 VSS 8.85605e-19 $X=0.513 $Y=0.063
c49 60 VSS 0.00358506f $X=0.513 $Y=0.114
c50 58 VSS 4.30151e-19 $X=0.513 $Y=0.189
c51 56 VSS 3.46932e-19 $X=0.5 $Y=0.198
c52 55 VSS 8.46035e-21 $X=0.468 $Y=0.198
c53 53 VSS 3.69675e-19 $X=0.431 $Y=0.198
c54 52 VSS 5.76352e-20 $X=0.379 $Y=0.198
c55 51 VSS 5.76656e-19 $X=0.342 $Y=0.198
c56 43 VSS 0.0021974f $X=0.504 $Y=0.198
c57 42 VSS 0.0176071f $X=0.468 $Y=0.036
c58 41 VSS 0.00359728f $X=0.288 $Y=0.036
c59 40 VSS 0.00354992f $X=0.486 $Y=0.036
c60 37 VSS 0.0176042f $X=0.252 $Y=0.036
c61 36 VSS 0.00257895f $X=0.072 $Y=0.036
c62 35 VSS 0.00480088f $X=0.27 $Y=0.036
c63 29 VSS 0.00359039f $X=0.054 $Y=0.036
c64 28 VSS 0.00223184f $X=0.054 $Y=0.036
c65 26 VSS 0.00709337f $X=0.504 $Y=0.036
c66 25 VSS 0.00215645f $X=0.432 $Y=0.2025
c67 21 VSS 7.35996e-19 $X=0.449 $Y=0.2025
c68 20 VSS 0.0025205f $X=0.324 $Y=0.2025
c69 16 VSS 6.53507e-19 $X=0.341 $Y=0.2025
c70 14 VSS 2.69461e-19 $X=0.484 $Y=0.0675
c71 6 VSS 5.38922e-19 $X=0.287 $Y=0.0675
c72 1 VSS 2.69461e-19 $X=0.071 $Y=0.0675
r73 63 64 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.171 $X2=0.513 $Y2=0.18
r74 61 62 1.73148 $w=1.8e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.063 $X2=0.513 $Y2=0.0885
r75 60 63 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.114 $X2=0.513 $Y2=0.171
r76 60 62 1.73148 $w=1.8e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.114 $X2=0.513 $Y2=0.0885
r77 58 64 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.513 $Y2=0.18
r78 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.063
r79 55 56 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.198 $X2=0.5 $Y2=0.198
r80 53 54 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.198 $X2=0.4315 $Y2=0.198
r81 52 53 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.198 $X2=0.431 $Y2=0.198
r82 51 52 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.379 $Y2=0.198
r83 49 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.468 $Y2=0.198
r84 49 54 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.4315 $Y2=0.198
r85 45 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.342 $Y2=0.198
r86 43 58 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.198 $X2=0.513 $Y2=0.189
r87 43 56 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.198 $X2=0.5 $Y2=0.198
r88 41 42 12.2222 $w=1.8e-08 $l=1.8e-07 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.468 $Y2=0.036
r89 39 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.468 $Y2=0.036
r90 39 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036 $X2=0.486
+ $Y2=0.036
r91 36 37 12.2222 $w=1.8e-08 $l=1.8e-07 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.252 $Y2=0.036
r92 34 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.288 $Y2=0.036
r93 34 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.252 $Y2=0.036
r94 34 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r95 28 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.072 $Y2=0.036
r96 28 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r97 26 57 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.036 $X2=0.513 $Y2=0.045
r98 26 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.486 $Y2=0.036
r99 25 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r100 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r101 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r102 20 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198
+ $X2=0.324 $Y2=0.198
r103 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r104 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r105 14 40 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.486 $Y=0.0675 $X2=0.486 $Y2=0.036
r106 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.484 $Y2=0.0675
r107 10 35 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r108 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r109 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r110 4 29 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r111 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./AOI22x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI22x1_ASAP7_75t_L  VSS VDD B2 B1 A2 A1 Y
* 
* Y	Y
* A1	A1
* A2	A2
* B1	B1
* B2	B2
M0 N_Y_M0_d N_B2_M0_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_9 N_B1_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_10 N_B1_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_Y_M3_d N_B2_M3_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_A2_M4_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_11 N_A1_M5_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_12 N_A1_M6_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_Y_M7_d N_A2_M7_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 VDD N_B2_M8_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M9 noxref_7 N_B1_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M10 noxref_7 N_B1_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M11 VDD N_B2_M11_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M12 N_Y_M12_d N_A2_M12_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M13 noxref_7 N_A1_M13_g N_Y_M13_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M14 noxref_7 N_A1_M14_g N_Y_M14_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M15 N_Y_M15_d N_A2_M15_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "AOI22x1_ASAP7_75t_L.pex.sp.AOI22X1_ASAP7_75T_L.pxi"
* BEGIN of "./AOI22x1_ASAP7_75t_L.pex.sp.AOI22X1_ASAP7_75T_L.pxi"
* File: AOI22x1_ASAP7_75t_L.pex.sp.AOI22X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:12:33 2017
* 
x_PM_AOI22X1_ASAP7_75T_L%B2 N_B2_M0_g N_B2_c_7_p N_B2_M8_g N_B2_M3_g N_B2_c_8_p
+ N_B2_M11_g B2 N_B2_c_13_p N_B2_c_11_p N_B2_c_21_p N_B2_c_30_p N_B2_c_26_p
+ N_B2_c_3_p N_B2_c_6_p N_B2_c_12_p N_B2_c_18_p N_B2_c_15_p VSS
+ PM_AOI22X1_ASAP7_75T_L%B2
x_PM_AOI22X1_ASAP7_75T_L%B1 N_B1_M1_g N_B1_M9_g N_B1_M2_g N_B1_c_41_n N_B1_M10_g
+ N_B1_c_44_n B1 VSS PM_AOI22X1_ASAP7_75T_L%B1
x_PM_AOI22X1_ASAP7_75T_L%A2 N_A2_M4_g N_A2_c_61_n N_A2_M12_g N_A2_M7_g
+ N_A2_c_74_p N_A2_M15_g A2 N_A2_c_63_n N_A2_c_64_n N_A2_c_88_p N_A2_c_65_n
+ N_A2_c_92_p N_A2_c_69_p N_A2_c_72_p N_A2_c_76_p N_A2_c_81_p VSS
+ PM_AOI22X1_ASAP7_75T_L%A2
x_PM_AOI22X1_ASAP7_75T_L%A1 N_A1_M5_g N_A1_M13_g N_A1_M6_g N_A1_c_106_n
+ N_A1_M14_g N_A1_c_109_n N_A1_c_110_n A1 VSS PM_AOI22X1_ASAP7_75T_L%A1
x_PM_AOI22X1_ASAP7_75T_L%Y N_Y_M0_d N_Y_M4_d N_Y_M3_d N_Y_M7_d N_Y_M13_s
+ N_Y_M12_d N_Y_c_146_n N_Y_M15_d N_Y_M14_s N_Y_c_134_n N_Y_c_127_n N_Y_c_128_n
+ N_Y_c_129_n N_Y_c_136_n N_Y_c_137_n N_Y_c_140_n N_Y_c_149_n N_Y_c_141_n
+ N_Y_c_142_n N_Y_c_167_n Y N_Y_c_145_n VSS PM_AOI22X1_ASAP7_75T_L%Y
cc_1 N_B2_M0_g N_B1_M1_g 0.00315405f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_B2_M3_g N_B1_M1_g 2.25374e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_3 N_B2_c_3_p N_B1_M1_g 3.97719e-19 $X=0.161 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_4 N_B2_M0_g N_B1_M2_g 2.25374e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_5 N_B2_M3_g N_B1_M2_g 0.00315405f $X=0.243 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_6 N_B2_c_6_p N_B1_M2_g 2.52885e-19 $X=0.198 $Y=0.072 $X2=0.189 $Y2=0.0675
cc_7 N_B2_c_7_p N_B1_c_41_n 0.00130109f $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_8 N_B2_c_8_p N_B1_c_41_n 9.59209e-19 $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.135
cc_9 N_B2_c_3_p N_B1_c_41_n 7.25985e-19 $X=0.161 $Y=0.072 $X2=0.189 $Y2=0.135
cc_10 B2 N_B1_c_44_n 8.58272e-19 $X=0.081 $Y=0.118 $X2=0.189 $Y2=0.135
cc_11 N_B2_c_11_p N_B1_c_44_n 3.88222e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_12 N_B2_c_12_p N_B1_c_44_n 0.00124457f $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.135
cc_13 N_B2_c_13_p B1 4.40275e-19 $X=0.081 $Y=0.117 $X2=0.183 $Y2=0.108
cc_14 N_B2_c_6_p B1 0.00373189f $X=0.198 $Y=0.072 $X2=0.183 $Y2=0.108
cc_15 N_B2_c_15_p B1 0.00124457f $X=0.243 $Y=0.117 $X2=0.183 $Y2=0.108
cc_16 N_B2_M3_g N_A2_M4_g 0.00353901f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_17 N_B2_c_8_p N_A2_c_61_n 8.87978e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_18 N_B2_c_18_p A2 9.57742e-19 $X=0.243 $Y=0.099 $X2=0.189 $Y2=0.135
cc_19 N_B2_c_12_p N_A2_c_63_n 9.57742e-19 $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.135
cc_20 N_B2_c_15_p N_A2_c_64_n 9.57742e-19 $X=0.243 $Y=0.117 $X2=0.183
+ $Y2=0.11225
cc_21 N_B2_c_21_p N_A2_c_65_n 9.57742e-19 $X=0.234 $Y=0.072 $X2=0 $Y2=0
cc_22 N_B2_M3_g N_A1_M5_g 2.949e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_23 VSS B2 8.25153e-19 $X=0.081 $Y=0.118 $X2=0.135 $Y2=0.135
cc_24 VSS N_B2_M0_g 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_25 VSS N_B2_c_11_p 0.00377207f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_26 VSS N_B2_c_26_p 2.48779e-19 $X=0.109 $Y=0.072 $X2=0 $Y2=0
cc_27 VSS N_B2_c_3_p 2.48779e-19 $X=0.161 $Y=0.072 $X2=0 $Y2=0
cc_28 VSS N_B2_M3_g 3.62717e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_29 VSS N_B2_c_12_p 4.46831e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_30 N_B2_c_30_p N_Y_c_127_n 0.0010499f $X=0.09 $Y=0.072 $X2=0.135 $Y2=0.135
cc_31 N_B2_c_21_p N_Y_c_128_n 0.00159517f $X=0.234 $Y=0.072 $X2=0 $Y2=0
cc_32 N_B2_M0_g N_Y_c_129_n 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_33 N_B2_M3_g N_Y_c_129_n 2.38303e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_34 N_B2_c_30_p N_Y_c_129_n 0.016433f $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_35 N_B1_M2_g N_A2_M4_g 2.60137e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_36 VSS N_B1_c_41_n 3.80455e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_37 VSS N_B1_c_41_n 8.00061e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_38 VSS N_B1_c_44_n 0.00205998f $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_39 VSS N_B1_M1_g 4.62717e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_40 VSS N_B1_c_41_n 3.50613e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.135
cc_41 VSS N_B1_M2_g 2.34993e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_42 VSS N_B1_c_44_n 0.00372108f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_43 N_B1_M1_g N_Y_c_129_n 2.64781e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.117
cc_44 N_B1_M2_g N_Y_c_129_n 2.38303e-19 $X=0.189 $Y=0.0675 $X2=0.243 $Y2=0.117
cc_45 N_A2_M4_g N_A1_M5_g 0.00358983f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_46 N_A2_M7_g N_A1_M5_g 2.6588e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_47 N_A2_c_69_p N_A1_M5_g 2.52885e-19 $X=0.379 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_48 N_A2_M4_g N_A1_M6_g 2.6588e-19 $X=0.297 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_49 N_A2_M7_g N_A1_M6_g 0.00364065f $X=0.459 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_50 N_A2_c_72_p N_A1_M6_g 3.99641e-19 $X=0.431 $Y=0.072 $X2=0.243 $Y2=0.0675
cc_51 N_A2_c_61_n N_A1_c_106_n 9.81317e-19 $X=0.297 $Y=0.135 $X2=0.243 $Y2=0.135
cc_52 N_A2_c_74_p N_A1_c_106_n 0.00129593f $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.135
cc_53 N_A2_c_72_p N_A1_c_106_n 6.92083e-19 $X=0.431 $Y=0.072 $X2=0.243 $Y2=0.135
cc_54 N_A2_c_76_p N_A1_c_109_n 5.64422e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_55 N_A2_c_63_n N_A1_c_110_n 0.00119724f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.118
cc_56 N_A2_c_64_n N_A1_c_110_n 0.00119724f $X=0.297 $Y=0.117 $X2=0.081 $Y2=0.118
cc_57 N_A2_c_69_p N_A1_c_110_n 0.00371882f $X=0.379 $Y=0.072 $X2=0.081 $Y2=0.118
cc_58 N_A2_c_76_p N_A1_c_110_n 4.71615e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.118
cc_59 N_A2_c_81_p N_A1_c_110_n 4.25941e-19 $X=0.459 $Y=0.117 $X2=0.081 $Y2=0.118
cc_60 VSS N_A2_c_76_p 2.73699e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.135
cc_61 VSS N_A2_M4_g 3.75866e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_62 VSS N_A2_c_63_n 4.38244e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_63 VSS N_A2_M7_g 2.38303e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_A2_c_76_p N_Y_c_134_n 0.0313705f $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.135
cc_65 N_A2_c_65_n N_Y_c_128_n 0.00159517f $X=0.306 $Y=0.072 $X2=0.243 $Y2=0.135
cc_66 N_A2_c_88_p N_Y_c_136_n 0.00158881f $X=0.45 $Y=0.072 $X2=0 $Y2=0
cc_67 N_A2_M4_g N_Y_c_137_n 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_68 N_A2_M7_g N_Y_c_137_n 2.38303e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_69 N_A2_c_65_n N_Y_c_137_n 0.0164209f $X=0.306 $Y=0.072 $X2=0 $Y2=0
cc_70 N_A2_c_92_p N_Y_c_140_n 3.65124e-19 $X=0.342 $Y=0.072 $X2=0 $Y2=0
cc_71 N_A2_c_72_p N_Y_c_141_n 3.65124e-19 $X=0.431 $Y=0.072 $X2=0 $Y2=0
cc_72 N_A2_M7_g N_Y_c_142_n 2.52885e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_73 N_A2_c_76_p N_Y_c_142_n 0.00371986f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_74 N_A2_c_81_p Y 0.00218861f $X=0.459 $Y=0.117 $X2=0 $Y2=0
cc_75 N_A2_c_88_p N_Y_c_145_n 0.00218861f $X=0.45 $Y=0.072 $X2=0 $Y2=0
cc_76 VSS N_A2_c_92_p 2.54007e-19 $X=0.342 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_77 VSS N_A1_c_106_n 3.78279e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_78 VSS N_A1_c_106_n 8.00061e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.118
cc_79 VSS N_A1_c_109_n 8.76024e-19 $X=0.351 $Y=0.153 $X2=0.081 $Y2=0.118
cc_80 VSS N_A1_M5_g 2.15135e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_81 VSS N_A1_M6_g 2.64781e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_82 N_A1_c_109_n N_Y_c_146_n 3.21662e-19 $X=0.351 $Y=0.153 $X2=0.081 $Y2=0.118
cc_83 N_A1_M5_g N_Y_c_137_n 2.38303e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_84 N_A1_M6_g N_Y_c_137_n 2.64781e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_85 N_A1_M5_g N_Y_c_149_n 2.56447e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_86 N_A1_c_109_n N_Y_c_149_n 0.00373962f $X=0.351 $Y=0.153 $X2=0 $Y2=0
cc_87 N_A1_M6_g N_Y_c_141_n 3.99641e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_88 N_A1_c_106_n N_Y_c_141_n 5.37025e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_89 VSS N_Y_c_146_n 0.00339475f $X=0.27 $Y=0.2025 $X2=0.081 $Y2=0.118
cc_90 VSS N_Y_c_146_n 0.0036466f $X=0.378 $Y=0.2025 $X2=0.081 $Y2=0.118
cc_91 VSS N_Y_c_146_n 0.00250965f $X=0.3435 $Y=0.234 $X2=0.081 $Y2=0.118
cc_92 VSS N_Y_c_134_n 0.00372512f $X=0.378 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_93 VSS N_Y_c_134_n 0.00384465f $X=0.484 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_94 VSS N_Y_c_134_n 0.00251378f $X=0.486 $Y=0.234 $X2=0.081 $Y2=0.135
cc_95 VSS N_Y_c_127_n 0.00107252f $X=0.056 $Y=0.2025 $X2=0.161 $Y2=0.072
cc_96 VSS N_Y_c_128_n 0.00107252f $X=0.27 $Y=0.2025 $X2=0.243 $Y2=0.135
cc_97 VSS N_Y_c_136_n 0.00138157f $X=0.484 $Y=0.2025 $X2=0 $Y2=0
cc_98 VSS N_Y_c_140_n 5.00406e-19 $X=0.27 $Y=0.2025 $X2=0 $Y2=0
cc_99 VSS N_Y_c_140_n 0.00796074f $X=0.3435 $Y=0.234 $X2=0 $Y2=0
cc_100 VSS N_Y_c_149_n 0.00128262f $X=0.378 $Y=0.2025 $X2=0 $Y2=0
cc_101 VSS N_Y_c_141_n 0.00107804f $X=0.378 $Y=0.2025 $X2=0 $Y2=0
cc_102 VSS N_Y_c_141_n 0.00796074f $X=0.486 $Y=0.234 $X2=0 $Y2=0
cc_103 VSS N_Y_c_167_n 0.00284922f $X=0.484 $Y=0.2025 $X2=0 $Y2=0
cc_104 VSS Y 2.85653e-19 $X=0.484 $Y=0.2025 $X2=0 $Y2=0
cc_105 VSS N_Y_c_129_n 2.27254e-19 $X=0.252 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_106 VSS N_Y_c_129_n 2.21722e-19 $X=0.252 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_107 VSS N_Y_c_137_n 2.27254e-19 $X=0.468 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_108 VSS N_Y_c_137_n 2.27254e-19 $X=0.468 $Y=0.036 $X2=0.081 $Y2=0.0675

* END of "./AOI22x1_ASAP7_75t_L.pex.sp.AOI22X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI22xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:12:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI22xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI22xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI22xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:12:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI22XP33_ASAP7_75T_L%A1 2 5 7 16 19 21 22 27 VSS
c16 27 VSS 0.0126747f $X=0.018 $Y=0.135
c17 22 VSS 7.38238e-19 $X=0.0635 $Y=0.135
c18 21 VSS 8.96246e-19 $X=0.046 $Y=0.135
c19 19 VSS 9.11762e-19 $X=0.081 $Y=0.135
c20 16 VSS 0.00527659f $X=0.018 $Y=0.151
c21 5 VSS 0.00273648f $X=0.081 $Y=0.135
c22 2 VSS 0.0646282f $X=0.081 $Y=0.054
r23 21 22 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r24 19 22 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r25 17 27 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r26 17 21 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.046 $Y2=0.135
r27 13 27 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r28 13 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.151
r29 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r30 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r31 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI22XP33_ASAP7_75T_L%A2 2 5 7 15 21 23 VSS
c18 23 VSS 1.81759e-19 $X=0.135 $Y=0.164
c19 21 VSS 0.00477153f $X=0.135 $Y=0.186
c20 15 VSS 0.00127134f $X=0.135 $Y=0.135
c21 5 VSS 0.00128502f $X=0.135 $Y=0.135
c22 2 VSS 0.0602909f $X=0.135 $Y=0.054
r23 22 23 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.164
r24 21 23 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.186 $X2=0.135 $Y2=0.164
r25 15 22 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r26 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI22XP33_ASAP7_75T_L%B2 2 5 7 10 VSS
c12 10 VSS 6.22747e-19 $X=0.188 $Y=0.115
c13 5 VSS 0.00110682f $X=0.189 $Y=0.135
c14 2 VSS 0.0604449f $X=0.189 $Y=0.054
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI22XP33_ASAP7_75T_L%B1 2 5 7 10 VSS
c10 10 VSS 9.28859e-19 $X=0.245 $Y=0.081
c11 5 VSS 0.00170643f $X=0.243 $Y=0.135
c12 2 VSS 0.0641824f $X=0.243 $Y=0.054
r13 10 13 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.135
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI22XP33_ASAP7_75T_L%Y 1 2 5 6 7 10 16 17 20 27 28 29 34 36 VSS
c19 38 VSS 7.1545e-19 $X=0.297 $Y=0.1765
c20 36 VSS 0.00101238f $X=0.297 $Y=0.092
c21 35 VSS 0.00131846f $X=0.297 $Y=0.07
c22 34 VSS 0.00327462f $X=0.297 $Y=0.114
c23 32 VSS 6.07272e-19 $X=0.297 $Y=0.189
c24 30 VSS 1.42799e-19 $X=0.286 $Y=0.198
c25 29 VSS 5.28464e-19 $X=0.284 $Y=0.198
c26 28 VSS 8.46035e-21 $X=0.252 $Y=0.198
c27 27 VSS 5.02599e-19 $X=0.234 $Y=0.198
c28 22 VSS 0.00199921f $X=0.288 $Y=0.198
c29 21 VSS 0.00332628f $X=0.27 $Y=0.036
c30 20 VSS 0.00142296f $X=0.252 $Y=0.036
c31 19 VSS 0.00311169f $X=0.234 $Y=0.036
c32 18 VSS 4.25461e-19 $X=0.202 $Y=0.036
c33 17 VSS 0.00146362f $X=0.198 $Y=0.036
c34 16 VSS 0.00393804f $X=0.18 $Y=0.036
c35 11 VSS 0.00630045f $X=0.288 $Y=0.036
c36 10 VSS 0.00219579f $X=0.216 $Y=0.216
c37 6 VSS 5.7036e-19 $X=0.233 $Y=0.216
c38 5 VSS 0.0042637f $X=0.162 $Y=0.054
c39 1 VSS 5.65078e-19 $X=0.179 $Y=0.054
r40 37 38 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.164 $X2=0.297 $Y2=0.1765
r41 35 36 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.07 $X2=0.297 $Y2=0.092
r42 34 37 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.114 $X2=0.297 $Y2=0.164
r43 34 36 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.114 $X2=0.297 $Y2=0.092
r44 32 38 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.1765
r45 31 35 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.07
r46 29 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.198 $X2=0.286 $Y2=0.198
r47 28 29 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.284 $Y2=0.198
r48 27 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.252 $Y2=0.198
r49 24 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.234 $Y2=0.198
r50 22 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.198 $X2=0.297 $Y2=0.189
r51 22 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.286 $Y2=0.198
r52 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.27 $Y2=0.036
r53 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r54 18 19 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.036 $X2=0.234 $Y2=0.036
r55 17 18 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.202 $Y2=0.036
r56 16 17 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r57 13 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r58 11 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r59 11 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.27 $Y2=0.036
r60 10 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r61 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.216 $X2=0.216 $Y2=0.216
r62 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.216 $X2=0.216 $Y2=0.216
r63 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r64 2 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.054 $X2=0.162 $Y2=0.054
r65 1 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.054 $X2=0.162 $Y2=0.054
.ends


* END of "./AOI22xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI22xp33_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 Y
* 
* Y	Y
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 noxref_9 N_A1_M0_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_Y_M1_d N_A2_M1_g noxref_9 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 noxref_10 N_B2_M2_g N_Y_M2_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.027
M3 VSS N_B1_M3_g noxref_10 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 VDD N_A1_M4_g noxref_7 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M5 noxref_7 N_A2_M5_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M6 N_Y_M6_d N_B2_M6_g noxref_7 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M7 noxref_7 N_B1_M7_g N_Y_M7_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
*
* 
* .include "AOI22xp33_ASAP7_75t_L.pex.sp.AOI22XP33_ASAP7_75T_L.pxi"
* BEGIN of "./AOI22xp33_ASAP7_75t_L.pex.sp.AOI22XP33_ASAP7_75T_L.pxi"
* File: AOI22xp33_ASAP7_75t_L.pex.sp.AOI22XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:12:55 2017
* 
x_PM_AOI22XP33_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M4_g A1 N_A1_c_3_p
+ N_A1_c_12_p N_A1_c_13_p N_A1_c_4_p VSS PM_AOI22XP33_ASAP7_75T_L%A1
x_PM_AOI22XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_18_n N_A2_M5_g N_A2_c_19_n A2
+ N_A2_c_24_n VSS PM_AOI22XP33_ASAP7_75T_L%A2
x_PM_AOI22XP33_ASAP7_75T_L%B2 N_B2_M2_g N_B2_c_37_n N_B2_M6_g B2 VSS
+ PM_AOI22XP33_ASAP7_75T_L%B2
x_PM_AOI22XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_49_n N_B1_M7_g B1 VSS
+ PM_AOI22XP33_ASAP7_75T_L%B1
x_PM_AOI22XP33_ASAP7_75T_L%Y N_Y_M2_s N_Y_M1_d N_Y_c_58_n N_Y_M7_s N_Y_M6_d
+ N_Y_c_69_n N_Y_c_57_n N_Y_c_61_n N_Y_c_63_n N_Y_c_59_n N_Y_c_65_n N_Y_c_75_n Y
+ N_Y_c_67_n VSS PM_AOI22XP33_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00315405f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A1_c_2_p N_A2_c_18_n 0.00120928f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p N_A2_c_19_n 8.78098e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A1_c_4_p N_A2_c_19_n 9.21192e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.135
cc_5 N_A1_M0_g A2 2.31533e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.186
cc_6 A1 A2 6.2884e-19 $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.186
cc_7 N_A1_c_3_p A2 3.4185e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.186
cc_8 A1 N_A2_c_24_n 8.11421e-19 $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.164
cc_9 N_A1_M0_g N_B2_M2_g 2.60137e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_10 VSS A1 0.00128285f $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.135
cc_11 VSS A1 7.45437e-19 $X=0.018 $Y=0.151 $X2=0 $Y2=0
cc_12 VSS N_A1_c_12_p 2.52895e-19 $X=0.046 $Y=0.135 $X2=0 $Y2=0
cc_13 VSS N_A1_c_13_p 2.52895e-19 $X=0.0635 $Y=0.135 $X2=0 $Y2=0
cc_14 VSS N_A1_M0_g 2.94699e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_15 VSS N_A1_c_3_p 2.52895e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_16 N_A1_c_4_p N_Y_c_57_n 2.6601e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.135
cc_17 N_A2_M1_g N_B2_M2_g 0.00353901f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_18 N_A2_c_18_n N_B2_c_37_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_19 N_A2_c_19_n B2 0.00443545f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_20 N_A2_M1_g N_B1_M3_g 2.949e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_21 VSS A2 3.93816e-19 $X=0.135 $Y=0.186 $X2=0.081 $Y2=0.135
cc_22 VSS A2 6.22427e-19 $X=0.135 $Y=0.186 $X2=0 $Y2=0
cc_23 VSS N_A2_M1_g 2.38303e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_24 VSS A2 0.00549565f $X=0.135 $Y=0.186 $X2=0 $Y2=0
cc_25 N_A2_c_19_n N_Y_c_58_n 3.87865e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_26 A2 N_Y_c_59_n 4.39597e-19 $X=0.135 $Y=0.186 $X2=0.018 $Y2=0.135
cc_27 N_B2_M2_g N_B1_M3_g 0.00358983f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_28 N_B2_c_37_n N_B1_c_49_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_29 B2 B1 0.00490704f $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_30 VSS N_B2_M2_g 3.57119e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_31 VSS B2 5.37372e-19 $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_32 B2 N_Y_c_58_n 3.87865e-19 $X=0.188 $Y=0.115 $X2=0.081 $Y2=0.135
cc_33 N_B2_M2_g N_Y_c_61_n 2.64276e-19 $X=0.189 $Y=0.054 $X2=0.027 $Y2=0.135
cc_34 B2 N_Y_c_61_n 0.00124805f $X=0.188 $Y=0.115 $X2=0.027 $Y2=0.135
cc_35 VSS N_B1_M3_g 2.08515e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_36 N_B1_M3_g N_Y_c_63_n 2.56935e-19 $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.186
cc_37 B1 N_Y_c_63_n 0.00123064f $X=0.245 $Y=0.081 $X2=0.135 $Y2=0.186
cc_38 N_B1_M3_g N_Y_c_65_n 2.76185e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_39 B1 N_Y_c_65_n 0.0012322f $X=0.245 $Y=0.081 $X2=0 $Y2=0
cc_40 B1 N_Y_c_67_n 0.00445461f $X=0.245 $Y=0.081 $X2=0 $Y2=0
cc_41 VSS N_Y_c_58_n 6.80422e-19 $X=0.162 $Y=0.216 $X2=0.081 $Y2=0.135
cc_42 VSS N_Y_c_69_n 0.00288888f $X=0.162 $Y=0.216 $X2=0 $Y2=0
cc_43 VSS N_Y_c_69_n 0.00302498f $X=0.268 $Y=0.216 $X2=0 $Y2=0
cc_44 VSS N_Y_c_69_n 0.00250965f $X=0.236 $Y=0.234 $X2=0 $Y2=0
cc_45 VSS N_Y_c_59_n 3.96143e-19 $X=0.162 $Y=0.216 $X2=0.018 $Y2=0.135
cc_46 VSS N_Y_c_59_n 0.00352873f $X=0.236 $Y=0.234 $X2=0.018 $Y2=0.135
cc_47 VSS N_Y_c_65_n 0.00352873f $X=0.27 $Y=0.234 $X2=0 $Y2=0
cc_48 VSS N_Y_c_75_n 0.00395609f $X=0.268 $Y=0.216 $X2=0 $Y2=0

* END of "./AOI22xp33_ASAP7_75t_L.pex.sp.AOI22XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI22xp5_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:13:17 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI22xp5_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI22xp5_ASAP7_75t_L.pex.sp.pex"
* File: AOI22xp5_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:13:17 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI22XP5_ASAP7_75T_L%A1 2 5 7 16 19 21 22 26 VSS
c14 26 VSS 0.0125858f $X=0.027 $Y=0.135
c15 22 VSS 5.72913e-19 $X=0.068 $Y=0.135
c16 21 VSS 8.17289e-19 $X=0.055 $Y=0.135
c17 19 VSS 7.99362e-19 $X=0.081 $Y=0.135
c18 16 VSS 0.00416161f $X=0.018 $Y=0.151
c19 5 VSS 0.00273954f $X=0.081 $Y=0.135
c20 2 VSS 0.0645488f $X=0.081 $Y=0.0675
r21 21 22 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.055
+ $Y=0.135 $X2=0.068 $Y2=0.135
r22 19 22 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.068 $Y2=0.135
r23 17 26 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.135 $X2=0.027 $Y2=0.135
r24 17 21 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.135 $X2=0.055 $Y2=0.135
r25 13 26 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.144 $X2=0.027 $Y2=0.135
r26 13 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.144 $X2=0.027 $Y2=0.151
r27 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r28 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r29 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI22XP5_ASAP7_75T_L%A2 2 5 7 11 17 19 VSS
c15 19 VSS 2.36257e-19 $X=0.135 $Y=0.164
c16 17 VSS 0.00288932f $X=0.135 $Y=0.186
c17 11 VSS 0.00139379f $X=0.135 $Y=0.135
c18 5 VSS 0.00128392f $X=0.135 $Y=0.135
c19 2 VSS 0.0602909f $X=0.135 $Y=0.0675
r20 18 19 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.164
r21 17 19 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.186 $X2=0.135 $Y2=0.164
r22 11 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r23 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r24 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r25 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI22XP5_ASAP7_75T_L%B2 2 5 7 10 VSS
c12 10 VSS 5.22847e-19 $X=0.188 $Y=0.115
c13 5 VSS 0.00110682f $X=0.189 $Y=0.135
c14 2 VSS 0.0604449f $X=0.189 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI22XP5_ASAP7_75T_L%B1 2 5 7 10 VSS
c10 10 VSS 0.00165942f $X=0.245 $Y=0.081
c11 5 VSS 0.00170643f $X=0.243 $Y=0.135
c12 2 VSS 0.0641824f $X=0.243 $Y=0.0675
r13 10 13 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.135
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI22XP5_ASAP7_75T_L%Y 1 2 6 7 10 14 16 17 19 20 27 28 29 34 36 VSS
c21 38 VSS 5.39703e-19 $X=0.297 $Y=0.1765
c22 36 VSS 0.00102781f $X=0.297 $Y=0.092
c23 35 VSS 0.00131846f $X=0.297 $Y=0.07
c24 34 VSS 0.00328923f $X=0.297 $Y=0.114
c25 32 VSS 6.07272e-19 $X=0.297 $Y=0.189
c26 30 VSS 1.42799e-19 $X=0.286 $Y=0.198
c27 29 VSS 5.14525e-19 $X=0.284 $Y=0.198
c28 28 VSS 8.46035e-21 $X=0.252 $Y=0.198
c29 27 VSS 4.59335e-19 $X=0.234 $Y=0.198
c30 22 VSS 0.00199921f $X=0.288 $Y=0.198
c31 21 VSS 0.00331385f $X=0.27 $Y=0.036
c32 20 VSS 0.00142296f $X=0.252 $Y=0.036
c33 19 VSS 0.00291823f $X=0.234 $Y=0.036
c34 18 VSS 4.13316e-19 $X=0.202 $Y=0.036
c35 17 VSS 0.00146362f $X=0.198 $Y=0.036
c36 16 VSS 0.00392404f $X=0.18 $Y=0.036
c37 14 VSS 0.00501635f $X=0.162 $Y=0.036
c38 11 VSS 0.0062054f $X=0.288 $Y=0.036
c39 10 VSS 0.00243084f $X=0.216 $Y=0.2025
c40 6 VSS 5.75997e-19 $X=0.233 $Y=0.2025
c41 1 VSS 5.72268e-19 $X=0.179 $Y=0.0675
r42 37 38 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.164 $X2=0.297 $Y2=0.1765
r43 35 36 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.07 $X2=0.297 $Y2=0.092
r44 34 37 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.114 $X2=0.297 $Y2=0.164
r45 34 36 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.114 $X2=0.297 $Y2=0.092
r46 32 38 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.1765
r47 31 35 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.07
r48 29 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.198 $X2=0.286 $Y2=0.198
r49 28 29 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.284 $Y2=0.198
r50 27 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.252 $Y2=0.198
r51 24 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.234 $Y2=0.198
r52 22 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.198 $X2=0.297 $Y2=0.189
r53 22 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.286 $Y2=0.198
r54 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.27 $Y2=0.036
r55 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r56 18 19 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.036 $X2=0.234 $Y2=0.036
r57 17 18 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.202 $Y2=0.036
r58 16 17 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r59 13 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r60 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r61 11 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r62 11 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.27 $Y2=0.036
r63 10 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r64 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r65 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r66 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r67 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.0675 $X2=0.162 $Y2=0.0675
r68 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.162 $Y2=0.0675
.ends


* END of "./AOI22xp5_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI22xp5_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 Y
* 
* Y	Y
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 noxref_9 N_A1_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_Y_M1_d N_A2_M1_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_10 N_B2_M2_g N_Y_M2_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_B1_M3_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 VDD N_A1_M4_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 noxref_7 N_A2_M5_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 N_Y_M6_d N_B2_M6_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M7 noxref_7 N_B1_M7_g N_Y_M7_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
*
* 
* .include "AOI22xp5_ASAP7_75t_L.pex.sp.AOI22XP5_ASAP7_75T_L.pxi"
* BEGIN of "./AOI22xp5_ASAP7_75t_L.pex.sp.AOI22XP5_ASAP7_75T_L.pxi"
* File: AOI22xp5_ASAP7_75t_L.pex.sp.AOI22XP5_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:13:17 2017
* 
x_PM_AOI22XP5_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M4_g A1 N_A1_c_3_p
+ N_A1_c_11_p N_A1_c_13_p N_A1_c_4_p VSS PM_AOI22XP5_ASAP7_75T_L%A1
x_PM_AOI22XP5_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_16_n N_A2_M5_g N_A2_c_17_n A2
+ N_A2_c_20_n VSS PM_AOI22XP5_ASAP7_75T_L%A2
x_PM_AOI22XP5_ASAP7_75T_L%B2 N_B2_M2_g N_B2_c_32_n N_B2_M6_g B2 VSS
+ PM_AOI22XP5_ASAP7_75T_L%B2
x_PM_AOI22XP5_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_44_n N_B1_M7_g B1 VSS
+ PM_AOI22XP5_ASAP7_75T_L%B1
x_PM_AOI22XP5_ASAP7_75T_L%Y N_Y_M2_s N_Y_M1_d N_Y_M7_s N_Y_M6_d N_Y_c_63_n
+ N_Y_c_53_n N_Y_c_52_n N_Y_c_56_n N_Y_c_72_p N_Y_c_58_n N_Y_c_54_n N_Y_c_60_n
+ N_Y_c_70_n Y N_Y_c_62_n VSS PM_AOI22XP5_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00315405f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_16_n 0.00120426f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p N_A2_c_17_n 8.76278e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A1_c_4_p N_A2_c_17_n 7.48762e-19 $X=0.027 $Y=0.135 $X2=0.135 $Y2=0.135
cc_5 A1 A2 3.88222e-19 $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.186
cc_6 A1 N_A2_c_20_n 5.23575e-19 $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.164
cc_7 N_A1_M0_g N_B2_M2_g 2.60137e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_8 VSS A1 2.0764e-19 $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.0675
cc_9 VSS A1 0.00259659f $X=0.018 $Y=0.151 $X2=0.135 $Y2=0.135
cc_10 VSS A1 0.0017083f $X=0.018 $Y=0.151 $X2=0 $Y2=0
cc_11 VSS N_A1_c_11_p 3.81942e-19 $X=0.055 $Y=0.135 $X2=0 $Y2=0
cc_12 VSS N_A1_M0_g 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_13 VSS N_A1_c_13_p 3.81942e-19 $X=0.068 $Y=0.135 $X2=0 $Y2=0
cc_14 N_A1_c_4_p N_Y_c_52_n 2.82062e-19 $X=0.027 $Y=0.135 $X2=0.135 $Y2=0.186
cc_15 N_A2_M1_g N_B2_M2_g 0.00353901f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_A2_c_16_n N_B2_c_32_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_17 N_A2_c_17_n B2 0.00388913f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_18 N_A2_M1_g N_B1_M3_g 2.949e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_19 VSS N_A2_c_20_n 0.00123935f $X=0.135 $Y=0.164 $X2=0 $Y2=0
cc_20 VSS N_A2_M1_g 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0.027 $Y2=0.135
cc_21 VSS A2 0.003771f $X=0.135 $Y=0.186 $X2=0.027 $Y2=0.135
cc_22 N_A2_c_17_n N_Y_c_53_n 0.0013399f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_23 A2 N_Y_c_54_n 4.25731e-19 $X=0.135 $Y=0.186 $X2=0 $Y2=0
cc_24 N_B2_M2_g N_B1_M3_g 0.00358983f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_25 N_B2_c_32_n N_B1_c_44_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_26 B2 B1 0.00477924f $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_27 VSS N_B2_M2_g 3.57119e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_28 VSS B2 5.37372e-19 $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_29 B2 N_Y_c_53_n 0.0013399f $X=0.188 $Y=0.115 $X2=0 $Y2=0
cc_30 N_B2_M2_g N_Y_c_56_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0.036 $Y2=0.135
cc_31 B2 N_Y_c_56_n 0.00124805f $X=0.188 $Y=0.115 $X2=0.036 $Y2=0.135
cc_32 VSS N_B1_M3_g 2.08515e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_33 N_B1_M3_g N_Y_c_58_n 2.56935e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_34 B1 N_Y_c_58_n 0.00123064f $X=0.245 $Y=0.081 $X2=0 $Y2=0
cc_35 N_B1_M3_g N_Y_c_60_n 2.76185e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_36 B1 N_Y_c_60_n 0.0012322f $X=0.245 $Y=0.081 $X2=0 $Y2=0
cc_37 B1 N_Y_c_62_n 0.00391435f $X=0.245 $Y=0.081 $X2=0 $Y2=0
cc_38 VSS N_Y_c_63_n 0.00369767f $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_39 VSS N_Y_c_63_n 0.00371662f $X=0.268 $Y=0.2025 $X2=0 $Y2=0
cc_40 VSS N_Y_c_63_n 0.00250965f $X=0.236 $Y=0.234 $X2=0 $Y2=0
cc_41 VSS N_Y_c_53_n 0.00107252f $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_42 VSS N_Y_c_54_n 3.96143e-19 $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_43 VSS N_Y_c_54_n 0.00352872f $X=0.236 $Y=0.234 $X2=0 $Y2=0
cc_44 VSS N_Y_c_60_n 0.00352872f $X=0.27 $Y=0.234 $X2=0 $Y2=0
cc_45 VSS N_Y_c_70_n 0.00284922f $X=0.268 $Y=0.2025 $X2=0 $Y2=0
cc_46 VSS Y 3.3721e-19 $X=0.268 $Y=0.2025 $X2=0 $Y2=0
cc_47 VSS N_Y_c_72_p 3.19955e-19 $X=0.234 $Y=0.036 $X2=0.081 $Y2=0.0675

* END of "./AOI22xp5_ASAP7_75t_L.pex.sp.AOI22XP5_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI311xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:13:40 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI311xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI311xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI311xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:13:40 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI311XP33_ASAP7_75T_L%A3 2 5 7 17 VSS
c5 17 VSS 0.0181247f $X=0.08 $Y=0.136
c6 5 VSS 0.00275452f $X=0.081 $Y=0.135
c7 2 VSS 0.0643308f $X=0.081 $Y=0.0675
r8 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r9 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r10 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI311XP33_ASAP7_75T_L%A2 2 5 7 17 VSS
c12 17 VSS 0.0040251f $X=0.134 $Y=0.136
c13 5 VSS 0.00131688f $X=0.135 $Y=0.135
c14 2 VSS 0.0597711f $X=0.135 $Y=0.0675
r15 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI311XP33_ASAP7_75T_L%A1 2 5 7 13 VSS
c13 13 VSS 0.0021029f $X=0.196 $Y=0.136
c14 5 VSS 0.00118479f $X=0.189 $Y=0.135
c15 2 VSS 0.0604741f $X=0.189 $Y=0.0675
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI311XP33_ASAP7_75T_L%B 2 5 7 13 VSS
c11 13 VSS 0.00135757f $X=0.247 $Y=0.134
c12 5 VSS 0.00123712f $X=0.243 $Y=0.135
c13 2 VSS 0.0620606f $X=0.243 $Y=0.054
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI311XP33_ASAP7_75T_L%C 2 5 7 10 VSS
c9 10 VSS 0.00137012f $X=0.297 $Y=0.134
c10 5 VSS 0.00179274f $X=0.297 $Y=0.135
c11 2 VSS 0.0660915f $X=0.297 $Y=0.054
r12 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r14 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AOI311XP33_ASAP7_75T_L%Y 2 3 5 8 15 18 23 26 27 28 34 39 45 VSS
c14 45 VSS 0.00384059f $X=0.342 $Y=0.234
c15 44 VSS 0.00278493f $X=0.351 $Y=0.234
c16 39 VSS 0.00565612f $X=0.351 $Y=0.2
c17 38 VSS 9.05161e-19 $X=0.351 $Y=0.07
c18 37 VSS 0.00126f $X=0.351 $Y=0.225
c19 35 VSS 4.19362e-19 $X=0.31 $Y=0.036
c20 34 VSS 0.00142296f $X=0.306 $Y=0.036
c21 33 VSS 0.00632503f $X=0.288 $Y=0.036
c22 32 VSS 0.00100794f $X=0.252 $Y=0.036
c23 28 VSS 6.7196e-19 $X=0.241 $Y=0.036
c24 27 VSS 0.00434692f $X=0.234 $Y=0.036
c25 23 VSS 0.00474875f $X=0.216 $Y=0.036
c26 20 VSS 0.00657518f $X=0.342 $Y=0.036
c27 18 VSS 0.00262708f $X=0.322 $Y=0.2025
c28 8 VSS 0.00574947f $X=0.322 $Y=0.054
c29 4 VSS 5.36031e-19 $X=0.216 $Y=0.0455
r30 45 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.3465 $Y2=0.234
r31 44 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.234 $X2=0.3465 $Y2=0.234
r32 41 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.342 $Y2=0.234
r33 38 39 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.07 $X2=0.351 $Y2=0.2
r34 37 44 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.234
r35 37 39 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.2
r36 36 38 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.07
r37 34 35 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.31 $Y2=0.036
r38 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r39 32 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r40 30 35 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.31 $Y2=0.036
r41 27 28 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.241 $Y2=0.036
r42 26 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.036 $X2=0.252 $Y2=0.036
r43 26 28 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.036 $X2=0.241 $Y2=0.036
r44 22 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.234 $Y2=0.036
r45 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r46 20 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.036 $X2=0.351 $Y2=0.045
r47 20 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.324 $Y2=0.036
r48 18 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r49 15 18 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.322 $Y2=0.2025
r50 14 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r51 8 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r52 5 8 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.054 $X2=0.322 $Y2=0.054
r53 3 4 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0455 $X2=0.216 $Y2=0.0455
r54 2 4 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0455 $X2=0.216 $Y2=0.0455
r55 1 14 3.12934 $w=6.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.216 $Y=0.064 $X2=0.199 $Y2=0.064
r56 1 4 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.216 $Y=0.064 $X2=0.216 $Y2=0.0455
.ends


* END of "./AOI311xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI311xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 B C Y
* 
* Y	Y
* C	C
* B	B
* A1	A1
* A2	A2
* A3	A3
M0 noxref_10 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_11 N_A2_M1_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_A1_M2_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_B_M3_g N_Y_M3_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_C_M4_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287 $Y=0.027
M5 noxref_8 N_A3_M5_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M6 VDD N_A2_M6_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 noxref_8 N_A1_M7_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M8 noxref_12 N_B_M8_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M9 N_Y_M9_d N_C_M9_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
*
* 
* .include "AOI311xp33_ASAP7_75t_L.pex.sp.AOI311XP33_ASAP7_75T_L.pxi"
* BEGIN of "./AOI311xp33_ASAP7_75t_L.pex.sp.AOI311XP33_ASAP7_75T_L.pxi"
* File: AOI311xp33_ASAP7_75t_L.pex.sp.AOI311XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:13:40 2017
* 
x_PM_AOI311XP33_ASAP7_75T_L%A3 N_A3_M0_g N_A3_c_2_p N_A3_M5_g A3 VSS
+ PM_AOI311XP33_ASAP7_75T_L%A3
x_PM_AOI311XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_7_n N_A2_M6_g A2 VSS
+ PM_AOI311XP33_ASAP7_75T_L%A2
x_PM_AOI311XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_20_n N_A1_M7_g A1 VSS
+ PM_AOI311XP33_ASAP7_75T_L%A1
x_PM_AOI311XP33_ASAP7_75T_L%B N_B_M3_g N_B_c_33_n N_B_M8_g B VSS
+ PM_AOI311XP33_ASAP7_75T_L%B
x_PM_AOI311XP33_ASAP7_75T_L%C N_C_M4_g N_C_c_44_n N_C_M9_g C VSS
+ PM_AOI311XP33_ASAP7_75T_L%C
x_PM_AOI311XP33_ASAP7_75T_L%Y N_Y_M3_s N_Y_M2_d N_Y_M4_d N_Y_c_57_n N_Y_M9_d
+ N_Y_c_58_n N_Y_c_51_n Y N_Y_c_52_n N_Y_c_56_n N_Y_c_59_n N_Y_c_61_n N_Y_c_64_n
+ VSS PM_AOI311XP33_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_A2_M1_g 0.00347357f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A3_c_2_p N_A2_c_7_n 0.00120426f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A3 A2 0.0026877f $X=0.08 $Y=0.136 $X2=0.134 $Y2=0.136
cc_4 N_A3_M0_g N_A1_M2_g 2.69148e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 VSS A3 2.10206e-19 $X=0.08 $Y=0.136 $X2=0 $Y2=0
cc_6 N_A2_M1_g N_A1_M2_g 0.00325575f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_7 N_A2_c_7_n N_A1_c_20_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_8 A2 A1 0.00564452f $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_9 N_A2_M1_g N_B_M3_g 2.69148e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_10 VSS A2 0.00132451f $X=0.134 $Y=0.136 $X2=0.081 $Y2=0.135
cc_11 VSS N_A2_M1_g 2.64276e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_12 VSS A2 0.00125674f $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_13 A2 N_Y_c_51_n 7.91188e-19 $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_14 A2 N_Y_c_52_n 4.76378e-19 $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_15 N_A1_M2_g N_B_M3_g 0.00359705f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_A1_c_20_n N_B_c_33_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_17 A1 B 0.00506253f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_18 N_A1_M2_g N_C_M4_g 2.69148e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_19 VSS A1 0.00114532f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_20 VSS N_A1_M2_g 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_21 VSS A1 0.00125352f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_22 A1 N_Y_c_51_n 0.0013295f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_23 N_A1_M2_g N_Y_c_52_n 2.80442e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 N_B_M3_g N_C_M4_g 0.00330657f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.0675
cc_25 N_B_c_33_n N_C_c_44_n 9.33263e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_26 B C 0.00624003f $X=0.247 $Y=0.134 $X2=0.135 $Y2=0.135
cc_27 VSS B 0.0013399f $X=0.247 $Y=0.134 $X2=0.135 $Y2=0.135
cc_28 VSS N_B_M3_g 3.06796e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_29 B N_Y_c_51_n 0.00127618f $X=0.247 $Y=0.134 $X2=0 $Y2=0
cc_30 B N_Y_c_56_n 0.00123604f $X=0.247 $Y=0.134 $X2=0 $Y2=0
cc_31 C N_Y_c_57_n 3.31541e-19 $X=0.297 $Y=0.134 $X2=0 $Y2=0
cc_32 C N_Y_c_58_n 0.0013399f $X=0.297 $Y=0.134 $X2=0 $Y2=0
cc_33 N_C_M4_g N_Y_c_59_n 2.56935e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_34 C N_Y_c_59_n 0.00123604f $X=0.297 $Y=0.134 $X2=0 $Y2=0
cc_35 C N_Y_c_61_n 0.00546796f $X=0.297 $Y=0.134 $X2=0 $Y2=0
cc_36 VSS N_Y_c_58_n 0.00147748f $X=0.216 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_37 VSS N_Y_c_51_n 0.00107252f $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_38 VSS N_Y_c_64_n 4.51619e-19 $X=0.216 $Y=0.234 $X2=0 $Y2=0

* END of "./AOI311xp33_ASAP7_75t_L.pex.sp.AOI311XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI31xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:14:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI31xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI31xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI31xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:14:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI31XP33_ASAP7_75T_L%A3 2 5 7 13 VSS
c5 13 VSS 0.00742663f $X=0.0855 $Y=0.1355
c6 5 VSS 0.00298625f $X=0.081 $Y=0.135
c7 2 VSS 0.0631569f $X=0.081 $Y=0.0675
r8 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.134 $X2=0.081
+ $Y2=0.134
r9 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r10 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI31XP33_ASAP7_75T_L%A2 2 5 7 15 VSS
c12 15 VSS 0.00230441f $X=0.1355 $Y=0.1355
c13 5 VSS 0.00178389f $X=0.135 $Y=0.135
c14 2 VSS 0.0597711f $X=0.135 $Y=0.0675
r15 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.134 $X2=0.135
+ $Y2=0.134
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI31XP33_ASAP7_75T_L%A1 2 5 7 13 VSS
c13 13 VSS 0.00151062f $X=0.1895 $Y=0.1355
c14 5 VSS 0.00178389f $X=0.189 $Y=0.135
c15 2 VSS 0.0607397f $X=0.189 $Y=0.0675
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.134 $X2=0.189
+ $Y2=0.134
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI31XP33_ASAP7_75T_L%B 2 5 7 10 VSS
c8 10 VSS 0.00118636f $X=0.2405 $Y=0.1355
c9 5 VSS 0.00234817f $X=0.243 $Y=0.135
c10 2 VSS 0.0655182f $X=0.243 $Y=0.054
r11 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.134 $X2=0.243
+ $Y2=0.134
r12 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r13 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI31XP33_ASAP7_75T_L%Y 2 3 6 10 13 20 22 27 29 31 37 VSS
c13 37 VSS 0.00203647f $X=0.288 $Y=0.198
c14 36 VSS 0.00163204f $X=0.297 $Y=0.198
c15 31 VSS 5.57912e-19 $X=0.297 $Y=0.1765
c16 29 VSS 9.04922e-19 $X=0.297 $Y=0.0905
c17 28 VSS 0.00142953f $X=0.297 $Y=0.07
c18 27 VSS 0.0032767f $X=0.299 $Y=0.111
c19 25 VSS 7.58409e-19 $X=0.297 $Y=0.189
c20 23 VSS 3.86697e-19 $X=0.256 $Y=0.036
c21 22 VSS 0.00142432f $X=0.252 $Y=0.036
c22 21 VSS 4.1452e-19 $X=0.234 $Y=0.036
c23 20 VSS 0.0039184f $X=0.23 $Y=0.036
c24 15 VSS 0.0088253f $X=0.288 $Y=0.036
c25 13 VSS 0.00174116f $X=0.268 $Y=0.216
c26 6 VSS 0.00531813f $X=0.205 $Y=0.028
r27 37 38 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.2925 $Y2=0.198
r28 36 38 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.198 $X2=0.2925 $Y2=0.198
r29 33 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.198 $X2=0.288 $Y2=0.198
r30 30 31 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.164 $X2=0.297 $Y2=0.1765
r31 28 29 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.07 $X2=0.297 $Y2=0.0905
r32 27 30 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.111 $X2=0.297 $Y2=0.164
r33 27 29 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.111 $X2=0.297 $Y2=0.0905
r34 25 36 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.198
r35 25 31 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.1765
r36 24 28 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.07
r37 22 23 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.256 $Y2=0.036
r38 21 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r39 20 21 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.036 $X2=0.234 $Y2=0.036
r40 17 20 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.23 $Y2=0.036
r41 15 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r42 15 23 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.256 $Y2=0.036
r43 13 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.198 $X2=0.27
+ $Y2=0.198
r44 10 13 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.216 $X2=0.268 $Y2=0.216
r45 6 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r46 3 6 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0455 $X2=0.216 $Y2=0.0455
r47 2 6 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0455 $X2=0.216 $Y2=0.0455
.ends


* END of "./AOI31xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI31xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 B Y
* 
* Y	Y
* B	B
* A1	A1
* A2	A2
* A3	A3
M0 noxref_9 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_10 N_A2_M1_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_A1_M2_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_B_M3_g N_Y_M3_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 noxref_7 N_A3_M4_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M5 VDD N_A2_M5_g noxref_7 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M6 noxref_7 N_A1_M6_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M7 N_Y_M7_d N_B_M7_g noxref_7 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
*
* 
* .include "AOI31xp33_ASAP7_75t_L.pex.sp.AOI31XP33_ASAP7_75T_L.pxi"
* BEGIN of "./AOI31xp33_ASAP7_75t_L.pex.sp.AOI31XP33_ASAP7_75T_L.pxi"
* File: AOI31xp33_ASAP7_75t_L.pex.sp.AOI31XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:14:03 2017
* 
x_PM_AOI31XP33_ASAP7_75T_L%A3 N_A3_M0_g N_A3_c_2_p N_A3_M4_g A3 VSS
+ PM_AOI31XP33_ASAP7_75T_L%A3
x_PM_AOI31XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_7_n N_A2_M5_g A2 VSS
+ PM_AOI31XP33_ASAP7_75T_L%A2
x_PM_AOI31XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_20_n N_A1_M6_g A1 VSS
+ PM_AOI31XP33_ASAP7_75T_L%A1
x_PM_AOI31XP33_ASAP7_75T_L%B N_B_M3_g N_B_c_33_n N_B_M7_g B VSS
+ PM_AOI31XP33_ASAP7_75T_L%B
x_PM_AOI31XP33_ASAP7_75T_L%Y N_Y_M3_s N_Y_M2_d N_Y_c_39_n N_Y_M7_d N_Y_c_49_n
+ N_Y_c_40_n N_Y_c_45_n Y N_Y_c_47_n N_Y_c_42_n N_Y_c_43_n VSS
+ PM_AOI31XP33_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_A2_M1_g 0.00347357f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A3_c_2_p N_A2_c_7_n 9.56181e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A3 A2 0.00802362f $X=0.0855 $Y=0.1355 $X2=0.1355 $Y2=0.1355
cc_4 N_A3_M0_g N_A1_M2_g 2.69148e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 VSS A3 3.31541e-19 $X=0.0855 $Y=0.1355 $X2=0.135 $Y2=0.135
cc_6 N_A2_M1_g N_A1_M2_g 0.00325575f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_7 N_A2_c_7_n N_A1_c_20_n 9.07968e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_8 A2 A1 0.00613955f $X=0.1355 $Y=0.1355 $X2=0.0855 $Y2=0.1355
cc_9 N_A2_M1_g N_B_M3_g 2.69148e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_10 VSS A2 3.31541e-19 $X=0.1355 $Y=0.1355 $X2=0.081 $Y2=0.135
cc_11 VSS N_A2_M1_g 2.64276e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_12 VSS A2 0.00125674f $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_13 A2 N_Y_c_39_n 7.56932e-19 $X=0.1355 $Y=0.1355 $X2=0.081 $Y2=0.216
cc_14 A2 N_Y_c_40_n 4.56622e-19 $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_15 N_A1_M2_g N_B_M3_g 0.00359705f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_A1_c_20_n N_B_c_33_n 9.56181e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_17 A1 B 0.00393834f $X=0.1895 $Y=0.1355 $X2=0.081 $Y2=0.134
cc_18 VSS A1 3.61412e-19 $X=0.1895 $Y=0.1355 $X2=0.081 $Y2=0.134
cc_19 VSS N_A1_M2_g 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_20 VSS A1 0.00125352f $X=0.1895 $Y=0.1355 $X2=0 $Y2=0
cc_21 A1 N_Y_c_39_n 0.0013295f $X=0.1895 $Y=0.1355 $X2=0.081 $Y2=0.216
cc_22 A1 N_Y_c_42_n 5.26804e-19 $X=0.1895 $Y=0.1355 $X2=0 $Y2=0
cc_23 A1 N_Y_c_43_n 2.59217e-19 $X=0.1895 $Y=0.1355 $X2=0 $Y2=0
cc_24 B N_Y_c_39_n 0.00127618f $X=0.2405 $Y=0.1355 $X2=0.135 $Y2=0.216
cc_25 N_B_M3_g N_Y_c_45_n 2.56935e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_26 B N_Y_c_45_n 0.00123064f $X=0.2405 $Y=0.1355 $X2=0 $Y2=0
cc_27 B N_Y_c_47_n 0.00441786f $X=0.2405 $Y=0.1355 $X2=0 $Y2=0
cc_28 VSS N_Y_c_39_n 9.28287e-19 $X=0.216 $Y=0.216 $X2=0.081 $Y2=0.216
cc_29 VSS N_Y_c_49_n 0.002591f $X=0.216 $Y=0.216 $X2=0.0855 $Y2=0.1355
cc_30 VSS N_Y_c_49_n 3.09692e-19 $X=0.216 $Y=0.234 $X2=0.0855 $Y2=0.1355
cc_31 VSS N_Y_c_43_n 3.59474e-19 $X=0.216 $Y=0.216 $X2=0 $Y2=0

* END of "./AOI31xp33_ASAP7_75t_L.pex.sp.AOI31XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI31xp67_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:14:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI31xp67_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI31xp67_ASAP7_75t_L.pex.sp.pex"
* File: AOI31xp67_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:14:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI31XP67_ASAP7_75T_L%A3 2 7 10 13 15 25 VSS
c18 25 VSS 0.0201929f $X=0.08 $Y=0.136
c19 13 VSS 0.0077404f $X=0.135 $Y=0.135
c20 10 VSS 0.063053f $X=0.135 $Y=0.0675
c21 2 VSS 0.0670913f $X=0.081 $Y=0.0675
r22 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r23 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r24 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r25 5 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI31XP67_ASAP7_75T_L%B 2 7 10 13 21 VSS
c31 21 VSS 0.00662363f $X=0.189 $Y=0.134
c32 10 VSS 0.0724844f $X=0.243 $Y=0.135
c33 2 VSS 0.0623453f $X=0.189 $Y=0.054
r34 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r35 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r36 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r37 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r38 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI31XP67_ASAP7_75T_L%A2 2 7 10 13 15 23 VSS
c29 23 VSS 0.0060928f $X=0.403 $Y=0.137
c30 13 VSS 0.00396437f $X=0.459 $Y=0.134
c31 10 VSS 0.0632471f $X=0.459 $Y=0.0675
c32 2 VSS 0.0665454f $X=0.405 $Y=0.0675
r33 13 15 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.134 $X2=0.459 $Y2=0.2025
r34 10 13 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.134
r35 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.134 $X2=0.459 $Y2=0.134
r36 5 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r37 5 7 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.134 $X2=0.405 $Y2=0.2025
r38 2 5 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.134
.ends

.subckt PM_AOI31XP67_ASAP7_75T_L%A1 2 7 10 13 15 22 VSS
c25 22 VSS 0.0108315f $X=0.569 $Y=0.137
c26 13 VSS 0.00311578f $X=0.567 $Y=0.135
c27 10 VSS 0.0668479f $X=0.567 $Y=0.0675
c28 2 VSS 0.0632472f $X=0.513 $Y=0.0675
r29 13 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r30 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r31 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r32 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r33 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r34 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AOI31XP67_ASAP7_75T_L%Y 1 4 6 7 11 12 15 18 19 20 22 23 24 25 26 27
+ 29 32 35 36 37 38 42 44 48 57 60 VSS
c62 66 VSS 1.77025e-19 $X=0.234 $Y=0.198
c63 60 VSS 4.02348e-20 $X=0.216 $Y=0.198
c64 57 VSS 1.58409e-19 $X=0.248 $Y=0.077
c65 54 VSS 2.67452e-19 $X=0.234 $Y=0.072
c66 48 VSS 4.77205e-19 $X=0.216 $Y=0.072
c67 44 VSS 0.00707584f $X=0.649 $Y=0.234
c68 42 VSS 0.00347422f $X=0.603 $Y=0.234
c69 41 VSS 6.42934e-19 $X=0.594 $Y=0.225
c70 38 VSS 0.00213769f $X=0.6285 $Y=0.036
c71 37 VSS 0.00695364f $X=0.608 $Y=0.036
c72 36 VSS 0.110791f $X=0.649 $Y=0.036
c73 35 VSS 0.00387584f $X=0.649 $Y=0.036
c74 32 VSS 0.00283143f $X=0.54 $Y=0.036
c75 29 VSS 4.75468e-19 $X=0.5695 $Y=0.198
c76 27 VSS 0.00277828f $X=0.553 $Y=0.198
c77 26 VSS 0.00413098f $X=0.419 $Y=0.198
c78 25 VSS 3.08827e-19 $X=0.306 $Y=0.198
c79 24 VSS 4.75287e-19 $X=0.288 $Y=0.198
c80 23 VSS 1.43629e-19 $X=0.252 $Y=0.198
c81 22 VSS 0.00248469f $X=0.585 $Y=0.198
c82 21 VSS 3.11686e-20 $X=0.243 $Y=0.1765
c83 20 VSS 2.87569e-19 $X=0.243 $Y=0.164
c84 18 VSS 3.66662e-19 $X=0.243 $Y=0.126
c85 17 VSS 6.69317e-20 $X=0.243 $Y=0.189
c86 15 VSS 0.00295586f $X=0.216 $Y=0.2025
c87 11 VSS 5.61665e-19 $X=0.233 $Y=0.2025
c88 6 VSS 5.98552e-19 $X=0.557 $Y=0.0675
c89 4 VSS 0.00597532f $X=0.214 $Y=0.054
r90 66 67 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.2385 $Y2=0.198
r91 65 67 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.198 $X2=0.2385 $Y2=0.198
r92 60 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.234 $Y2=0.198
r93 54 55 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.2385 $Y2=0.072
r94 53 57 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.072 $X2=0.248 $Y2=0.072
r95 53 55 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.072 $X2=0.2385 $Y2=0.072
r96 48 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.072 $X2=0.234 $Y2=0.072
r97 44 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.649 $Y=0.234 $X2=0.649
+ $Y2=0.234
r98 42 44 3.12346 $w=1.8e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.603
+ $Y=0.234 $X2=0.649 $Y2=0.234
r99 41 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.594 $Y=0.225 $X2=0.603 $Y2=0.234
r100 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.207 $X2=0.594 $Y2=0.225
r101 37 38 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.608
+ $Y=0.036 $X2=0.6285 $Y2=0.036
r102 36 45 170.893 $w=2.4e-08 $l=1.98e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.649 $Y=0.036 $X2=0.649 $Y2=0.234
r103 35 38 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.649
+ $Y=0.036 $X2=0.6285 $Y2=0.036
r104 35 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.649 $Y=0.036
+ $X2=0.649 $Y2=0.036
r105 31 37 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.608 $Y2=0.036
r106 31 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r107 28 29 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.554
+ $Y=0.198 $X2=0.5695 $Y2=0.198
r108 27 28 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.553
+ $Y=0.198 $X2=0.554 $Y2=0.198
r109 26 27 9.09877 $w=1.8e-08 $l=1.34e-07 $layer=M1 $thickness=3.6e-08 $X=0.419
+ $Y=0.198 $X2=0.553 $Y2=0.198
r110 25 26 7.67284 $w=1.8e-08 $l=1.13e-07 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.198 $X2=0.419 $Y2=0.198
r111 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.306 $Y2=0.198
r112 23 65 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.243 $Y2=0.198
r113 23 24 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.288 $Y2=0.198
r114 22 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.585 $Y=0.198 $X2=0.594 $Y2=0.207
r115 22 29 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.198 $X2=0.5695 $Y2=0.198
r116 20 21 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.164 $X2=0.243 $Y2=0.1765
r117 19 20 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.144 $X2=0.243 $Y2=0.164
r118 18 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.144
r119 17 65 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.198
r120 17 21 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.1765
r121 16 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.072
r122 16 18 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.126
r123 15 60 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198
+ $X2=0.216 $Y2=0.198
r124 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r125 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r126 10 32 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r127 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r128 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r129 4 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072 $X2=0.216
+ $Y2=0.072
r130 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.054 $X2=0.214 $Y2=0.054
.ends


* END of "./AOI31xp67_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI31xp67_ASAP7_75t_L  VSS VDD A3 B A2 A1 Y
* 
* Y	Y
* A1	A1
* A2	A2
* B	B
* A3	A3
M0 noxref_8 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_8 N_A3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_B_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 noxref_8 N_A2_M3_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 noxref_8 N_A2_M4_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M5 N_Y_M5_d N_A1_M5_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M6 N_Y_M6_d N_A1_M6_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M7 VDD N_A3_M7_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M8 VDD N_A3_M8_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M9 N_Y_M9_d N_B_M9_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M10 N_Y_M10_d N_B_M10_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M11 noxref_7 N_A2_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M12 noxref_7 N_A2_M12_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M13 noxref_7 N_A1_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M14 noxref_7 N_A1_M14_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
*
* 
* .include "AOI31xp67_ASAP7_75t_L.pex.sp.AOI31XP67_ASAP7_75T_L.pxi"
* BEGIN of "./AOI31xp67_ASAP7_75t_L.pex.sp.AOI31XP67_ASAP7_75T_L.pxi"
* File: AOI31xp67_ASAP7_75t_L.pex.sp.AOI31XP67_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:14:25 2017
* 
x_PM_AOI31XP67_ASAP7_75T_L%A3 N_A3_M0_g N_A3_M7_g N_A3_M1_g N_A3_c_4_p N_A3_M8_g
+ A3 VSS PM_AOI31XP67_ASAP7_75T_L%A3
x_PM_AOI31XP67_ASAP7_75T_L%B N_B_M2_g N_B_M9_g N_B_c_21_n N_B_M10_g B VSS
+ PM_AOI31XP67_ASAP7_75T_L%B
x_PM_AOI31XP67_ASAP7_75T_L%A2 N_A2_M3_g N_A2_M11_g N_A2_M4_g N_A2_c_53_p
+ N_A2_M12_g A2 VSS PM_AOI31XP67_ASAP7_75T_L%A2
x_PM_AOI31XP67_ASAP7_75T_L%A1 N_A1_M5_g N_A1_M13_g N_A1_M6_g N_A1_c_82_n
+ N_A1_M14_g A1 VSS PM_AOI31XP67_ASAP7_75T_L%A1
x_PM_AOI31XP67_ASAP7_75T_L%Y N_Y_M2_d N_Y_c_104_n N_Y_M6_d N_Y_M5_d N_Y_M10_d
+ N_Y_M9_d N_Y_c_106_n N_Y_c_107_n N_Y_c_109_n N_Y_c_111_n N_Y_c_127_n
+ N_Y_c_144_n N_Y_c_145_n N_Y_c_120_n N_Y_c_121_n N_Y_c_124_n N_Y_c_130_n
+ N_Y_c_132_n N_Y_c_133_n N_Y_c_134_n N_Y_c_136_n N_Y_c_138_n N_Y_c_149_n
+ N_Y_c_139_n N_Y_c_113_n Y N_Y_c_115_n VSS PM_AOI31XP67_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_B_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.054
cc_2 N_A3_M1_g N_B_M2_g 0.00323392f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.054
cc_3 N_A3_M1_g N_B_c_21_n 2.69148e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_4 N_A3_c_4_p N_B_c_21_n 0.00149358f $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_5 N_A3_M1_g B 5.93459e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.134
cc_6 N_A3_c_4_p B 0.0032047f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.134
cc_7 A3 B 0.002207f $X=0.08 $Y=0.136 $X2=0.189 $Y2=0.134
cc_8 VSS A3 2.23359e-19 $X=0.08 $Y=0.136 $X2=0.189 $Y2=0.054
cc_9 VSS A3 0.00225004f $X=0.08 $Y=0.136 $X2=0.189 $Y2=0.135
cc_10 VSS A3 0.00179824f $X=0.08 $Y=0.136 $X2=0 $Y2=0
cc_11 VSS N_A3_M0_g 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_12 VSS N_A3_c_4_p 3.08494e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_13 VSS A3 2.73034e-19 $X=0.08 $Y=0.136 $X2=0 $Y2=0
cc_14 VSS N_A3_M1_g 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 VSS N_A3_c_4_p 3.80277e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.054
cc_16 VSS A3 5.97636e-19 $X=0.08 $Y=0.136 $X2=0.243 $Y2=0.2025
cc_17 VSS N_A3_c_4_p 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.2025
cc_18 VSS N_A3_M1_g 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 VSS B 0.00154715f $X=0.189 $Y=0.134 $X2=0.135 $Y2=0.0675
cc_20 VSS B 0.00375052f $X=0.189 $Y=0.134 $X2=0.081 $Y2=0.135
cc_21 VSS B 5.19988e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_22 VSS N_B_M2_g 4.28653e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_23 VSS B 5.19988e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_24 VSS N_B_c_21_n 2.08515e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_25 VSS B 0.002132f $X=0.189 $Y=0.134 $X2=0.135 $Y2=0.135
cc_26 VSS B 0.00374737f $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_27 VSS N_B_M2_g 4.28653e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_28 VSS B 0.00104433f $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_29 VSS N_B_c_21_n 2.34993e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_30 N_B_c_21_n N_Y_c_104_n 3.82299e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_31 N_B_c_21_n N_Y_M10_d 3.8028e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_32 N_B_c_21_n N_Y_c_106_n 9.18375e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_33 N_B_c_21_n N_Y_c_107_n 7.54008e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_34 B N_Y_c_107_n 6.4382e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_35 N_B_c_21_n N_Y_c_109_n 0.00127415f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_36 B N_Y_c_109_n 8.41056e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_37 N_B_c_21_n N_Y_c_111_n 4.86057e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_38 B N_Y_c_111_n 5.36365e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_39 N_B_c_21_n N_Y_c_113_n 4.02804e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_40 B N_Y_c_113_n 3.57329e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_41 N_B_c_21_n N_Y_c_115_n 4.39606e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_42 B N_Y_c_115_n 3.72423e-19 $X=0.189 $Y=0.134 $X2=0 $Y2=0
cc_43 N_A2_M3_g N_A1_M5_g 2.74891e-19 $X=0.405 $Y=0.0675 $X2=0.189 $Y2=0.054
cc_44 N_A2_M4_g N_A1_M5_g 0.00335739f $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.054
cc_45 N_A2_M4_g N_A1_M6_g 2.74891e-19 $X=0.459 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_46 N_A2_c_53_p N_A1_c_82_n 0.00160986f $X=0.459 $Y=0.134 $X2=0.243 $Y2=0.2025
cc_47 VSS N_A2_c_53_p 3.74175e-19 $X=0.459 $Y=0.134 $X2=0 $Y2=0
cc_48 VSS N_A2_c_53_p 7.60428e-19 $X=0.459 $Y=0.134 $X2=0 $Y2=0
cc_49 VSS N_A2_M3_g 2.65027e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_50 VSS N_A2_M4_g 2.65027e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_51 VSS A2 3.34314e-19 $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_52 VSS N_A2_c_53_p 4.31323e-19 $X=0.459 $Y=0.134 $X2=0.189 $Y2=0.2025
cc_53 VSS N_A2_M3_g 3.32113e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_54 VSS A2 3.79597e-19 $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_55 VSS N_A2_c_53_p 8.43851e-19 $X=0.459 $Y=0.134 $X2=0 $Y2=0
cc_56 VSS A2 0.00410107f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_57 VSS A2 3.79597e-19 $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_58 VSS A2 8.62688e-19 $X=0.403 $Y=0.137 $X2=0.189 $Y2=0.135
cc_59 VSS N_A2_M3_g 3.42779e-19 $X=0.405 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_60 VSS N_A2_c_53_p 9.74713e-19 $X=0.459 $Y=0.134 $X2=0.189 $Y2=0.135
cc_61 VSS A2 0.00362146f $X=0.403 $Y=0.137 $X2=0.189 $Y2=0.135
cc_62 VSS N_A2_M4_g 4.86079e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_63 A2 N_Y_c_107_n 0.00126829f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_64 A2 N_Y_c_109_n 0.00126829f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_65 A2 N_Y_c_111_n 0.00126829f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_66 A2 N_Y_c_120_n 0.00125876f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_67 N_A2_M3_g N_Y_c_121_n 3.33408e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_68 N_A2_c_53_p N_Y_c_121_n 7.41207e-19 $X=0.459 $Y=0.134 $X2=0 $Y2=0
cc_69 A2 N_Y_c_121_n 0.00408842f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_70 N_A2_M4_g N_Y_c_124_n 3.98183e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_71 A2 Y 0.00126829f $X=0.403 $Y=0.137 $X2=0 $Y2=0
cc_72 VSS N_A1_c_82_n 3.80413e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_73 VSS N_A1_c_82_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_74 VSS N_A1_M5_g 2.64781e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_75 VSS N_A1_M6_g 3.44437e-19 $X=0.567 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_76 VSS A1 0.0034871f $X=0.569 $Y=0.137 $X2=0.405 $Y2=0.135
cc_77 VSS N_A1_M5_g 4.89467e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_78 VSS N_A1_c_82_n 9.79091e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_79 N_A1_c_82_n N_Y_M6_d 4.22601e-19 $X=0.567 $Y=0.135 $X2=0.405 $Y2=0.2025
cc_80 A1 N_Y_c_127_n 2.13112e-19 $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_81 N_A1_M5_g N_Y_c_124_n 3.95247e-19 $X=0.513 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_82 N_A1_c_82_n N_Y_c_124_n 7.66668e-19 $X=0.567 $Y=0.135 $X2=0.405 $Y2=0.135
cc_83 N_A1_M6_g N_Y_c_130_n 2.69508e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_84 A1 N_Y_c_130_n 0.00159015f $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_85 N_A1_c_82_n N_Y_c_132_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_86 A1 N_Y_c_133_n 4.07063e-19 $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_87 N_A1_c_82_n N_Y_c_134_n 8.21731e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_88 A1 N_Y_c_134_n 0.00862815f $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_89 N_A1_M6_g N_Y_c_136_n 3.32713e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_90 A1 N_Y_c_136_n 4.07063e-19 $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_91 A1 N_Y_c_138_n 4.07063e-19 $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_92 A1 N_Y_c_139_n 0.00116925f $X=0.569 $Y=0.137 $X2=0 $Y2=0
cc_93 VSS N_Y_c_106_n 0.00392515f $X=0.162 $Y=0.2025 $X2=0.135 $Y2=0.2025
cc_94 VSS N_Y_c_106_n 0.00345036f $X=0.268 $Y=0.2025 $X2=0.135 $Y2=0.2025
cc_95 VSS N_Y_c_106_n 0.00249183f $X=0.236 $Y=0.234 $X2=0.135 $Y2=0.2025
cc_96 VSS N_Y_c_111_n 5.0548e-19 $X=0.268 $Y=0.2025 $X2=0 $Y2=0
cc_97 VSS N_Y_c_144_n 0.0143431f $X=0.54 $Y=0.234 $X2=0 $Y2=0
cc_98 VSS N_Y_c_145_n 0.00294986f $X=0.268 $Y=0.2025 $X2=0 $Y2=0
cc_99 VSS N_Y_c_124_n 0.00222139f $X=0.432 $Y=0.2025 $X2=0 $Y2=0
cc_100 VSS N_Y_c_124_n 0.00222139f $X=0.54 $Y=0.2025 $X2=0 $Y2=0
cc_101 VSS N_Y_c_132_n 0.00169333f $X=0.54 $Y=0.2025 $X2=0 $Y2=0
cc_102 VSS N_Y_c_149_n 9.49966e-19 $X=0.54 $Y=0.234 $X2=0 $Y2=0
cc_103 VSS N_Y_c_115_n 3.96872e-19 $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_104 VSS N_Y_c_115_n 0.0143431f $X=0.236 $Y=0.234 $X2=0 $Y2=0
cc_105 VSS N_Y_c_104_n 0.00319086f $X=0.252 $Y=0.036 $X2=0.081 $Y2=0.135
cc_106 VSS N_Y_c_145_n 2.3841e-19 $X=0.288 $Y=0.036 $X2=0 $Y2=0
cc_107 VSS N_Y_c_121_n 2.3841e-19 $X=0.364 $Y=0.036 $X2=0 $Y2=0
cc_108 VSS N_Y_c_136_n 3.11971e-19 $X=0.432 $Y=0.036 $X2=0.081 $Y2=0.135
cc_109 VSS N_Y_c_113_n 0.00462434f $X=0.252 $Y=0.036 $X2=0 $Y2=0
cc_110 VSS N_Y_c_121_n 6.54052e-19 $X=0.419 $Y=0.09 $X2=0.405 $Y2=0.135
cc_111 VSS N_Y_c_124_n 6.54052e-19 $X=0.526 $Y=0.09 $X2=0.405 $Y2=0.135
cc_112 VSS N_Y_c_132_n 0.00322402f $X=0.486 $Y=0.0675 $X2=0 $Y2=0
cc_113 VSS N_Y_c_132_n 0.00354269f $X=0.592 $Y=0.0675 $X2=0 $Y2=0
cc_114 VSS N_Y_c_132_n 0.00228824f $X=0.553 $Y=0.09 $X2=0 $Y2=0
cc_115 VSS N_Y_c_134_n 0.0044312f $X=0.592 $Y=0.0675 $X2=0 $Y2=0
cc_116 VSS N_Y_c_136_n 4.45555e-19 $X=0.486 $Y=0.0675 $X2=0 $Y2=0
cc_117 VSS N_Y_c_136_n 0.00268693f $X=0.592 $Y=0.0675 $X2=0 $Y2=0
cc_118 VSS N_Y_c_136_n 0.00364017f $X=0.553 $Y=0.09 $X2=0 $Y2=0

* END of "./AOI31xp67_ASAP7_75t_L.pex.sp.AOI31XP67_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI321xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:14:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI321xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI321xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI321xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:14:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI321XP33_ASAP7_75T_L%A3 2 5 7 19 VSS
c5 19 VSS 0.0184885f $X=0.08 $Y=0.136
c6 5 VSS 0.00275452f $X=0.081 $Y=0.135
c7 2 VSS 0.0643308f $X=0.081 $Y=0.0675
r8 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r9 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r10 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI321XP33_ASAP7_75T_L%A2 2 5 7 17 VSS
c11 17 VSS 0.00290906f $X=0.134 $Y=0.136
c12 5 VSS 0.00132829f $X=0.135 $Y=0.135
c13 2 VSS 0.0599065f $X=0.135 $Y=0.0675
r14 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI321XP33_ASAP7_75T_L%A1 2 5 7 13 VSS
c12 13 VSS 0.00103414f $X=0.196 $Y=0.136
c13 5 VSS 0.00119626f $X=0.189 $Y=0.135
c14 2 VSS 0.0606095f $X=0.189 $Y=0.0675
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI321XP33_ASAP7_75T_L%C 2 5 7 10 VSS
c11 10 VSS 0.00128201f $X=0.243 $Y=0.134
c12 5 VSS 0.00120688f $X=0.243 $Y=0.135
c13 2 VSS 0.0616439f $X=0.243 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI321XP33_ASAP7_75T_L%B1 2 5 7 10 VSS
c11 10 VSS 9.49292e-19 $X=0.296 $Y=0.134
c12 5 VSS 0.00113128f $X=0.297 $Y=0.135
c13 2 VSS 0.0619909f $X=0.297 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AOI321XP33_ASAP7_75T_L%B2 2 5 7 10 VSS
c11 10 VSS 5.93188e-19 $X=0.348 $Y=0.134
c12 5 VSS 0.00170643f $X=0.351 $Y=0.135
c13 2 VSS 0.066866f $X=0.351 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.054 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AOI321XP33_ASAP7_75T_L%Y 2 3 5 8 15 16 19 23 26 27 32 35 38 40 45 46
+ 50 VSS
c27 50 VSS 0.00423691f $X=0.405 $Y=0.164
c28 49 VSS 0.00112176f $X=0.405 $Y=0.07
c29 48 VSS 0.00112176f $X=0.405 $Y=0.189
c30 46 VSS 8.46035e-21 $X=0.36 $Y=0.198
c31 45 VSS 4.59335e-19 $X=0.342 $Y=0.198
c32 40 VSS 0.00240073f $X=0.396 $Y=0.198
c33 39 VSS 8.90106e-19 $X=0.369 $Y=0.036
c34 38 VSS 0.00142296f $X=0.36 $Y=0.036
c35 37 VSS 0.00310342f $X=0.342 $Y=0.036
c36 36 VSS 4.3113e-19 $X=0.31 $Y=0.036
c37 35 VSS 0.00146362f $X=0.306 $Y=0.036
c38 34 VSS 0.00554947f $X=0.288 $Y=0.036
c39 33 VSS 4.31197e-19 $X=0.256 $Y=0.036
c40 32 VSS 0.00142296f $X=0.252 $Y=0.036
c41 28 VSS 4.19362e-19 $X=0.234 $Y=0.036
c42 27 VSS 0.00376122f $X=0.23 $Y=0.036
c43 23 VSS 0.00474306f $X=0.216 $Y=0.036
c44 20 VSS 0.00614869f $X=0.396 $Y=0.036
c45 19 VSS 0.00233317f $X=0.324 $Y=0.2025
c46 15 VSS 5.75997e-19 $X=0.341 $Y=0.2025
c47 8 VSS 0.00345731f $X=0.376 $Y=0.054
c48 4 VSS 5.22702e-19 $X=0.216 $Y=0.0455
r49 49 50 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.07 $X2=0.405 $Y2=0.164
r50 48 50 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.164
r51 47 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.07
r52 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r53 42 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.342 $Y2=0.198
r54 40 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.198 $X2=0.405 $Y2=0.189
r55 40 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.36 $Y2=0.198
r56 38 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.369 $Y2=0.036
r57 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r58 36 37 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.31
+ $Y=0.036 $X2=0.342 $Y2=0.036
r59 35 36 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.31 $Y2=0.036
r60 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r61 33 34 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.036 $X2=0.288 $Y2=0.036
r62 32 33 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.256 $Y2=0.036
r63 30 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.369 $Y2=0.036
r64 27 28 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.036 $X2=0.234 $Y2=0.036
r65 26 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.036 $X2=0.252 $Y2=0.036
r66 26 28 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.036 $X2=0.234 $Y2=0.036
r67 22 27 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.23 $Y2=0.036
r68 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r69 20 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r70 20 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.378 $Y2=0.036
r71 19 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198 $X2=0.324
+ $Y2=0.198
r72 16 19 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r73 15 19 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r74 14 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r75 8 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r76 5 8 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.054 $X2=0.376 $Y2=0.054
r77 3 4 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0455 $X2=0.216 $Y2=0.0455
r78 2 4 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0455 $X2=0.216 $Y2=0.0455
r79 1 14 3.12934 $w=6.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.216 $Y=0.064 $X2=0.199 $Y2=0.064
r80 1 4 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.216 $Y=0.064 $X2=0.216 $Y2=0.0455
.ends


* END of "./AOI321xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI321xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 C B1 B2 Y
* 
* Y	Y
* B2	B2
* B1	B1
* C	C
* A1	A1
* A2	A2
* A3	A3
M0 noxref_12 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_13 N_A2_M1_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_A1_M2_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_C_M3_g N_Y_M3_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 noxref_14 N_B1_M4_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.027
M5 N_Y_M5_d N_B2_M5_g noxref_14 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341
+ $Y=0.027
M6 noxref_9 N_A3_M6_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 VDD N_A2_M7_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 noxref_9 N_A1_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 noxref_10 N_C_M9_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 N_Y_M10_d N_B1_M10_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M11 noxref_10 N_B2_M11_g N_Y_M11_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
*
* 
* .include "AOI321xp33_ASAP7_75t_L.pex.sp.AOI321XP33_ASAP7_75T_L.pxi"
* BEGIN of "./AOI321xp33_ASAP7_75t_L.pex.sp.AOI321XP33_ASAP7_75T_L.pxi"
* File: AOI321xp33_ASAP7_75t_L.pex.sp.AOI321XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:14:48 2017
* 
x_PM_AOI321XP33_ASAP7_75T_L%A3 N_A3_M0_g N_A3_c_2_p N_A3_M6_g A3 VSS
+ PM_AOI321XP33_ASAP7_75T_L%A3
x_PM_AOI321XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_7_n N_A2_M7_g A2 VSS
+ PM_AOI321XP33_ASAP7_75T_L%A2
x_PM_AOI321XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_19_n N_A1_M8_g A1 VSS
+ PM_AOI321XP33_ASAP7_75T_L%A1
x_PM_AOI321XP33_ASAP7_75T_L%C N_C_M3_g N_C_c_31_n N_C_M9_g C VSS
+ PM_AOI321XP33_ASAP7_75T_L%C
x_PM_AOI321XP33_ASAP7_75T_L%B1 N_B1_M4_g N_B1_c_42_n N_B1_M10_g B1 VSS
+ PM_AOI321XP33_ASAP7_75T_L%B1
x_PM_AOI321XP33_ASAP7_75T_L%B2 N_B2_M5_g N_B2_c_53_n N_B2_M11_g B2 VSS
+ PM_AOI321XP33_ASAP7_75T_L%B2
x_PM_AOI321XP33_ASAP7_75T_L%Y N_Y_M3_s N_Y_M2_d N_Y_M5_d N_Y_c_71_n N_Y_M11_s
+ N_Y_M10_d N_Y_c_81_n N_Y_c_62_n Y N_Y_c_63_n N_Y_c_67_n N_Y_c_69_n N_Y_c_72_n
+ N_Y_c_84_n N_Y_c_79_n N_Y_c_74_n N_Y_c_76_n VSS PM_AOI321XP33_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_A2_M1_g 0.00347357f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A3_c_2_p N_A2_c_7_n 0.00120426f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A3 A2 0.00247926f $X=0.08 $Y=0.136 $X2=0.134 $Y2=0.136
cc_4 N_A3_M0_g N_A1_M2_g 2.69148e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 VSS A3 3.43147e-19 $X=0.08 $Y=0.136 $X2=0 $Y2=0
cc_6 N_A2_M1_g N_A1_M2_g 0.00325575f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_7 N_A2_c_7_n N_A1_c_19_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_8 A2 A1 0.00464813f $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_9 N_A2_M1_g N_C_M3_g 2.69148e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_10 VSS N_A2_M1_g 3.62029e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_11 VSS A2 0.0012376f $X=0.134 $Y=0.136 $X2=0.081 $Y2=0.135
cc_12 A2 N_Y_c_62_n 6.88222e-19 $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_13 A2 N_Y_c_63_n 4.76861e-19 $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_14 N_A1_M2_g N_C_M3_g 0.00359705f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_15 N_A1_c_19_n N_C_c_31_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_16 A1 C 0.00406615f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_17 N_A1_M2_g N_B1_M4_g 2.69148e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_18 VSS N_A1_M2_g 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_19 VSS A1 0.0012322f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_20 A1 N_Y_c_62_n 0.0013295f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_21 N_A1_M2_g N_Y_c_63_n 2.84579e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_22 N_C_M3_g N_B1_M4_g 0.00330657f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.0675
cc_23 N_C_c_31_n N_B1_c_42_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_24 C B1 0.00453023f $X=0.243 $Y=0.134 $X2=0.135 $Y2=0.135
cc_25 N_C_M3_g N_B2_M5_g 2.74891e-19 $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.0675
cc_26 C N_Y_c_62_n 0.00127618f $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_27 N_C_M3_g N_Y_c_67_n 2.56935e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_28 C N_Y_c_67_n 0.00123064f $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_29 N_B1_M4_g N_B2_M5_g 0.00372052f $X=0.297 $Y=0.054 $X2=0.189 $Y2=0.0675
cc_30 N_B1_c_42_n N_B2_c_53_n 9.33263e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_31 B1 B2 0.00484406f $X=0.296 $Y=0.134 $X2=0.189 $Y2=0.135
cc_32 VSS N_B1_M4_g 3.57119e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_33 VSS B1 5.37372e-19 $X=0.296 $Y=0.134 $X2=0 $Y2=0
cc_34 N_B1_M4_g N_Y_c_69_n 2.64276e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_35 B1 N_Y_c_69_n 0.00124805f $X=0.296 $Y=0.134 $X2=0 $Y2=0
cc_36 VSS N_B2_M5_g 2.08515e-19 $X=0.351 $Y=0.054 $X2=0 $Y2=0
cc_37 B2 N_Y_c_71_n 3.87865e-19 $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_38 N_B2_M5_g N_Y_c_72_n 2.56935e-19 $X=0.351 $Y=0.054 $X2=0 $Y2=0
cc_39 B2 N_Y_c_72_n 0.00123064f $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_40 N_B2_M5_g N_Y_c_74_n 2.76185e-19 $X=0.351 $Y=0.054 $X2=0 $Y2=0
cc_41 B2 N_Y_c_74_n 0.0012322f $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_42 B2 N_Y_c_76_n 0.00441847f $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_43 VSS N_Y_c_62_n 0.00138157f $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_44 VSS N_Y_c_63_n 2.10682e-19 $X=0.216 $Y=0.198 $X2=0 $Y2=0
cc_45 VSS N_Y_c_79_n 2.88175e-19 $X=0.216 $Y=0.198 $X2=0 $Y2=0
cc_46 VSS N_Y_c_71_n 9.98826e-19 $X=0.376 $Y=0.2025 $X2=0 $Y2=0
cc_47 VSS N_Y_c_81_n 0.0033367f $X=0.27 $Y=0.2025 $X2=0 $Y2=0
cc_48 VSS N_Y_c_81_n 0.00371671f $X=0.376 $Y=0.2025 $X2=0 $Y2=0
cc_49 VSS N_Y_c_81_n 0.00250965f $X=0.344 $Y=0.234 $X2=0 $Y2=0
cc_50 VSS N_Y_c_84_n 0.00284922f $X=0.376 $Y=0.2025 $X2=0 $Y2=0
cc_51 VSS N_Y_c_79_n 4.49388e-19 $X=0.27 $Y=0.2025 $X2=0 $Y2=0
cc_52 VSS N_Y_c_79_n 0.00369159f $X=0.344 $Y=0.234 $X2=0 $Y2=0
cc_53 VSS N_Y_c_74_n 0.00369159f $X=0.378 $Y=0.234 $X2=0 $Y2=0
cc_54 VSS N_Y_c_76_n 3.97918e-19 $X=0.376 $Y=0.2025 $X2=0 $Y2=0

* END of "./AOI321xp33_ASAP7_75t_L.pex.sp.AOI321XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI322xp5_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:15:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI322xp5_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI322xp5_ASAP7_75t_L.pex.sp.pex"
* File: AOI322xp5_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:15:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI322XP5_ASAP7_75T_L%B2 2 5 7 10 VSS
c8 10 VSS 0.00502923f $X=0.075 $Y=0.134
c9 5 VSS 0.00230059f $X=0.081 $Y=0.135
c10 2 VSS 0.0649001f $X=0.081 $Y=0.054
r11 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r12 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r13 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI322XP5_ASAP7_75T_L%B1 2 5 7 10 VSS
c10 10 VSS 0.00111927f $X=0.131 $Y=0.134
c11 5 VSS 0.00123757f $X=0.135 $Y=0.135
c12 2 VSS 0.0618615f $X=0.135 $Y=0.054
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI322XP5_ASAP7_75T_L%A1 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.187 $Y=0.136
c14 5 VSS 0.00111823f $X=0.189 $Y=0.135
c15 2 VSS 0.0618966f $X=0.189 $Y=0.0675
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI322XP5_ASAP7_75T_L%A2 2 5 7 13 VSS
c13 13 VSS 4.81053e-19 $X=0.247 $Y=0.136
c14 5 VSS 0.00112315f $X=0.243 $Y=0.135
c15 2 VSS 0.0623167f $X=0.243 $Y=0.0675
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI322XP5_ASAP7_75T_L%A3 2 5 7 13 VSS
c12 13 VSS 7.62261e-19 $X=0.296 $Y=0.136
c13 5 VSS 0.00110907f $X=0.297 $Y=0.135
c14 2 VSS 0.0620895f $X=0.297 $Y=0.0675
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AOI322XP5_ASAP7_75T_L%C2 2 5 7 10 VSS
c11 10 VSS 0.00116759f $X=0.348 $Y=0.134
c12 5 VSS 0.00113128f $X=0.351 $Y=0.135
c13 2 VSS 0.0624109f $X=0.351 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.054 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AOI322XP5_ASAP7_75T_L%C1 2 5 7 10 VSS
c11 10 VSS 5.93188e-19 $X=0.405 $Y=0.134
c12 5 VSS 0.00170643f $X=0.405 $Y=0.135
c13 2 VSS 0.066866f $X=0.405 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.054 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AOI322XP5_ASAP7_75T_L%Y 2 3 5 8 15 16 19 23 26 27 28 29 30 34 35 37
+ 39 42 44 49 50 54 VSS
c34 56 VSS 5.02308e-19 $X=0.459 $Y=0.177
c35 54 VSS 0.00418428f $X=0.459 $Y=0.164
c36 53 VSS 0.00112176f $X=0.459 $Y=0.07
c37 52 VSS 5.81969e-19 $X=0.459 $Y=0.189
c38 50 VSS 8.46035e-21 $X=0.414 $Y=0.198
c39 49 VSS 4.59335e-19 $X=0.396 $Y=0.198
c40 44 VSS 0.00240073f $X=0.45 $Y=0.198
c41 43 VSS 8.90106e-19 $X=0.423 $Y=0.036
c42 42 VSS 0.00142296f $X=0.414 $Y=0.036
c43 41 VSS 0.00310342f $X=0.396 $Y=0.036
c44 40 VSS 4.17449e-19 $X=0.364 $Y=0.036
c45 39 VSS 0.00146362f $X=0.36 $Y=0.036
c46 38 VSS 0.00666605f $X=0.342 $Y=0.036
c47 37 VSS 0.00146362f $X=0.306 $Y=0.036
c48 36 VSS 4.17449e-19 $X=0.288 $Y=0.036
c49 35 VSS 0.00307159f $X=0.284 $Y=0.036
c50 34 VSS 8.53778e-19 $X=0.252 $Y=0.036
c51 30 VSS 7.04757e-19 $X=0.241 $Y=0.036
c52 29 VSS 0.00340162f $X=0.234 $Y=0.036
c53 28 VSS 0.00146362f $X=0.198 $Y=0.036
c54 27 VSS 0.0039381f $X=0.18 $Y=0.036
c55 23 VSS 0.00305925f $X=0.162 $Y=0.036
c56 20 VSS 0.00615748f $X=0.45 $Y=0.036
c57 19 VSS 0.00234286f $X=0.378 $Y=0.2025
c58 15 VSS 5.75997e-19 $X=0.395 $Y=0.2025
c59 8 VSS 0.00345731f $X=0.43 $Y=0.054
c60 4 VSS 5.57323e-19 $X=0.162 $Y=0.0455
r61 55 56 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.177
r62 54 55 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.164 $X2=0.459 $Y2=0.165
r63 53 54 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.07 $X2=0.459 $Y2=0.164
r64 52 56 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.189 $X2=0.459 $Y2=0.177
r65 51 53 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.07
r66 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.414 $Y2=0.198
r67 46 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.198 $X2=0.396 $Y2=0.198
r68 44 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.198 $X2=0.459 $Y2=0.189
r69 44 50 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.198 $X2=0.414 $Y2=0.198
r70 42 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.423 $Y2=0.036
r71 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r72 40 41 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.364
+ $Y=0.036 $X2=0.396 $Y2=0.036
r73 39 40 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.364 $Y2=0.036
r74 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r75 37 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.342 $Y2=0.036
r76 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r77 35 36 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.036 $X2=0.288 $Y2=0.036
r78 34 35 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.284 $Y2=0.036
r79 32 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.423 $Y2=0.036
r80 29 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.241 $Y2=0.036
r81 28 29 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.234 $Y2=0.036
r82 27 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r83 26 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.036 $X2=0.252 $Y2=0.036
r84 26 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.036 $X2=0.241 $Y2=0.036
r85 22 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r86 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r87 20 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r88 20 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.432 $Y2=0.036
r89 19 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.198 $X2=0.378
+ $Y2=0.198
r90 16 19 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r91 15 19 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r92 14 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r93 8 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r94 5 8 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.054 $X2=0.43 $Y2=0.054
r95 3 4 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.0455 $X2=0.162 $Y2=0.0455
r96 2 4 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0455 $X2=0.162 $Y2=0.0455
r97 1 14 3.12934 $w=6.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.162 $Y=0.064 $X2=0.145 $Y2=0.064
r98 1 4 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.162 $Y=0.064 $X2=0.162 $Y2=0.0455
.ends


* END of "./AOI322xp5_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI322xp5_ASAP7_75t_L  VSS VDD B2 B1 A1 A2 A3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
M0 noxref_13 N_B2_M0_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_Y_M1_d N_B1_M1_g noxref_13 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 noxref_14 N_A1_M2_g N_Y_M2_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_15 N_A2_M3_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 VSS N_A3_M4_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_16 N_C2_M5_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341
+ $Y=0.027
M6 N_Y_M6_d N_C1_M6_g noxref_16 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.395
+ $Y=0.027
M7 VDD N_B2_M7_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M8 noxref_10 N_B1_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M9 noxref_11 N_A1_M9_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M10 noxref_10 N_A2_M10_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M11 noxref_11 N_A3_M11_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M12 N_Y_M12_d N_C2_M12_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M13 noxref_11 N_C1_M13_g N_Y_M13_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
*
* 
* .include "AOI322xp5_ASAP7_75t_L.pex.sp.AOI322XP5_ASAP7_75T_L.pxi"
* BEGIN of "./AOI322xp5_ASAP7_75t_L.pex.sp.AOI322XP5_ASAP7_75T_L.pxi"
* File: AOI322xp5_ASAP7_75t_L.pex.sp.AOI322XP5_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:15:10 2017
* 
x_PM_AOI322XP5_ASAP7_75T_L%B2 N_B2_M0_g N_B2_c_2_p N_B2_M7_g B2 VSS
+ PM_AOI322XP5_ASAP7_75T_L%B2
x_PM_AOI322XP5_ASAP7_75T_L%B1 N_B1_M1_g N_B1_c_10_n N_B1_M8_g B1 VSS
+ PM_AOI322XP5_ASAP7_75T_L%B1
x_PM_AOI322XP5_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_21_n N_A1_M9_g A1 VSS
+ PM_AOI322XP5_ASAP7_75T_L%A1
x_PM_AOI322XP5_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_34_n N_A2_M10_g A2 VSS
+ PM_AOI322XP5_ASAP7_75T_L%A2
x_PM_AOI322XP5_ASAP7_75T_L%A3 N_A3_M4_g N_A3_c_47_n N_A3_M11_g A3 VSS
+ PM_AOI322XP5_ASAP7_75T_L%A3
x_PM_AOI322XP5_ASAP7_75T_L%C2 N_C2_M5_g N_C2_c_59_n N_C2_M12_g C2 VSS
+ PM_AOI322XP5_ASAP7_75T_L%C2
x_PM_AOI322XP5_ASAP7_75T_L%C1 N_C1_M6_g N_C1_c_70_n N_C1_M13_g C1 VSS
+ PM_AOI322XP5_ASAP7_75T_L%C1
x_PM_AOI322XP5_ASAP7_75T_L%Y N_Y_M2_s N_Y_M1_d N_Y_M6_d N_Y_c_91_n N_Y_M13_s
+ N_Y_M12_d N_Y_c_103_n N_Y_c_79_n Y N_Y_c_80_n N_Y_c_83_n N_Y_c_99_n N_Y_c_85_n
+ N_Y_c_86_n N_Y_c_100_n N_Y_c_87_n N_Y_c_89_n N_Y_c_92_n N_Y_c_106_n
+ N_Y_c_101_n N_Y_c_94_n N_Y_c_96_n VSS PM_AOI322XP5_ASAP7_75T_L%Y
cc_1 N_B2_M0_g N_B1_M1_g 0.00323392f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_B2_c_2_p N_B1_c_10_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 B2 B1 0.00464555f $X=0.075 $Y=0.134 $X2=0.131 $Y2=0.134
cc_4 N_B2_M0_g N_A1_M2_g 2.69148e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 VSS N_B2_M0_g 3.62029e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_6 VSS B2 0.0012376f $X=0.075 $Y=0.134 $X2=0 $Y2=0
cc_7 B2 N_Y_c_79_n 4.85822e-19 $X=0.075 $Y=0.134 $X2=0 $Y2=0
cc_8 B2 N_Y_c_80_n 4.5241e-19 $X=0.075 $Y=0.134 $X2=0 $Y2=0
cc_9 N_B1_M1_g N_A1_M2_g 0.0036697f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_10 N_B1_c_10_n N_A1_c_21_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_11 B1 A1 0.00406615f $X=0.131 $Y=0.134 $X2=0.075 $Y2=0.134
cc_12 N_B1_M1_g N_A2_M3_g 3.09654e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_13 VSS N_B1_M1_g 3.62029e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_14 VSS B1 0.0012322f $X=0.131 $Y=0.134 $X2=0 $Y2=0
cc_15 B1 N_Y_c_79_n 0.00133251f $X=0.131 $Y=0.134 $X2=0 $Y2=0
cc_16 N_A1_M2_g N_A2_M3_g 0.00374235f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_17 N_A1_c_21_n N_A2_c_34_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_18 A1 A2 0.00483372f $X=0.187 $Y=0.136 $X2=0.081 $Y2=0.135
cc_19 N_A1_M2_g N_A3_M4_g 3.09654e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_20 VSS N_A1_M2_g 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_21 VSS A1 0.0012322f $X=0.187 $Y=0.136 $X2=0 $Y2=0
cc_22 A1 N_Y_c_79_n 0.0013295f $X=0.187 $Y=0.136 $X2=0 $Y2=0
cc_23 N_A1_M2_g N_Y_c_83_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 A1 N_Y_c_83_n 0.00124805f $X=0.187 $Y=0.136 $X2=0 $Y2=0
cc_25 N_A2_M3_g N_A3_M4_g 0.00372052f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_26 N_A2_c_34_n N_A3_c_47_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_27 A2 A3 0.00481174f $X=0.247 $Y=0.136 $X2=0.135 $Y2=0.135
cc_28 N_A2_M3_g N_C2_M5_g 2.74891e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_29 VSS N_A2_M3_g 2.68514e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_30 VSS A2 0.00121543f $X=0.247 $Y=0.136 $X2=0 $Y2=0
cc_31 VSS N_A2_M3_g 2.38303e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_32 A2 N_Y_c_85_n 0.00123064f $X=0.247 $Y=0.136 $X2=0 $Y2=0
cc_33 N_A2_M3_g N_Y_c_86_n 2.03357e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_34 N_A3_M4_g N_C2_M5_g 0.00335739f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_35 N_A3_c_47_n N_C2_c_59_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_36 A3 C2 0.00407881f $X=0.296 $Y=0.136 $X2=0.187 $Y2=0.136
cc_37 N_A3_M4_g N_C1_M6_g 2.74891e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_38 VSS N_A3_M4_g 3.45454e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_39 VSS A3 5.39731e-19 $X=0.296 $Y=0.136 $X2=0 $Y2=0
cc_40 N_A3_M4_g N_Y_c_87_n 2.64276e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_41 A3 N_Y_c_87_n 0.00124825f $X=0.296 $Y=0.136 $X2=0 $Y2=0
cc_42 N_C2_M5_g N_C1_M6_g 0.00372052f $X=0.351 $Y=0.054 $X2=0.243 $Y2=0.0675
cc_43 N_C2_c_59_n N_C1_c_70_n 9.33263e-19 $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_44 C2 C1 0.00479746f $X=0.348 $Y=0.134 $X2=0.243 $Y2=0.135
cc_45 VSS N_C2_M5_g 3.55324e-19 $X=0.351 $Y=0.054 $X2=0 $Y2=0
cc_46 VSS C2 5.47169e-19 $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_47 N_C2_M5_g N_Y_c_89_n 2.64276e-19 $X=0.351 $Y=0.054 $X2=0 $Y2=0
cc_48 C2 N_Y_c_89_n 0.00124825f $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_49 VSS N_C1_M6_g 2.08515e-19 $X=0.405 $Y=0.054 $X2=0 $Y2=0
cc_50 C1 N_Y_c_91_n 3.87865e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_51 N_C1_M6_g N_Y_c_92_n 2.56935e-19 $X=0.405 $Y=0.054 $X2=0 $Y2=0
cc_52 C1 N_Y_c_92_n 0.00123064f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_53 N_C1_M6_g N_Y_c_94_n 2.76185e-19 $X=0.405 $Y=0.054 $X2=0 $Y2=0
cc_54 C1 N_Y_c_94_n 0.0012322f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_55 C1 N_Y_c_96_n 0.00441564f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_56 VSS N_Y_c_79_n 0.00138157f $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_57 VSS N_Y_c_80_n 2.83966e-19 $X=0.1545 $Y=0.198 $X2=0 $Y2=0
cc_58 VSS N_Y_c_99_n 2.83966e-19 $X=0.202 $Y=0.198 $X2=0 $Y2=0
cc_59 VSS N_Y_c_100_n 2.83966e-19 $X=0.261 $Y=0.198 $X2=0 $Y2=0
cc_60 VSS N_Y_c_101_n 2.91395e-19 $X=0.27 $Y=0.198 $X2=0 $Y2=0
cc_61 VSS N_Y_c_91_n 9.98826e-19 $X=0.43 $Y=0.2025 $X2=0 $Y2=0
cc_62 VSS N_Y_c_103_n 0.00334511f $X=0.324 $Y=0.2025 $X2=0 $Y2=0
cc_63 VSS N_Y_c_103_n 0.00373054f $X=0.43 $Y=0.2025 $X2=0 $Y2=0
cc_64 VSS N_Y_c_103_n 0.00250965f $X=0.398 $Y=0.234 $X2=0 $Y2=0
cc_65 VSS N_Y_c_106_n 0.00284922f $X=0.43 $Y=0.2025 $X2=0 $Y2=0
cc_66 VSS N_Y_c_101_n 4.49388e-19 $X=0.324 $Y=0.2025 $X2=0 $Y2=0
cc_67 VSS N_Y_c_101_n 0.00369159f $X=0.398 $Y=0.234 $X2=0 $Y2=0
cc_68 VSS N_Y_c_94_n 0.00369159f $X=0.432 $Y=0.234 $X2=0 $Y2=0
cc_69 VSS N_Y_c_96_n 3.8442e-19 $X=0.43 $Y=0.2025 $X2=0 $Y2=0
cc_70 VSS N_Y_c_99_n 3.48201e-19 $X=0.234 $Y=0.036 $X2=0.081 $Y2=0.054
cc_71 VSS N_Y_c_100_n 3.19955e-19 $X=0.284 $Y=0.036 $X2=0.081 $Y2=0.054

* END of "./AOI322xp5_ASAP7_75t_L.pex.sp.AOI322XP5_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI32xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:15:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI32xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI32xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI32xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:15:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI32XP33_ASAP7_75T_L%A1 2 5 7 13 17 24 28 VSS
c12 30 VSS 4.23379e-19 $X=0.0315 $Y=0.234
c13 29 VSS 0.00314823f $X=0.027 $Y=0.234
c14 28 VSS 0.00378304f $X=0.036 $Y=0.2345
c15 24 VSS 0.00544585f $X=0.018 $Y=0.135
c16 20 VSS 3.39266e-19 $X=0.0565 $Y=0.135
c17 19 VSS 0.00110334f $X=0.049 $Y=0.135
c18 17 VSS 4.57556e-19 $X=0.064 $Y=0.135
c19 14 VSS 0.00105698f $X=0.018 $Y=0.207
c20 13 VSS 0.00255236f $X=0.018 $Y=0.189
c21 12 VSS 0.00110018f $X=0.018 $Y=0.225
c22 5 VSS 0.00503773f $X=0.081 $Y=0.135
c23 2 VSS 0.0656689f $X=0.081 $Y=0.0675
r24 29 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.0315 $Y2=0.234
r25 28 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.0315 $Y2=0.234
r26 25 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.234 $X2=0.027 $Y2=0.234
r27 19 20 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.049
+ $Y=0.135 $X2=0.0565 $Y2=0.135
r28 17 20 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.135 $X2=0.0565 $Y2=0.135
r29 17 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r30 15 24 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r31 15 19 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.049 $Y2=0.135
r32 13 14 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.207
r33 12 25 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.234
r34 12 14 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.207
r35 11 24 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r36 11 13 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.189
r37 5 18 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r38 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r39 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI32XP33_ASAP7_75T_L%A2 2 5 7 12 14 15 19 VSS
c21 19 VSS 5.21783e-19 $X=0.135 $Y=0.0785
c22 15 VSS 1.98685e-20 $X=0.135 $Y=0.1305
c23 14 VSS 2.62055e-19 $X=0.135 $Y=0.126
c24 12 VSS 0.00171912f $X=0.135 $Y=0.135
c25 5 VSS 0.00110641f $X=0.135 $Y=0.135
c26 2 VSS 0.0606055f $X=0.135 $Y=0.0675
r27 14 15 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.1305
r28 12 15 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.1305
r29 9 19 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.081 $X2=0.135 $Y2=0.072
r30 9 14 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.081 $X2=0.135 $Y2=0.126
r31 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r32 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r33 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI32XP33_ASAP7_75T_L%A3 2 5 7 11 15 17 18 VSS
c17 18 VSS 3.22517e-19 $X=0.201 $Y=0.189
c18 17 VSS 0.001236f $X=0.187 $Y=0.1945
c19 15 VSS 3.2206e-19 $X=0.189 $Y=0.1765
c20 11 VSS 5.70856e-19 $X=0.189 $Y=0.135
c21 5 VSS 0.00109247f $X=0.189 $Y=0.135
c22 2 VSS 0.0604511f $X=0.189 $Y=0.0675
r23 17 18 0.447408 $w=4.2e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.201
+ $Y=0.1945 $X2=0.201 $Y2=0.189
r24 15 18 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.1765 $X2=0.189 $Y2=0.189
r25 14 15 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.1765
r26 11 14 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.164
r27 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r28 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r29 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI32XP33_ASAP7_75T_L%B1 2 5 7 10 VSS
c11 10 VSS 9.97444e-19 $X=0.243 $Y=0.1195
c12 5 VSS 0.00113686f $X=0.243 $Y=0.135
c13 2 VSS 0.0617155f $X=0.243 $Y=0.054
r14 10 13 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.1195 $X2=0.243 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI32XP33_ASAP7_75T_L%B2 2 5 7 10 VSS
c11 10 VSS 4.87963e-19 $X=0.297 $Y=0.1335
c12 5 VSS 0.00170409f $X=0.297 $Y=0.135
c13 2 VSS 0.066446f $X=0.297 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AOI32XP33_ASAP7_75T_L%Y 1 6 9 11 12 15 18 19 26 29 30 31 34 37 43 44
+ 45 51 54 VSS
c27 52 VSS 7.16962e-19 $X=0.351 $Y=0.1765
c28 51 VSS 0.00417529f $X=0.351 $Y=0.164
c29 50 VSS 2.67033e-19 $X=0.351 $Y=0.07
c30 49 VSS 8.85605e-19 $X=0.351 $Y=0.063
c31 48 VSS 6.07272e-19 $X=0.351 $Y=0.189
c32 47 VSS 0.00338949f $X=0.351 $Y=0.045
c33 46 VSS 1.42799e-19 $X=0.34 $Y=0.198
c34 45 VSS 3.90732e-19 $X=0.338 $Y=0.198
c35 44 VSS 8.46035e-21 $X=0.306 $Y=0.198
c36 43 VSS 5.02599e-19 $X=0.288 $Y=0.198
c37 38 VSS 0.00199921f $X=0.342 $Y=0.198
c38 37 VSS 0.00146362f $X=0.306 $Y=0.036
c39 36 VSS 0.0030651f $X=0.288 $Y=0.036
c40 35 VSS 4.99302e-19 $X=0.256 $Y=0.036
c41 34 VSS 0.00142296f $X=0.252 $Y=0.036
c42 33 VSS 0.00242556f $X=0.234 $Y=0.036
c43 32 VSS 0.00455239f $X=0.222 $Y=0.036
c44 31 VSS 0.00146362f $X=0.198 $Y=0.036
c45 30 VSS 0.00339397f $X=0.18 $Y=0.036
c46 29 VSS 0.00340784f $X=0.144 $Y=0.036
c47 28 VSS 0.00111752f $X=0.104 $Y=0.036
c48 27 VSS 0.00162508f $X=0.094 $Y=0.036
c49 26 VSS 0.0023503f $X=0.078 $Y=0.036
c50 19 VSS 0.00338979f $X=0.054 $Y=0.036
c51 18 VSS 0.00236514f $X=0.054 $Y=0.036
c52 16 VSS 0.00365978f $X=0.342 $Y=0.036
c53 15 VSS 0.00220204f $X=0.27 $Y=0.216
c54 11 VSS 5.70405e-19 $X=0.287 $Y=0.216
c55 9 VSS 0.00345862f $X=0.322 $Y=0.054
c56 1 VSS 4.5957e-19 $X=0.071 $Y=0.0675
r57 51 52 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.164 $X2=0.351 $Y2=0.1765
r58 50 51 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.07 $X2=0.351 $Y2=0.164
r59 49 50 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.063 $X2=0.351 $Y2=0.07
r60 48 52 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.1765
r61 47 54 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.036
r62 47 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.063
r63 45 46 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.198 $X2=0.34 $Y2=0.198
r64 44 45 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.198 $X2=0.338 $Y2=0.198
r65 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.306 $Y2=0.198
r66 40 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.198 $X2=0.288 $Y2=0.198
r67 38 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.198 $X2=0.351 $Y2=0.189
r68 38 46 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.34 $Y2=0.198
r69 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r70 35 36 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.036 $X2=0.288 $Y2=0.036
r71 34 35 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.256 $Y2=0.036
r72 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r73 32 33 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.222
+ $Y=0.036 $X2=0.234 $Y2=0.036
r74 31 32 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.222 $Y2=0.036
r75 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r76 29 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.18 $Y2=0.036
r77 28 29 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.104
+ $Y=0.036 $X2=0.144 $Y2=0.036
r78 27 28 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.036 $X2=0.104 $Y2=0.036
r79 26 27 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.036 $X2=0.094 $Y2=0.036
r80 24 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.306 $Y2=0.036
r81 18 26 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.078 $Y2=0.036
r82 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r83 16 54 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.351 $Y2=0.036
r84 16 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.324 $Y2=0.036
r85 15 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.198 $X2=0.27
+ $Y2=0.198
r86 12 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.216 $X2=0.27 $Y2=0.216
r87 11 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.216 $X2=0.27 $Y2=0.216
r88 9 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r89 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.054 $X2=0.322 $Y2=0.054
r90 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r91 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./AOI32xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI32xp33_ASAP7_75t_L  VSS VDD A1 A2 A3 B1 B2 Y
* 
* Y	Y
* B2	B2
* B1	B1
* A3	A3
* A2	A2
* A1	A1
M0 noxref_10 N_A1_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_11 N_A2_M1_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_A3_M2_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_12 N_B1_M3_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_B2_M4_g noxref_12 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.027
M5 noxref_8 N_A1_M5_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M6 VDD N_A2_M6_g noxref_8 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M7 noxref_8 N_A3_M7_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M8 N_Y_M8_d N_B1_M8_g noxref_8 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M9 noxref_8 N_B2_M9_g N_Y_M9_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.189
*
* 
* .include "AOI32xp33_ASAP7_75t_L.pex.sp.AOI32XP33_ASAP7_75T_L.pxi"
* BEGIN of "./AOI32xp33_ASAP7_75t_L.pex.sp.AOI32XP33_ASAP7_75T_L.pxi"
* File: AOI32xp33_ASAP7_75t_L.pex.sp.AOI32XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:15:33 2017
* 
x_PM_AOI32XP33_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M5_g N_A1_c_3_p
+ N_A1_c_5_p N_A1_c_4_p A1 VSS PM_AOI32XP33_ASAP7_75T_L%A1
x_PM_AOI32XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_14_n N_A2_M6_g N_A2_c_15_n
+ N_A2_c_16_n N_A2_c_17_n A2 VSS PM_AOI32XP33_ASAP7_75T_L%A2
x_PM_AOI32XP33_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_36_n N_A3_M7_g N_A3_c_37_n
+ N_A3_c_38_n A3 N_A3_c_40_n VSS PM_AOI32XP33_ASAP7_75T_L%A3
x_PM_AOI32XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_53_n N_B1_M8_g B1 VSS
+ PM_AOI32XP33_ASAP7_75T_L%B1
x_PM_AOI32XP33_ASAP7_75T_L%B2 N_B2_M4_g N_B2_c_64_n N_B2_M9_g B2 VSS
+ PM_AOI32XP33_ASAP7_75T_L%B2
x_PM_AOI32XP33_ASAP7_75T_L%Y N_Y_M0_s N_Y_M4_d N_Y_c_86_n N_Y_M9_s N_Y_M8_d
+ N_Y_c_93_n N_Y_c_74_n N_Y_c_75_n N_Y_c_76_n N_Y_c_79_n N_Y_c_99_p N_Y_c_81_n
+ N_Y_c_84_n N_Y_c_87_n N_Y_c_83_n N_Y_c_89_n N_Y_c_98_n N_Y_c_91_n Y VSS
+ PM_AOI32XP33_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00354623f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_14_n 0.0010528f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p N_A2_c_15_n 8.09446e-19 $X=0.018 $Y=0.189 $X2=0.135 $Y2=0.135
cc_4 N_A1_c_4_p N_A2_c_16_n 5.60591e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.126
cc_5 N_A1_c_5_p N_A2_c_17_n 4.18081e-19 $X=0.064 $Y=0.135 $X2=0.135 $Y2=0.1305
cc_6 N_A1_c_4_p A2 4.92635e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.0785
cc_7 N_A1_M0_g N_A3_M2_g 2.69148e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_8 VSS A1 5.7877e-19 $X=0.036 $Y=0.2345 $X2=0 $Y2=0
cc_9 N_A1_c_4_p N_Y_M0_s 2.23359e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_10 N_A1_c_4_p N_Y_c_74_n 9.06393e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.072
cc_11 N_A1_c_4_p N_Y_c_75_n 0.00225778f $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.0785
cc_12 N_A1_c_2_p N_Y_c_76_n 3.06588e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_13 N_A2_M1_g N_A3_M2_g 0.00323392f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_A2_c_14_n N_A3_c_36_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 A2 N_A3_c_37_n 0.00161862f $X=0.135 $Y=0.0785 $X2=0.018 $Y2=0.144
cc_16 N_A2_c_16_n N_A3_c_38_n 0.00161862f $X=0.135 $Y=0.126 $X2=0.027 $Y2=0.135
cc_17 N_A2_c_15_n A3 0.00161862f $X=0.135 $Y=0.135 $X2=0.064 $Y2=0.135
cc_18 N_A2_c_15_n N_A3_c_40_n 0.00161862f $X=0.135 $Y=0.135 $X2=0.064 $Y2=0.135
cc_19 N_A2_M1_g N_B1_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_20 VSS N_A2_c_15_n 0.00215958f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 VSS N_A2_c_15_n 0.00401037f $X=0.135 $Y=0.135 $X2=0.064 $Y2=0.135
cc_22 VSS N_A2_M1_g 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0.018 $Y2=0.234
cc_23 N_A2_c_16_n N_Y_c_75_n 7.60168e-19 $X=0.135 $Y=0.126 $X2=0.049 $Y2=0.135
cc_24 A2 N_Y_c_75_n 6.40333e-19 $X=0.135 $Y=0.0785 $X2=0.049 $Y2=0.135
cc_25 N_A2_M1_g N_Y_c_79_n 3.27325e-19 $X=0.135 $Y=0.0675 $X2=0.027 $Y2=0.234
cc_26 A2 N_Y_c_79_n 0.00424732f $X=0.135 $Y=0.0785 $X2=0.027 $Y2=0.234
cc_27 VSS A2 3.27354e-19 $X=0.135 $Y=0.0785 $X2=0.081 $Y2=0.0675
cc_28 N_A3_M2_g N_B1_M3_g 0.00323392f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_29 N_A3_c_36_n N_B1_c_53_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_30 N_A3_c_37_n B1 0.00383317f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_31 N_A3_M2_g N_B2_M4_g 2.69148e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_32 VSS A3 0.00222856f $X=0.187 $Y=0.1945 $X2=0 $Y2=0
cc_33 VSS N_A3_M2_g 2.34993e-19 $X=0.189 $Y=0.0675 $X2=0.0315 $Y2=0.234
cc_34 VSS A3 0.00413281f $X=0.187 $Y=0.1945 $X2=0.0315 $Y2=0.234
cc_35 N_A3_M2_g N_Y_c_81_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_A3_c_37_n N_Y_c_81_n 0.00125427f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_37 A3 N_Y_c_83_n 7.98429e-19 $X=0.187 $Y=0.1945 $X2=0 $Y2=0
cc_38 N_B1_M3_g N_B2_M4_g 0.0036697f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.0675
cc_39 N_B1_c_53_n N_B2_c_64_n 9.33263e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_40 B1 B2 0.00487321f $X=0.243 $Y=0.1195 $X2=0 $Y2=0
cc_41 VSS N_B1_M3_g 3.47199e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_42 VSS B1 5.30079e-19 $X=0.243 $Y=0.1195 $X2=0 $Y2=0
cc_43 N_B1_M3_g N_Y_c_84_n 2.56935e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_44 B1 N_Y_c_84_n 0.00123064f $X=0.243 $Y=0.1195 $X2=0 $Y2=0
cc_45 VSS N_B2_M4_g 2.38303e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_46 B2 N_Y_c_86_n 3.87865e-19 $X=0.297 $Y=0.1335 $X2=0.189 $Y2=0.189
cc_47 N_B2_M4_g N_Y_c_87_n 2.64276e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_48 B2 N_Y_c_87_n 0.00124805f $X=0.297 $Y=0.1335 $X2=0 $Y2=0
cc_49 N_B2_M4_g N_Y_c_89_n 2.76185e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_50 B2 N_Y_c_89_n 0.0012322f $X=0.297 $Y=0.1335 $X2=0 $Y2=0
cc_51 B2 N_Y_c_91_n 0.00445407f $X=0.297 $Y=0.1335 $X2=0 $Y2=0
cc_52 VSS N_Y_c_86_n 4.54531e-19 $X=0.322 $Y=0.216 $X2=0 $Y2=0
cc_53 VSS N_Y_c_93_n 0.00288888f $X=0.216 $Y=0.216 $X2=0.027 $Y2=0.135
cc_54 VSS N_Y_c_93_n 0.00302498f $X=0.322 $Y=0.216 $X2=0.027 $Y2=0.135
cc_55 VSS N_Y_c_93_n 0.00250965f $X=0.324 $Y=0.234 $X2=0.027 $Y2=0.135
cc_56 VSS N_Y_c_83_n 2.56435e-19 $X=0.216 $Y=0.216 $X2=0 $Y2=0
cc_57 VSS N_Y_c_83_n 0.00705732f $X=0.324 $Y=0.234 $X2=0 $Y2=0
cc_58 VSS N_Y_c_98_n 0.00391824f $X=0.322 $Y=0.216 $X2=0 $Y2=0
cc_59 VSS N_Y_c_99_p 4.8755e-19 $X=0.18 $Y=0.036 $X2=0.081 $Y2=0.0675

* END of "./AOI32xp33_ASAP7_75t_L.pex.sp.AOI32XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI331xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:15:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI331xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI331xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI331xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:15:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
* File: AOI331xp33_ASAP7_75t_SL.pex.netlist.pex
* Created: Fri Sep  8 15:43:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI331xp33_ASAP7_75t_SL%A3 2 5 7 10 VSS
c11 10 VSS 0.00760948f
c12 5 VSS 0.00156103f
c13 2 VSS 0.0591573f
r14 10 13 1.35802
r15 5 13 6.07099 $a=3.24e-16
r16 5 7 252.889
r17 2 5 252.889
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%A2 2 5 7 10 VSS
c12 10 VSS 0.00281637f
c13 5 VSS 0.00105303f
c14 2 VSS 0.0597431f
r15 10 15 1.35802
r16 5 15 6.07099 $a=3.24e-16
r17 5 7 252.889
r18 2 5 252.889
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%A1 2 5 7 10 13 VSS
c13 13 VSS 0.00115482f
c14 10 VSS 9.20655e-19
c15 5 VSS 0.00120113f
c16 2 VSS 0.0607001f
r17 10 13 1.35802
r18 5 13 6.07099 $a=3.24e-16
r19 5 7 252.889
r20 2 5 252.889
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%B1 2 5 7 10 VSS
c13 10 VSS 5.11375e-19
c14 5 VSS 0.00110017f
c15 2 VSS 0.0616432f
r16 10 13 1.29012
r17 5 13 6.07099 $a=3.24e-16
r18 5 7 252.889
r19 2 5 252.889
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%B2 2 5 7 10 VSS
c13 10 VSS 4.81053e-19
c14 5 VSS 0.00112057f
c15 2 VSS 0.0616432f
r16 10 13 1.35802
r17 5 13 6.07099 $a=3.24e-16
r18 5 7 252.889
r19 2 5 252.889
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%B3 2 5 7 10 VSS
c11 10 VSS 6.93937e-19
c12 5 VSS 9.76227e-19
c13 2 VSS 0.0619588f
r14 10 13 1.35802
r15 5 13 6.07099 $a=3.24e-16
r16 5 7 252.889
r17 2 5 252.889
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%C1 2 5 7 10 VSS
c12 10 VSS 0.0022532f
c13 5 VSS 0.00126988f
c14 2 VSS 0.0618014f
r15 10 13 1.35802
r16 5 13 6.07099 $a=3.24e-16
r17 5 7 252.889
r18 2 5 252.889
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%net031 1 2 5 6 7 10 11 12 15 24 26 30 33 35
+ VSS
c22 35 VSS 0.00277595f
c23 33 VSS 0.00160383f
c24 32 VSS 0.00251354f
c25 30 VSS 0.00445081f
c26 28 VSS 8.81722e-19
c27 26 VSS 0.00164964f
c28 25 VSS 0.00672353f
c29 24 VSS 0.00146362f
c30 23 VSS 0.00474634f
c31 15 VSS 0.00240395f
c32 11 VSS 6.28007e-19
c33 10 VSS 0.00597448f
c34 6 VSS 5.25448e-19
c35 5 VSS 0.0102025f
c36 1 VSS 5.37876e-19
r37 33 35 2.51235
r38 32 33 1.22222
r39 30 35 2.37654
r40 26 28 0.712963
r41 25 26 1.22222
r42 24 25 2.44444
r43 23 24 1.22222
r44 21 32 1.22222
r45 21 28 0.509259
r46 17 23 1.22222
r47 15 30 6.07099 $a=3.24e-16
r48 12 15 8.39506
r49 11 15 8.39506
r50 10 21 6.07099 $a=3.24e-16
r51 7 10 8.39506
r52 6 10 8.39506
r53 5 17 6.07099 $a=3.24e-16
r54 2 5 8.39506
r55 1 5 8.39506
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%net030 1 2 5 6 7 10 16 18 19 20 22 23 VSS
c21 23 VSS 4.305e-19
c22 22 VSS 5.36594e-19
c23 20 VSS 4.85415e-19
c24 19 VSS 8.46035e-21
c25 18 VSS 4.82421e-19
c26 16 VSS 0.0014984f
c27 10 VSS 0.00249476f
c28 6 VSS 6.65915e-19
c29 5 VSS 0.00259461f
c30 1 VSS 5.77541e-19
r31 22 23 0.611111
r32 20 22 1.42593
r33 19 20 2.24074
r34 18 19 1.22222
r35 16 23 0.611111
r36 12 18 1.22222
r37 10 16 6.07099 $a=3.24e-16
r38 7 10 8.39506
r39 6 10 8.39506
r40 5 12 6.07099 $a=3.24e-16
r41 2 5 8.39506
r42 1 5 8.39506
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%Y 1 2 6 11 14 16 19 23 24 25 27 28 29 30 31
+ 33 39 40 41 43 44 50 51 VSS
c34 51 VSS 0.00385307f
c35 50 VSS 0.00286577f
c36 45 VSS 6.83364e-19
c37 44 VSS 4.05647e-19
c38 43 VSS 5.76058e-19
c39 41 VSS 6.56706e-19
c40 40 VSS 5.64537e-19
c41 39 VSS 0.00168412f
c42 35 VSS 7.50497e-19
c43 33 VSS 0.00167953f
c44 31 VSS 0.00627688f
c45 30 VSS 0.00142296f
c46 29 VSS 0.00343941f
c47 28 VSS 0.00142296f
c48 27 VSS 0.00326561f
c49 25 VSS 0.00167697f
c50 24 VSS 0.00428544f
c51 23 VSS 0.00676142f
c52 19 VSS 0.00218628f
c53 16 VSS 0.00562693f
c54 14 VSS 0.00259367f
c55 9 VSS 2.55988e-19
c56 1 VSS 5.61153e-19
r57 51 52 0.305556
r58 50 52 0.305556
r59 47 51 1.22222
r60 45 50 0.682891
r61 44 45 0.611111
r62 43 44 1.22222
r63 42 43 1.69753
r64 40 41 1.93519
r65 39 42 2.51235
r66 39 41 1.93519
r67 36 40 1.69753
r68 33 35 0.712963
r69 31 33 1.42593
r70 30 31 2.24074
r71 29 30 1.22222
r72 28 29 2.44444
r73 27 28 1.22222
r74 25 27 2.44444
r75 24 25 1.22222
r76 22 35 0.509259
r77 22 23 6.07099 $a=3.24e-16
r78 18 24 1.22222
r79 18 19 6.07099 $a=3.24e-16
r80 16 36 0.682891
r81 16 22 1.22222
r82 14 47 6.07099 $a=3.24e-16
r83 11 14 7.40741
r84 9 23 27.1875
r85 6 9 7.40741
r86 5 19 27.1875
r87 2 5 8.39506
r88 1 5 8.39506
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%net25 1 2 VSS
c0 1 VSS 0.00221026f
r1 1 2 16.7901
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%net26 1 2 VSS
c0 1 VSS 0.00221026f
r1 1 2 16.7901
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%net063 1 2 VSS
c1 1 VSS 0.00181886f
r2 1 2 16.7901
.ends

.subckt PM_AOI331xp33_ASAP7_75t_SL%net064 1 2 VSS
c1 1 VSS 0.00183233f
r2 1 2 16.7901
.ends


* END of "./AOI331xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI331xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C1 Y
* 
* Y	Y
* C1	C1
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
MM3 N_net25_MM3_d N_A3_MM3_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=0.071
+ $Y=0.027
MM2 N_net26_MM2_d N_A2_MM2_g N_net25_MM2_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
+ $X=0.125 $Y=0.027
MM14 N_Y_MM14_d N_A1_MM14_g N_net26_MM14_s VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
+ $X=0.179 $Y=0.027
MM12 N_Y_MM12_d N_B1_MM12_g N_net063_MM12_s VSS nmos_rvt L=2e-08 W=8.1e-08
+ nfin=3 $X=0.233 $Y=0.027
MM11 N_net063_MM11_d N_B2_MM11_g N_net064_MM11_s VSS nmos_rvt L=2e-08 W=8.1e-08
+ nfin=3 $X=0.287 $Y=0.027
MM10 N_net064_MM10_d N_B3_MM10_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3
+ $X=0.341 $Y=0.027
MM17 N_Y_MM17_d N_C1_MM17_g VSS VSS nmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=0.395
+ $Y=0.027
MM7 N_net031_MM7_d N_A3_MM7_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=0.071
+ $Y=0.162
MM8 N_net031_MM8_d N_A2_MM8_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=0.125
+ $Y=0.162
MM9 N_net031_MM9_d N_A1_MM9_g VDD VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3 $X=0.179
+ $Y=0.162
MM6 N_net030_MM6_d N_B1_MM6_g N_net031_MM6_s VDD pmos_rvt L=2e-08 W=8.1e-08
+ nfin=3 $X=0.233 $Y=0.162
MM5 N_net030_MM5_d N_B2_MM5_g N_net031_MM5_s VDD pmos_rvt L=2e-08 W=8.1e-08
+ nfin=3 $X=0.287 $Y=0.162
MM4 N_net030_MM4_d N_B3_MM4_g N_net031_MM4_s VDD pmos_rvt L=2e-08 W=8.1e-08
+ nfin=3 $X=0.341 $Y=0.162
MM1 N_Y_MM1_d N_C1_MM1_g N_net030_MM1_s VDD pmos_rvt L=2e-08 W=8.1e-08 nfin=3
+ $X=0.395 $Y=0.162
*
* 
* File: AOI331xp33_ASAP7_75t_SL.pex.netlist.AOI331xp33_ASAP7_75t_SL.pxi
* Created: Fri Sep  8 15:43:41 2017
* 
x_PM_AOI331xp33_ASAP7_75t_SL%A3 N_A3_MM3_g N_A3_c_2_p N_A3_MM7_g A3 vss!
+ PM_AOI331xp33_ASAP7_75t_SL%A3
x_PM_AOI331xp33_ASAP7_75t_SL%A2 N_A2_MM2_g N_A2_c_13_n N_A2_MM8_g A2 vss!
+ PM_AOI331xp33_ASAP7_75t_SL%A2
x_PM_AOI331xp33_ASAP7_75t_SL%A1 N_A1_MM14_g N_A1_c_26_n N_A1_MM9_g A1
+ N_A1_c_34_p vss! PM_AOI331xp33_ASAP7_75t_SL%A1
x_PM_AOI331xp33_ASAP7_75t_SL%B1 N_B1_MM12_g N_B1_c_39_n N_B1_MM6_g B1 vss!
+ PM_AOI331xp33_ASAP7_75t_SL%B1
x_PM_AOI331xp33_ASAP7_75t_SL%B2 N_B2_MM11_g N_B2_c_52_n N_B2_MM5_g B2 vss!
+ PM_AOI331xp33_ASAP7_75t_SL%B2
x_PM_AOI331xp33_ASAP7_75t_SL%B3 N_B3_MM10_g N_B3_c_65_n N_B3_MM4_g B3 vss!
+ PM_AOI331xp33_ASAP7_75t_SL%B3
x_PM_AOI331xp33_ASAP7_75t_SL%C1 N_C1_MM17_g N_C1_c_76_n N_C1_MM1_g C1 vss!
+ PM_AOI331xp33_ASAP7_75t_SL%C1
x_PM_AOI331xp33_ASAP7_75t_SL%net031 N_net031_MM8_d N_net031_MM7_d
+ N_net031_c_86_n N_net031_MM6_s N_net031_MM9_d N_net031_c_90_n N_net031_MM4_s
+ N_net031_MM5_s N_net031_c_97_p N_net031_c_88_n N_net031_c_91_n N_net031_c_95_n
+ N_net031_c_93_n N_net031_c_98_p vss! PM_AOI331xp33_ASAP7_75t_SL%net031
x_PM_AOI331xp33_ASAP7_75t_SL%net030 N_net030_MM5_d N_net030_MM6_d
+ N_net030_c_113_n N_net030_MM1_s N_net030_MM4_d N_net030_c_116_n
+ N_net030_c_123_p N_net030_c_108_n N_net030_c_109_n N_net030_c_121_n
+ N_net030_c_111_n N_net030_c_126_p vss! PM_AOI331xp33_ASAP7_75t_SL%net030
x_PM_AOI331xp33_ASAP7_75t_SL%Y N_Y_MM12_d N_Y_MM14_d N_Y_MM17_d N_Y_MM1_d
+ N_Y_c_143_n N_Y_c_155_p N_Y_c_129_n N_Y_c_139_n N_Y_c_130_n N_Y_c_133_n
+ N_Y_c_148_n N_Y_c_135_n N_Y_c_149_n N_Y_c_137_n N_Y_c_150_n N_Y_c_140_n Y
+ N_Y_c_157_p N_Y_c_142_n N_Y_c_160_p N_Y_c_151_n N_Y_c_162_p N_Y_c_145_n vss!
+ PM_AOI331xp33_ASAP7_75t_SL%Y
x_PM_AOI331xp33_ASAP7_75t_SL%net25 N_net25_MM2_s N_net25_MM3_d vss!
+ PM_AOI331xp33_ASAP7_75t_SL%net25
x_PM_AOI331xp33_ASAP7_75t_SL%net26 N_net26_MM14_s N_net26_MM2_d vss!
+ PM_AOI331xp33_ASAP7_75t_SL%net26
x_PM_AOI331xp33_ASAP7_75t_SL%net063 N_net063_MM11_d N_net063_MM12_s vss!
+ PM_AOI331xp33_ASAP7_75t_SL%net063
x_PM_AOI331xp33_ASAP7_75t_SL%net064 N_net064_MM10_d N_net064_MM11_s vss!
+ PM_AOI331xp33_ASAP7_75t_SL%net064
cc_1 N_A3_MM3_g N_A2_MM2_g 0.00344695f
cc_2 N_A3_c_2_p N_A2_c_13_n 9.33263e-19
cc_3 A3 A2 0.00752842f
cc_4 N_A3_MM3_g N_A1_MM14_g 2.66145e-19
cc_5 A3 N_net031_c_86_n 0.00114532f
cc_6 vss! N_A3_MM3_g 0.00149874f
cc_7 vss! N_A3_c_2_p 5.63328e-19
cc_8 vss! A3 2.01978e-19
cc_9 vss! N_A3_MM3_g 0.00149874f
cc_10 vss! N_A3_c_2_p 5.50525e-19
cc_11 vss! A3 2.01978e-19
cc_12 N_A2_MM2_g N_A1_MM14_g 0.00327995f
cc_13 N_A2_c_13_n N_A1_c_26_n 8.86777e-19
cc_14 A2 A1 0.00564665f
cc_15 N_A2_MM2_g N_B1_MM12_g 2.71887e-19
cc_16 A2 N_net031_c_86_n 0.00114532f
cc_17 N_A2_MM2_g N_net031_c_88_n 2.64276e-19
cc_18 A2 N_net031_c_88_n 0.00125674f
cc_19 A2 N_Y_c_129_n 5.87506e-19
cc_20 A2 N_Y_c_130_n 4.59602e-19
cc_21 N_A1_MM14_g N_B1_MM12_g 0.0036939f
cc_22 N_A1_c_26_n N_B1_c_39_n 8.86777e-19
cc_23 A1 B1 0.00389755f
cc_24 N_A1_MM14_g N_B2_MM11_g 3.06651e-19
cc_25 A1 N_net031_c_90_n 8.72546e-19
cc_26 N_A1_MM14_g N_net031_c_91_n 2.64276e-19
cc_27 N_A1_c_34_p N_net031_c_91_n 0.00125352f
cc_28 N_A1_c_34_p N_net030_c_108_n 2.75021e-19
cc_29 A1 N_Y_c_129_n 0.0013295f
cc_30 N_B1_MM12_g N_B2_MM11_g 0.00371573f
cc_31 N_B1_c_39_n N_B2_c_52_n 8.86777e-19
cc_32 B1 B2 0.00483372f
cc_33 N_B1_MM12_g N_B3_MM10_g 3.06651e-19
cc_34 N_B1_MM12_g N_net031_c_93_n 3.57119e-19
cc_35 B1 N_net031_c_93_n 5.37372e-19
cc_36 B1 N_Y_c_129_n 0.0013295f
cc_37 N_B1_MM12_g N_Y_c_133_n 2.64276e-19
cc_38 B1 N_Y_c_133_n 0.00124805f
cc_39 N_B2_MM11_g N_B3_MM10_g 0.0036939f
cc_40 N_B2_c_52_n N_B3_c_65_n 8.86777e-19
cc_41 B2 B3 0.00483372f
cc_42 N_B2_MM11_g N_C1_MM17_g 2.71887e-19
cc_43 N_B2_MM11_g N_net031_c_95_n 2.21754e-19
cc_44 N_B2_MM11_g N_net030_c_109_n 2.76185e-19
cc_45 B2 N_net030_c_109_n 0.0012322f
cc_46 N_B2_MM11_g N_Y_c_135_n 3.38929e-19
cc_47 B2 N_Y_c_135_n 0.00123064f
cc_48 N_B3_MM10_g N_C1_MM17_g 0.00333077f
cc_49 N_B3_c_65_n N_C1_c_76_n 9.33263e-19
cc_50 B3 C1 0.00406322f
cc_51 N_B3_MM10_g N_net030_c_111_n 3.51973e-19
cc_52 B3 N_net030_c_111_n 0.00121543f
cc_53 N_B3_MM10_g N_Y_c_137_n 2.56935e-19
cc_54 B3 N_Y_c_137_n 0.00123064f
cc_55 C1 N_Y_c_139_n 0.00114532f
cc_56 N_C1_MM17_g N_Y_c_140_n 2.64276e-19
cc_57 C1 N_Y_c_140_n 0.00124805f
cc_58 C1 N_Y_c_142_n 0.00391435f
cc_59 vss! N_C1_MM17_g 0.00188828f
cc_60 vss! N_C1_c_76_n 4.4617e-19
cc_61 vss! N_C1_MM17_g 0.00201175f
cc_62 vss! N_C1_c_76_n 4.3603e-19
cc_63 N_net031_c_90_n N_net030_c_113_n 0.00364173f
cc_64 N_net031_c_97_p N_net030_c_113_n 0.00355395f
cc_65 N_net031_c_98_p N_net030_c_113_n 0.00250965f
cc_66 N_net031_c_97_p N_net030_c_116_n 0.00323383f
cc_67 N_net031_c_95_n N_net030_c_116_n 4.54631e-19
cc_68 N_net031_c_90_n N_net030_c_108_n 3.69901e-19
cc_69 N_net031_c_98_p N_net030_c_108_n 0.00365081f
cc_70 N_net031_c_95_n N_net030_c_109_n 0.00365081f
cc_71 N_net031_c_97_p N_net030_c_121_n 0.00233206f
cc_72 N_net031_c_97_p N_Y_c_143_n 2.24644e-19
cc_73 N_net031_c_90_n N_Y_c_129_n 0.00107252f
cc_74 N_net031_c_95_n N_Y_c_145_n 2.83845e-19
cc_75 N_net030_c_116_n N_Y_c_143_n 0.0036142f
cc_76 N_net030_c_123_p N_Y_c_143_n 3.99913e-19
cc_77 N_net030_c_108_n N_Y_c_148_n 3.03225e-19
cc_78 N_net030_c_121_n N_Y_c_149_n 3.03225e-19
cc_79 N_net030_c_126_p N_Y_c_150_n 3.03225e-19
cc_80 N_net030_c_123_p N_Y_c_151_n 3.49487e-19
cc_81 N_net030_c_116_n N_Y_c_145_n 4.47506e-19
cc_82 N_Y_c_148_n N_net063_MM11_d 3.48201e-19
cc_83 N_Y_c_149_n N_net064_MM10_d 3.34078e-19
cc_84 vss! N_Y_c_155_p 3.1415e-19
cc_85 vss! Y 7.0789e-19
cc_86 vss! N_Y_c_157_p 2.46707e-19
cc_87 vss! N_Y_c_142_n 5.21182e-19
cc_88 vss! Y 5.58472e-19
cc_89 vss! N_Y_c_160_p 4.86009e-19
cc_90 vss! N_Y_c_151_n 2.60982e-19
cc_91 vss! N_Y_c_162_p 2.64997e-19

* END of "./AOI331xp33_ASAP7_75t_L.pex.sp.AOI331XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI332xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:16:17 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI332xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI332xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI332xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:16:17 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI332XP33_ASAP7_75T_L%A3 2 5 7 10 VSS
c4 10 VSS 0.00613146f $X=0.081 $Y=0.115
c5 5 VSS 0.00238289f $X=0.081 $Y=0.135
c6 2 VSS 0.062704f $X=0.081 $Y=0.0675
r7 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.115 $X2=0.081 $Y2=0.135
r8 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r9 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r10 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI332XP33_ASAP7_75T_L%A2 2 5 7 10 VSS
c11 10 VSS 0.00174706f $X=0.135 $Y=0.115
c12 5 VSS 0.00123757f $X=0.135 $Y=0.135
c13 2 VSS 0.0598541f $X=0.135 $Y=0.0675
r14 10 15 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.115 $X2=0.135 $Y2=0.135
r15 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI332XP33_ASAP7_75T_L%A1 2 5 7 10 VSS
c11 10 VSS 0.00101969f $X=0.189 $Y=0.115
c12 5 VSS 0.00121257f $X=0.189 $Y=0.135
c13 2 VSS 0.0608354f $X=0.189 $Y=0.0675
r14 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI332XP33_ASAP7_75T_L%B1 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.243 $Y=0.116
c14 5 VSS 0.00111336f $X=0.243 $Y=0.135
c15 2 VSS 0.0617786f $X=0.243 $Y=0.0675
r16 10 13 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.116 $X2=0.243 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI332XP33_ASAP7_75T_L%B2 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.296 $Y=0.115
c14 5 VSS 0.00112198f $X=0.297 $Y=0.135
c15 2 VSS 0.0616432f $X=0.297 $Y=0.0675
r16 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.115 $X2=0.297 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AOI332XP33_ASAP7_75T_L%B3 2 5 7 10 VSS
c12 10 VSS 7.27237e-19 $X=0.349 $Y=0.115
c13 5 VSS 0.00111185f $X=0.351 $Y=0.135
c14 2 VSS 0.0615515f $X=0.351 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.115 $X2=0.351 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AOI332XP33_ASAP7_75T_L%C2 2 5 7 10 VSS
c11 10 VSS 0.00167719f $X=0.406 $Y=0.114
c12 5 VSS 0.00113407f $X=0.405 $Y=0.135
c13 2 VSS 0.0618699f $X=0.405 $Y=0.0675
r14 10 13 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.114 $X2=0.405 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AOI332XP33_ASAP7_75T_L%C1 2 5 7 10 VSS
c11 10 VSS 4.90626e-19 $X=0.459 $Y=0.115
c12 5 VSS 0.00170409f $X=0.459 $Y=0.135
c13 2 VSS 0.0662985f $X=0.459 $Y=0.0675
r14 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.115 $X2=0.459 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AOI332XP33_ASAP7_75T_L%Y 1 2 6 11 12 15 19 23 24 25 26 27 28 30 32 34
+ 35 41 42 43 48 50 VSS
c35 52 VSS 5.10117e-19 $X=0.513 $Y=0.1765
c36 50 VSS 0.00117789f $X=0.513 $Y=0.0985
c37 49 VSS 0.00112176f $X=0.513 $Y=0.07
c38 48 VSS 0.00292471f $X=0.512 $Y=0.127
c39 46 VSS 6.07272e-19 $X=0.513 $Y=0.189
c40 44 VSS 4.93718e-20 $X=0.503 $Y=0.198
c41 43 VSS 4.1269e-19 $X=0.502 $Y=0.198
c42 42 VSS 8.46035e-21 $X=0.468 $Y=0.198
c43 41 VSS 4.70878e-19 $X=0.45 $Y=0.198
c44 36 VSS 0.0019286f $X=0.504 $Y=0.198
c45 35 VSS 0.00146362f $X=0.468 $Y=0.036
c46 34 VSS 0.00296425f $X=0.45 $Y=0.036
c47 33 VSS 3.35992e-19 $X=0.417 $Y=0.036
c48 32 VSS 0.00142296f $X=0.414 $Y=0.036
c49 31 VSS 0.00672869f $X=0.396 $Y=0.036
c50 30 VSS 0.00142296f $X=0.36 $Y=0.036
c51 29 VSS 3.35992e-19 $X=0.342 $Y=0.036
c52 28 VSS 0.00311761f $X=0.339 $Y=0.036
c53 27 VSS 0.00146362f $X=0.306 $Y=0.036
c54 26 VSS 0.00340162f $X=0.288 $Y=0.036
c55 25 VSS 0.00146362f $X=0.252 $Y=0.036
c56 24 VSS 0.00418453f $X=0.234 $Y=0.036
c57 23 VSS 0.00357414f $X=0.486 $Y=0.036
c58 19 VSS 0.00220422f $X=0.216 $Y=0.036
c59 16 VSS 0.00700674f $X=0.504 $Y=0.036
c60 15 VSS 0.0023085f $X=0.432 $Y=0.2025
c61 11 VSS 5.70099e-19 $X=0.449 $Y=0.2025
c62 9 VSS 2.69461e-19 $X=0.484 $Y=0.0675
c63 1 VSS 5.61153e-19 $X=0.233 $Y=0.0675
r64 51 52 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.164 $X2=0.513 $Y2=0.1765
r65 49 50 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.07 $X2=0.513 $Y2=0.0985
r66 48 51 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.127 $X2=0.513 $Y2=0.164
r67 48 50 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.127 $X2=0.513 $Y2=0.0985
r68 46 52 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.513 $Y2=0.1765
r69 45 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.07
r70 43 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.502
+ $Y=0.198 $X2=0.503 $Y2=0.198
r71 42 43 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.198 $X2=0.502 $Y2=0.198
r72 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.198 $X2=0.468 $Y2=0.198
r73 38 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.45 $Y2=0.198
r74 36 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.198 $X2=0.513 $Y2=0.189
r75 36 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.198 $X2=0.503 $Y2=0.198
r76 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r77 33 34 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.417
+ $Y=0.036 $X2=0.45 $Y2=0.036
r78 32 33 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.417 $Y2=0.036
r79 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r80 30 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.396 $Y2=0.036
r81 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r82 28 29 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.339
+ $Y=0.036 $X2=0.342 $Y2=0.036
r83 27 28 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.339 $Y2=0.036
r84 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r85 25 26 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r86 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r87 22 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.468 $Y2=0.036
r88 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036 $X2=0.486
+ $Y2=0.036
r89 18 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.234 $Y2=0.036
r90 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r91 16 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.036 $X2=0.513 $Y2=0.045
r92 16 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.486 $Y2=0.036
r93 15 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r94 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r95 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r96 9 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0675 $X2=0.486 $Y2=0.036
r97 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.0675 $X2=0.484 $Y2=0.0675
r98 5 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r99 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r100 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./AOI332xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI332xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 noxref_14 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_15 N_A2_M1_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_A1_M2_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_16 N_B1_M3_g N_Y_M3_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_17 N_B2_M4_g noxref_16 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 VSS N_B3_M5_g noxref_17 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_18 N_C2_M6_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_Y_M7_d N_C1_M7_g noxref_18 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 noxref_11 N_A3_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M9 VDD N_A2_M9_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M10 noxref_11 N_A1_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M11 noxref_12 N_B1_M11_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M12 noxref_11 N_B2_M12_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M13 noxref_12 N_B3_M13_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M14 N_Y_M14_d N_C2_M14_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M15 noxref_12 N_C1_M15_g N_Y_M15_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
*
* 
* .include "AOI332xp33_ASAP7_75t_L.pex.sp.AOI332XP33_ASAP7_75T_L.pxi"
* BEGIN of "./AOI332xp33_ASAP7_75t_L.pex.sp.AOI332XP33_ASAP7_75T_L.pxi"
* File: AOI332xp33_ASAP7_75t_L.pex.sp.AOI332XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:16:17 2017
* 
x_PM_AOI332XP33_ASAP7_75T_L%A3 N_A3_M0_g N_A3_c_2_p N_A3_M8_g A3 VSS
+ PM_AOI332XP33_ASAP7_75T_L%A3
x_PM_AOI332XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_6_n N_A2_M9_g A2 VSS
+ PM_AOI332XP33_ASAP7_75T_L%A2
x_PM_AOI332XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_18_n N_A1_M10_g A1 VSS
+ PM_AOI332XP33_ASAP7_75T_L%A1
x_PM_AOI332XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_29_n N_B1_M11_g B1 VSS
+ PM_AOI332XP33_ASAP7_75T_L%B1
x_PM_AOI332XP33_ASAP7_75T_L%B2 N_B2_M4_g N_B2_c_42_n N_B2_M12_g B2 VSS
+ PM_AOI332XP33_ASAP7_75T_L%B2
x_PM_AOI332XP33_ASAP7_75T_L%B3 N_B3_M5_g N_B3_c_55_n N_B3_M13_g B3 VSS
+ PM_AOI332XP33_ASAP7_75T_L%B3
x_PM_AOI332XP33_ASAP7_75T_L%C2 N_C2_M6_g N_C2_c_67_n N_C2_M14_g C2 VSS
+ PM_AOI332XP33_ASAP7_75T_L%C2
x_PM_AOI332XP33_ASAP7_75T_L%C1 N_C1_M7_g N_C1_c_78_n N_C1_M15_g C1 VSS
+ PM_AOI332XP33_ASAP7_75T_L%C1
x_PM_AOI332XP33_ASAP7_75T_L%Y N_Y_M3_s N_Y_M2_d N_Y_M7_d N_Y_M15_s N_Y_M14_d
+ N_Y_c_110_n N_Y_c_87_n N_Y_c_99_n N_Y_c_88_n N_Y_c_91_n N_Y_c_107_n N_Y_c_93_n
+ N_Y_c_108_n N_Y_c_95_n N_Y_c_97_n N_Y_c_121_p N_Y_c_100_n N_Y_c_109_n
+ N_Y_c_102_n N_Y_c_117_n Y N_Y_c_104_n VSS PM_AOI332XP33_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_A2_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A3_c_2_p N_A2_c_6_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A3 A2 0.00653171f $X=0.081 $Y=0.115 $X2=0.135 $Y2=0.115
cc_4 N_A3_M0_g N_A1_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 N_A2_M1_g N_A1_M2_g 0.00327995f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_6 N_A2_c_6_n N_A1_c_18_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_7 A2 A1 0.00466039f $X=0.135 $Y=0.115 $X2=0.081 $Y2=0.115
cc_8 N_A2_M1_g N_B1_M3_g 2.71887e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_9 VSS N_A2_M1_g 3.62029e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_10 VSS A2 0.0012376f $X=0.135 $Y=0.115 $X2=0 $Y2=0
cc_11 A2 N_Y_c_87_n 5.87506e-19 $X=0.135 $Y=0.115 $X2=0 $Y2=0
cc_12 A2 N_Y_c_88_n 4.59821e-19 $X=0.135 $Y=0.115 $X2=0 $Y2=0
cc_13 N_A1_M2_g N_B1_M3_g 0.0036939f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_A1_c_18_n N_B1_c_29_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 A1 B1 0.00406615f $X=0.189 $Y=0.115 $X2=0.081 $Y2=0.115
cc_16 N_A1_M2_g N_B2_M4_g 3.06651e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 VSS N_A1_M2_g 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_18 VSS A1 0.0012322f $X=0.189 $Y=0.115 $X2=0 $Y2=0
cc_19 A1 N_Y_c_87_n 0.0013295f $X=0.189 $Y=0.115 $X2=0 $Y2=0
cc_20 N_B1_M3_g N_B2_M4_g 0.00371573f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_21 N_B1_c_29_n N_B2_c_42_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_22 B1 B2 0.00483372f $X=0.243 $Y=0.116 $X2=0.135 $Y2=0.115
cc_23 N_B1_M3_g N_B3_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_24 VSS N_B1_M3_g 3.62029e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_25 VSS B1 0.0012322f $X=0.243 $Y=0.116 $X2=0 $Y2=0
cc_26 B1 N_Y_c_87_n 0.0013295f $X=0.243 $Y=0.116 $X2=0 $Y2=0
cc_27 N_B1_M3_g N_Y_c_91_n 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_28 B1 N_Y_c_91_n 0.00124805f $X=0.243 $Y=0.116 $X2=0 $Y2=0
cc_29 N_B2_M4_g N_B3_M5_g 0.0036939f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_30 N_B2_c_42_n N_B3_c_55_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_31 B2 B3 0.00483372f $X=0.296 $Y=0.115 $X2=0.189 $Y2=0.115
cc_32 N_B2_M4_g N_C2_M6_g 2.71887e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_33 VSS N_B2_M4_g 2.68514e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_34 VSS B2 0.00121543f $X=0.296 $Y=0.115 $X2=0 $Y2=0
cc_35 VSS N_B2_M4_g 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B2_M4_g N_Y_c_93_n 3.48613e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_37 B2 N_Y_c_93_n 0.00124805f $X=0.296 $Y=0.115 $X2=0 $Y2=0
cc_38 N_B3_M5_g N_C2_M6_g 0.00333077f $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_39 N_B3_c_55_n N_C2_c_67_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_40 B3 C2 0.00406615f $X=0.349 $Y=0.115 $X2=0.243 $Y2=0.116
cc_41 N_B3_M5_g N_C1_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_42 VSS N_B3_M5_g 3.47199e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_43 VSS B3 5.30079e-19 $X=0.349 $Y=0.115 $X2=0 $Y2=0
cc_44 N_B3_M5_g N_Y_c_95_n 2.56935e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_45 B3 N_Y_c_95_n 0.00123064f $X=0.349 $Y=0.115 $X2=0 $Y2=0
cc_46 N_C2_M6_g N_C1_M7_g 0.0036939f $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_47 N_C2_c_67_n N_C1_c_78_n 9.33263e-19 $X=0.405 $Y=0.135 $X2=0.297 $Y2=0.135
cc_48 C2 C1 0.00477924f $X=0.406 $Y=0.114 $X2=0.296 $Y2=0.115
cc_49 VSS N_C2_M6_g 3.57119e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_50 VSS C2 5.37372e-19 $X=0.406 $Y=0.114 $X2=0 $Y2=0
cc_51 N_C2_M6_g N_Y_c_97_n 2.56935e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_52 C2 N_Y_c_97_n 0.00123064f $X=0.406 $Y=0.114 $X2=0 $Y2=0
cc_53 VSS N_C1_M7_g 2.15135e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_54 C1 N_Y_c_99_n 0.0013399f $X=0.459 $Y=0.115 $X2=0 $Y2=0
cc_55 N_C1_M7_g N_Y_c_100_n 2.64276e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_56 C1 N_Y_c_100_n 0.00124805f $X=0.459 $Y=0.115 $X2=0 $Y2=0
cc_57 N_C1_M7_g N_Y_c_102_n 2.76185e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_58 C1 N_Y_c_102_n 0.0012322f $X=0.459 $Y=0.115 $X2=0 $Y2=0
cc_59 C1 N_Y_c_104_n 0.00391435f $X=0.459 $Y=0.115 $X2=0 $Y2=0
cc_60 VSS N_Y_c_87_n 0.00138157f $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_61 VSS N_Y_c_88_n 2.88662e-19 $X=0.2085 $Y=0.198 $X2=0 $Y2=0
cc_62 VSS N_Y_c_107_n 2.88662e-19 $X=0.254 $Y=0.198 $X2=0 $Y2=0
cc_63 VSS N_Y_c_108_n 2.88662e-19 $X=0.315 $Y=0.198 $X2=0 $Y2=0
cc_64 VSS N_Y_c_109_n 2.99055e-19 $X=0.324 $Y=0.198 $X2=0 $Y2=0
cc_65 VSS N_Y_c_110_n 0.00333582f $X=0.378 $Y=0.2025 $X2=0 $Y2=0
cc_66 VSS N_Y_c_110_n 0.00371671f $X=0.484 $Y=0.2025 $X2=0 $Y2=0
cc_67 VSS N_Y_c_110_n 0.00250965f $X=0.4515 $Y=0.234 $X2=0 $Y2=0
cc_68 VSS N_Y_c_99_n 0.00138157f $X=0.484 $Y=0.2025 $X2=0 $Y2=0
cc_69 VSS N_Y_c_109_n 4.54465e-19 $X=0.378 $Y=0.2025 $X2=0 $Y2=0
cc_70 VSS N_Y_c_109_n 0.00365373f $X=0.4515 $Y=0.234 $X2=0 $Y2=0
cc_71 VSS N_Y_c_102_n 0.00365373f $X=0.486 $Y=0.234 $X2=0 $Y2=0
cc_72 VSS N_Y_c_117_n 0.00284922f $X=0.484 $Y=0.2025 $X2=0 $Y2=0
cc_73 VSS Y 4.01247e-19 $X=0.484 $Y=0.2025 $X2=0 $Y2=0
cc_74 VSS N_Y_c_107_n 3.48201e-19 $X=0.288 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_75 VSS N_Y_c_108_n 3.30547e-19 $X=0.339 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_76 VSS N_Y_c_121_p 3.30547e-19 $X=0.45 $Y=0.036 $X2=0.135 $Y2=0.0675

* END of "./AOI332xp33_ASAP7_75t_L.pex.sp.AOI332XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI333xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:16:40 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI333xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI333xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI333xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:16:40 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI333XP33_ASAP7_75T_L%C3 2 5 7 10 VSS
c4 10 VSS 0.00613146f $X=0.073 $Y=0.114
c5 5 VSS 0.00238289f $X=0.081 $Y=0.135
c6 2 VSS 0.062704f $X=0.081 $Y=0.0675
r7 10 13 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.114 $X2=0.081 $Y2=0.135
r8 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r9 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r10 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI333XP33_ASAP7_75T_L%C2 2 5 7 10 VSS
c11 10 VSS 0.00174706f $X=0.129 $Y=0.116
c12 5 VSS 0.00123757f $X=0.135 $Y=0.135
c13 2 VSS 0.0598541f $X=0.135 $Y=0.0675
r14 10 15 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.116 $X2=0.135 $Y2=0.135
r15 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI333XP33_ASAP7_75T_L%C1 2 5 7 10 VSS
c11 10 VSS 0.00101969f $X=0.187 $Y=0.115
c12 5 VSS 0.00121257f $X=0.189 $Y=0.135
c13 2 VSS 0.0608354f $X=0.189 $Y=0.0675
r14 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI333XP33_ASAP7_75T_L%B1 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.243 $Y=0.116
c14 5 VSS 0.00111336f $X=0.243 $Y=0.135
c15 2 VSS 0.0617786f $X=0.243 $Y=0.0675
r16 10 13 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.116 $X2=0.243 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI333XP33_ASAP7_75T_L%B2 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.296 $Y=0.115
c14 5 VSS 0.00112198f $X=0.297 $Y=0.135
c15 2 VSS 0.0616432f $X=0.297 $Y=0.0675
r16 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.115 $X2=0.297 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AOI333XP33_ASAP7_75T_L%B3 2 5 7 10 VSS
c12 10 VSS 7.27237e-19 $X=0.346 $Y=0.115
c13 5 VSS 0.00111185f $X=0.351 $Y=0.135
c14 2 VSS 0.0615515f $X=0.351 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.115 $X2=0.351 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AOI333XP33_ASAP7_75T_L%A3 2 5 7 10 VSS
c12 10 VSS 7.27237e-19 $X=0.408 $Y=0.115
c13 5 VSS 0.00111774f $X=0.405 $Y=0.135
c14 2 VSS 0.0615416f $X=0.405 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.115 $X2=0.405 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AOI333XP33_ASAP7_75T_L%A2 2 5 7 10 VSS
c12 10 VSS 4.78074e-19 $X=0.457 $Y=0.115
c13 5 VSS 0.00114557f $X=0.459 $Y=0.135
c14 2 VSS 0.0623815f $X=0.459 $Y=0.0675
r15 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.115 $X2=0.459 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_AOI333XP33_ASAP7_75T_L%A1 2 5 7 10 VSS
c9 10 VSS 4.90626e-19 $X=0.521 $Y=0.115
c10 5 VSS 0.00171677f $X=0.513 $Y=0.135
c11 2 VSS 0.0671256f $X=0.513 $Y=0.0675
r12 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.115 $X2=0.513 $Y2=0.135
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_AOI333XP33_ASAP7_75T_L%Y 1 2 6 11 12 15 16 19 24 28 29 30 31 32 33 35
+ 37 38 39 40 41 45 54 55 56 62 64 VSS
c38 66 VSS 5.10117e-19 $X=0.567 $Y=0.1765
c39 64 VSS 0.00117789f $X=0.567 $Y=0.0985
c40 63 VSS 0.00112176f $X=0.567 $Y=0.07
c41 62 VSS 0.00292471f $X=0.572 $Y=0.127
c42 60 VSS 6.07272e-19 $X=0.567 $Y=0.189
c43 58 VSS 4.0892e-19 $X=0.531 $Y=0.198
c44 57 VSS 3.28227e-19 $X=0.522 $Y=0.198
c45 56 VSS 1.7724e-19 $X=0.515 $Y=0.198
c46 55 VSS 4.2636e-19 $X=0.504 $Y=0.198
c47 54 VSS 8.46035e-21 $X=0.468 $Y=0.198
c48 53 VSS 3.93699e-19 $X=0.45 $Y=0.198
c49 45 VSS 3.25927e-19 $X=0.432 $Y=0.198
c50 43 VSS 0.00335467f $X=0.558 $Y=0.198
c51 42 VSS 8.36318e-19 $X=0.531 $Y=0.036
c52 41 VSS 0.00142296f $X=0.522 $Y=0.036
c53 40 VSS 0.00344621f $X=0.504 $Y=0.036
c54 39 VSS 0.00142296f $X=0.468 $Y=0.036
c55 38 VSS 0.00329285f $X=0.45 $Y=0.036
c56 37 VSS 0.00142296f $X=0.414 $Y=0.036
c57 36 VSS 0.00688205f $X=0.396 $Y=0.036
c58 35 VSS 0.00142296f $X=0.36 $Y=0.036
c59 34 VSS 2.83817e-19 $X=0.342 $Y=0.036
c60 33 VSS 0.00320869f $X=0.34 $Y=0.036
c61 32 VSS 0.00146362f $X=0.306 $Y=0.036
c62 31 VSS 0.00340162f $X=0.288 $Y=0.036
c63 30 VSS 0.00146362f $X=0.252 $Y=0.036
c64 29 VSS 0.0041898f $X=0.234 $Y=0.036
c65 28 VSS 0.00224055f $X=0.54 $Y=0.036
c66 24 VSS 0.00220422f $X=0.216 $Y=0.036
c67 21 VSS 0.00607902f $X=0.558 $Y=0.036
c68 19 VSS 0.00113516f $X=0.538 $Y=0.2025
c69 15 VSS 0.0023085f $X=0.432 $Y=0.2025
c70 11 VSS 5.91014e-19 $X=0.449 $Y=0.2025
c71 9 VSS 2.69461e-19 $X=0.538 $Y=0.0675
c72 1 VSS 5.61153e-19 $X=0.233 $Y=0.0675
r73 65 66 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.164 $X2=0.567 $Y2=0.1765
r74 63 64 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.07 $X2=0.567 $Y2=0.0985
r75 62 65 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.127 $X2=0.567 $Y2=0.164
r76 62 64 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.127 $X2=0.567 $Y2=0.0985
r77 60 66 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.567 $Y2=0.1765
r78 59 63 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.045 $X2=0.567 $Y2=0.07
r79 57 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.198 $X2=0.531 $Y2=0.198
r80 56 57 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.515
+ $Y=0.198 $X2=0.522 $Y2=0.198
r81 55 56 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.198 $X2=0.515 $Y2=0.198
r82 54 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.198 $X2=0.504 $Y2=0.198
r83 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.198 $X2=0.468 $Y2=0.198
r84 51 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.198 $X2=0.531 $Y2=0.198
r85 45 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.45 $Y2=0.198
r86 43 60 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.198 $X2=0.567 $Y2=0.189
r87 43 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.198 $X2=0.54 $Y2=0.198
r88 41 42 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.531 $Y2=0.036
r89 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.522 $Y2=0.036
r90 39 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.504 $Y2=0.036
r91 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r92 37 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.45 $Y2=0.036
r93 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r94 35 36 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.396 $Y2=0.036
r95 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r96 33 34 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.34
+ $Y=0.036 $X2=0.342 $Y2=0.036
r97 32 33 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.34 $Y2=0.036
r98 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r99 30 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r100 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r101 27 42 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.531 $Y2=0.036
r102 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r103 23 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.234 $Y2=0.036
r104 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r105 21 59 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.036 $X2=0.567 $Y2=0.045
r106 21 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.54 $Y2=0.036
r107 19 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.198 $X2=0.54
+ $Y2=0.198
r108 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.538 $Y2=0.2025
r109 15 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198
+ $X2=0.432 $Y2=0.198
r110 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r111 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r112 9 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r113 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.538 $Y2=0.0675
r114 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r115 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r116 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./AOI333xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI333xp33_ASAP7_75t_L  VSS VDD C3 C2 C1 B1 B2 B3 A3 A2 A1 Y
* 
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* B3	B3
* B2	B2
* B1	B1
* C1	C1
* C2	C2
* C3	C3
M0 noxref_15 N_C3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_16 N_C2_M1_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_C1_M2_g noxref_16 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_17 N_B1_M3_g N_Y_M3_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_18 N_B2_M4_g noxref_17 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 VSS N_B3_M5_g noxref_18 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_19 N_A3_M6_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_20 N_A2_M7_g noxref_19 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_Y_M8_d N_A1_M8_g noxref_20 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 noxref_12 N_C3_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M10 VDD N_C2_M10_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M11 noxref_12 N_C1_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M12 noxref_13 N_B1_M12_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M13 noxref_12 N_B2_M13_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M14 noxref_13 N_B3_M14_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M15 N_Y_M15_d N_A3_M15_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M16 noxref_13 N_A2_M16_g N_Y_M16_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M17 N_Y_M17_d N_A1_M17_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
*
* 
* .include "AOI333xp33_ASAP7_75t_L.pex.sp.AOI333XP33_ASAP7_75T_L.pxi"
* BEGIN of "./AOI333xp33_ASAP7_75t_L.pex.sp.AOI333XP33_ASAP7_75T_L.pxi"
* File: AOI333xp33_ASAP7_75t_L.pex.sp.AOI333XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:16:40 2017
* 
x_PM_AOI333XP33_ASAP7_75T_L%C3 N_C3_M0_g N_C3_c_2_p N_C3_M9_g C3 VSS
+ PM_AOI333XP33_ASAP7_75T_L%C3
x_PM_AOI333XP33_ASAP7_75T_L%C2 N_C2_M1_g N_C2_c_6_n N_C2_M10_g C2 VSS
+ PM_AOI333XP33_ASAP7_75T_L%C2
x_PM_AOI333XP33_ASAP7_75T_L%C1 N_C1_M2_g N_C1_c_18_n N_C1_M11_g C1 VSS
+ PM_AOI333XP33_ASAP7_75T_L%C1
x_PM_AOI333XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_29_n N_B1_M12_g B1 VSS
+ PM_AOI333XP33_ASAP7_75T_L%B1
x_PM_AOI333XP33_ASAP7_75T_L%B2 N_B2_M4_g N_B2_c_42_n N_B2_M13_g B2 VSS
+ PM_AOI333XP33_ASAP7_75T_L%B2
x_PM_AOI333XP33_ASAP7_75T_L%B3 N_B3_M5_g N_B3_c_55_n N_B3_M14_g B3 VSS
+ PM_AOI333XP33_ASAP7_75T_L%B3
x_PM_AOI333XP33_ASAP7_75T_L%A3 N_A3_M6_g N_A3_c_67_n N_A3_M15_g A3 VSS
+ PM_AOI333XP33_ASAP7_75T_L%A3
x_PM_AOI333XP33_ASAP7_75T_L%A2 N_A2_M7_g N_A2_c_79_n N_A2_M16_g A2 VSS
+ PM_AOI333XP33_ASAP7_75T_L%A2
x_PM_AOI333XP33_ASAP7_75T_L%A1 N_A1_M8_g N_A1_c_91_n N_A1_M17_g A1 VSS
+ PM_AOI333XP33_ASAP7_75T_L%A1
x_PM_AOI333XP33_ASAP7_75T_L%Y N_Y_M3_s N_Y_M2_d N_Y_M8_d N_Y_M16_s N_Y_M15_d
+ N_Y_c_124_n N_Y_M17_d N_Y_c_127_n N_Y_c_98_n N_Y_c_114_n N_Y_c_99_n
+ N_Y_c_102_n N_Y_c_121_n N_Y_c_104_n N_Y_c_122_n N_Y_c_106_n N_Y_c_108_n
+ N_Y_c_134_p N_Y_c_110_n N_Y_c_135_p N_Y_c_115_n N_Y_c_123_n N_Y_c_112_n
+ N_Y_c_131_n N_Y_c_117_n Y N_Y_c_118_n VSS PM_AOI333XP33_ASAP7_75T_L%Y
cc_1 N_C3_M0_g N_C2_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_C3_c_2_p N_C2_c_6_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 C3 C2 0.00653171f $X=0.073 $Y=0.114 $X2=0.129 $Y2=0.116
cc_4 N_C3_M0_g N_C1_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 N_C2_M1_g N_C1_M2_g 0.00327995f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_6 N_C2_c_6_n N_C1_c_18_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_7 C2 C1 0.00466039f $X=0.129 $Y=0.116 $X2=0.073 $Y2=0.114
cc_8 N_C2_M1_g N_B1_M3_g 2.71887e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_9 VSS N_C2_M1_g 3.62029e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_10 VSS C2 0.0012376f $X=0.129 $Y=0.116 $X2=0 $Y2=0
cc_11 C2 N_Y_c_98_n 5.87506e-19 $X=0.129 $Y=0.116 $X2=0 $Y2=0
cc_12 C2 N_Y_c_99_n 4.59979e-19 $X=0.129 $Y=0.116 $X2=0 $Y2=0
cc_13 N_C1_M2_g N_B1_M3_g 0.0036939f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_C1_c_18_n N_B1_c_29_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 C1 B1 0.00406615f $X=0.187 $Y=0.115 $X2=0.073 $Y2=0.114
cc_16 N_C1_M2_g N_B2_M4_g 3.06651e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 VSS N_C1_M2_g 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_18 VSS C1 0.0012322f $X=0.187 $Y=0.115 $X2=0 $Y2=0
cc_19 C1 N_Y_c_98_n 0.0013295f $X=0.187 $Y=0.115 $X2=0 $Y2=0
cc_20 N_B1_M3_g N_B2_M4_g 0.00371573f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_21 N_B1_c_29_n N_B2_c_42_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_22 B1 B2 0.00483372f $X=0.243 $Y=0.116 $X2=0.129 $Y2=0.116
cc_23 N_B1_M3_g N_B3_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_24 VSS N_B1_M3_g 3.62029e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_25 VSS B1 0.0012322f $X=0.243 $Y=0.116 $X2=0 $Y2=0
cc_26 B1 N_Y_c_98_n 0.0013295f $X=0.243 $Y=0.116 $X2=0 $Y2=0
cc_27 N_B1_M3_g N_Y_c_102_n 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_28 B1 N_Y_c_102_n 0.00124805f $X=0.243 $Y=0.116 $X2=0 $Y2=0
cc_29 N_B2_M4_g N_B3_M5_g 0.0036939f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_30 N_B2_c_42_n N_B3_c_55_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_31 B2 B3 0.00483372f $X=0.296 $Y=0.115 $X2=0.187 $Y2=0.115
cc_32 N_B2_M4_g N_A3_M6_g 2.71887e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_33 VSS N_B2_M4_g 2.68514e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_34 VSS B2 0.00121543f $X=0.296 $Y=0.115 $X2=0 $Y2=0
cc_35 VSS N_B2_M4_g 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B2_M4_g N_Y_c_104_n 3.48613e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_37 B2 N_Y_c_104_n 0.00124805f $X=0.296 $Y=0.115 $X2=0 $Y2=0
cc_38 N_B3_M5_g N_A3_M6_g 0.00333077f $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_39 N_B3_c_55_n N_A3_c_67_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_40 B3 A3 0.00406615f $X=0.346 $Y=0.115 $X2=0.243 $Y2=0.116
cc_41 N_B3_M5_g N_A2_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_42 VSS N_B3_M5_g 3.47199e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_43 VSS B3 5.30079e-19 $X=0.346 $Y=0.115 $X2=0 $Y2=0
cc_44 N_B3_M5_g N_Y_c_106_n 2.56935e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_45 B3 N_Y_c_106_n 0.00123064f $X=0.346 $Y=0.115 $X2=0 $Y2=0
cc_46 N_A3_M6_g N_A2_M7_g 0.0036939f $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_47 N_A3_c_67_n N_A2_c_79_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.297 $Y2=0.135
cc_48 A3 A2 0.00483372f $X=0.408 $Y=0.115 $X2=0.296 $Y2=0.115
cc_49 N_A3_M6_g N_A1_M8_g 3.06651e-19 $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_50 VSS N_A3_M6_g 3.37279e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_51 VSS A3 5.22785e-19 $X=0.408 $Y=0.115 $X2=0 $Y2=0
cc_52 N_A3_M6_g N_Y_c_108_n 2.45924e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_53 A3 N_Y_c_108_n 0.00123064f $X=0.408 $Y=0.115 $X2=0 $Y2=0
cc_54 N_A2_M7_g N_A1_M8_g 0.00376655f $X=0.459 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_55 N_A2_c_79_n N_A1_c_91_n 9.33263e-19 $X=0.459 $Y=0.135 $X2=0.351 $Y2=0.135
cc_56 A2 A1 0.0048308f $X=0.457 $Y=0.115 $X2=0.346 $Y2=0.115
cc_57 VSS N_A2_M7_g 2.38303e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_A2_M7_g N_Y_c_110_n 3.38929e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_59 A2 N_Y_c_110_n 0.00123064f $X=0.457 $Y=0.115 $X2=0 $Y2=0
cc_60 N_A2_M7_g N_Y_c_112_n 2.76185e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_61 A2 N_Y_c_112_n 0.0012322f $X=0.457 $Y=0.115 $X2=0 $Y2=0
cc_62 A1 N_Y_c_114_n 0.0013295f $X=0.521 $Y=0.115 $X2=0 $Y2=0
cc_63 N_A1_M8_g N_Y_c_115_n 2.56935e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_64 A1 N_Y_c_115_n 0.00123064f $X=0.521 $Y=0.115 $X2=0 $Y2=0
cc_65 A1 N_Y_c_117_n 0.00121543f $X=0.521 $Y=0.115 $X2=0 $Y2=0
cc_66 A1 N_Y_c_118_n 0.00391435f $X=0.521 $Y=0.115 $X2=0 $Y2=0
cc_67 VSS N_Y_c_98_n 0.00138157f $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_68 VSS N_Y_c_99_n 2.9391e-19 $X=0.2085 $Y=0.198 $X2=0 $Y2=0
cc_69 VSS N_Y_c_121_n 2.9391e-19 $X=0.254 $Y=0.198 $X2=0 $Y2=0
cc_70 VSS N_Y_c_122_n 2.9391e-19 $X=0.315 $Y=0.198 $X2=0 $Y2=0
cc_71 VSS N_Y_c_123_n 3.22079e-19 $X=0.324 $Y=0.198 $X2=0 $Y2=0
cc_72 VSS N_Y_c_124_n 0.003332f $X=0.378 $Y=0.2025 $X2=0 $Y2=0
cc_73 VSS N_Y_c_124_n 0.00355403f $X=0.486 $Y=0.2025 $X2=0 $Y2=0
cc_74 VSS N_Y_c_124_n 0.00250965f $X=0.486 $Y=0.234 $X2=0 $Y2=0
cc_75 VSS N_Y_c_127_n 0.00337424f $X=0.486 $Y=0.2025 $X2=0 $Y2=0
cc_76 VSS N_Y_c_127_n 3.14809e-19 $X=0.486 $Y=0.234 $X2=0 $Y2=0
cc_77 VSS N_Y_c_123_n 4.6373e-19 $X=0.378 $Y=0.2025 $X2=0 $Y2=0
cc_78 VSS N_Y_c_123_n 0.00881219f $X=0.486 $Y=0.234 $X2=0 $Y2=0
cc_79 VSS N_Y_c_131_n 0.00233206f $X=0.486 $Y=0.2025 $X2=0 $Y2=0
cc_80 VSS N_Y_c_121_n 3.48201e-19 $X=0.288 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_81 VSS N_Y_c_122_n 3.4467e-19 $X=0.34 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_82 VSS N_Y_c_134_p 3.48201e-19 $X=0.45 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_83 VSS N_Y_c_135_p 3.48201e-19 $X=0.504 $Y=0.036 $X2=0.135 $Y2=0.0675

* END of "./AOI333xp33_ASAP7_75t_L.pex.sp.AOI333XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: AOI33xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:17:02 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AOI33xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./AOI33xp33_ASAP7_75t_L.pex.sp.pex"
* File: AOI33xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:17:02 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AOI33XP33_ASAP7_75T_L%A1 2 5 7 12 18 20 VSS
c8 20 VSS 0.00201554f $X=0.063 $Y=0.135
c9 18 VSS 8.46268e-19 $X=0.027 $Y=0.135
c10 12 VSS 0.0137164f $X=0.027 $Y=0.08
c11 5 VSS 0.0103458f $X=0.081 $Y=0.135
c12 2 VSS 0.0605822f $X=0.081 $Y=0.0675
r13 20 21 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.063 $Y=0.135 $X2=0.063
+ $Y2=0.135
r14 18 20 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.063 $Y2=0.135
r15 10 18 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.126 $X2=0.027 $Y2=0.135
r16 10 12 3.12346 $w=1.8e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.08
r17 5 21 22.5 $w=1.6e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.063 $Y2=0.135
r18 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AOI33XP33_ASAP7_75T_L%A2 2 5 7 11 12 13 14 15 16 20 22 29 31 VSS
c24 31 VSS 0.00618103f $X=0.024 $Y=0.233
c25 29 VSS 4.48164e-19 $X=0.135 $Y=0.1665
c26 22 VSS 0.0055343f $X=0.135 $Y=0.135
c27 20 VSS 5.91281e-19 $X=0.135 $Y=0.189
c28 16 VSS 1.77619e-19 $X=0.1125 $Y=0.198
c29 15 VSS 5.2199e-19 $X=0.099 $Y=0.198
c30 14 VSS 0.0013652f $X=0.09 $Y=0.198
c31 13 VSS 0.00303979f $X=0.064 $Y=0.198
c32 12 VSS 9.00122e-19 $X=0.027 $Y=0.198
c33 11 VSS 9.14602e-19 $X=0.126 $Y=0.198
c34 10 VSS 0.00360474f $X=0.018 $Y=0.225
c35 5 VSS 0.00101464f $X=0.135 $Y=0.135
c36 2 VSS 0.0576487f $X=0.135 $Y=0.0675
r37 28 29 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.1665
r38 22 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r39 20 29 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.135 $Y2=0.1665
r40 15 16 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.198 $X2=0.1125 $Y2=0.198
r41 14 15 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.198 $X2=0.099 $Y2=0.198
r42 13 14 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.198 $X2=0.09 $Y2=0.198
r43 12 13 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.198 $X2=0.064 $Y2=0.198
r44 11 20 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.126 $Y=0.198 $X2=0.135 $Y2=0.189
r45 11 16 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.198 $X2=0.1125 $Y2=0.198
r46 10 31 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.234
r47 9 12 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.207 $X2=0.027 $Y2=0.198
r48 9 10 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.207 $X2=0.018 $Y2=0.225
r49 5 22 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r50 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r51 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AOI33XP33_ASAP7_75T_L%A3 2 5 7 11 15 17 18 VSS
c15 18 VSS 3.22517e-19 $X=0.2015 $Y=0.189
c16 17 VSS 0.00115008f $X=0.186 $Y=0.198
c17 15 VSS 3.09574e-19 $X=0.189 $Y=0.1765
c18 11 VSS 7.79063e-19 $X=0.189 $Y=0.135
c19 5 VSS 0.00101548f $X=0.189 $Y=0.135
c20 2 VSS 0.0585669f $X=0.189 $Y=0.0675
r21 17 18 0.533258 $w=4.3e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.2015
+ $Y=0.198 $X2=0.2015 $Y2=0.189
r22 15 18 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.1765 $X2=0.189 $Y2=0.189
r23 14 15 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.1765
r24 11 14 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.164
r25 5 11 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r26 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AOI33XP33_ASAP7_75T_L%B1 2 5 7 11 VSS
c14 11 VSS 0.00130981f $X=0.238 $Y=0.115
c15 5 VSS 9.30047e-19 $X=0.243 $Y=0.135
c16 2 VSS 0.0593517f $X=0.243 $Y=0.0675
r17 11 15 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.115 $X2=0.243 $Y2=0.135
r18 5 15 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r19 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r20 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AOI33XP33_ASAP7_75T_L%B2 2 5 7 10 VSS
c12 10 VSS 3.66617e-19 $X=0.303 $Y=0.122
c13 5 VSS 9.83461e-19 $X=0.297 $Y=0.135
c14 2 VSS 0.0593926f $X=0.297 $Y=0.0675
r15 10 13 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.122 $X2=0.297 $Y2=0.135
r16 5 13 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AOI33XP33_ASAP7_75T_L%B3 2 5 7 10 VSS
c9 10 VSS 6.52219e-19 $X=0.353 $Y=0.122
c10 5 VSS 0.00139335f $X=0.351 $Y=0.135
c11 2 VSS 0.0629245f $X=0.351 $Y=0.0675
r12 10 13 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.122 $X2=0.351 $Y2=0.135
r13 5 13 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.216
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_AOI33XP33_ASAP7_75T_L%Y 1 2 6 7 10 11 14 18 19 23 25 26 27 28 37 38
+ 39 41 47 50 VSS
c26 48 VSS 7.1665e-19 $X=0.405 $Y=0.1765
c27 47 VSS 0.0043346f $X=0.405 $Y=0.164
c28 46 VSS 4.39352e-19 $X=0.405 $Y=0.07
c29 45 VSS 8.85605e-19 $X=0.405 $Y=0.063
c30 44 VSS 6.07272e-19 $X=0.405 $Y=0.189
c31 43 VSS 0.00336642f $X=0.405 $Y=0.045
c32 42 VSS 4.63286e-19 $X=0.369 $Y=0.198
c33 41 VSS 5.16928e-19 $X=0.36 $Y=0.198
c34 40 VSS 2.26742e-19 $X=0.342 $Y=0.198
c35 39 VSS 4.06957e-19 $X=0.338 $Y=0.198
c36 38 VSS 7.99121e-21 $X=0.306 $Y=0.198
c37 37 VSS 5.00504e-19 $X=0.288 $Y=0.198
c38 29 VSS 0.00354587f $X=0.396 $Y=0.198
c39 28 VSS 0.00146362f $X=0.36 $Y=0.036
c40 27 VSS 0.00325271f $X=0.342 $Y=0.036
c41 26 VSS 0.00146362f $X=0.306 $Y=0.036
c42 25 VSS 0.00287879f $X=0.288 $Y=0.036
c43 24 VSS 4.33098e-19 $X=0.256 $Y=0.036
c44 23 VSS 0.00312887f $X=0.252 $Y=0.036
c45 19 VSS 0.00234273f $X=0.216 $Y=0.036
c46 18 VSS 0.00164743f $X=0.216 $Y=0.036
c47 16 VSS 0.00628666f $X=0.396 $Y=0.036
c48 14 VSS 0.00169758f $X=0.376 $Y=0.216
c49 10 VSS 0.0022026f $X=0.27 $Y=0.216
c50 6 VSS 5.70405e-19 $X=0.287 $Y=0.216
c51 1 VSS 8.77547e-19 $X=0.233 $Y=0.0675
r52 47 48 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.164 $X2=0.405 $Y2=0.1765
r53 46 47 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.07 $X2=0.405 $Y2=0.164
r54 45 46 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.063 $X2=0.405 $Y2=0.07
r55 44 48 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.1765
r56 43 50 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.036
r57 43 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.063
r58 41 42 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.198 $X2=0.369 $Y2=0.198
r59 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r60 39 40 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.198 $X2=0.342 $Y2=0.198
r61 38 39 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.198 $X2=0.338 $Y2=0.198
r62 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.306 $Y2=0.198
r63 35 42 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.198 $X2=0.369 $Y2=0.198
r64 31 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.198 $X2=0.288 $Y2=0.198
r65 29 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.198 $X2=0.405 $Y2=0.189
r66 29 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.378 $Y2=0.198
r67 27 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r68 26 27 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.342 $Y2=0.036
r69 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r70 24 25 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.036 $X2=0.288 $Y2=0.036
r71 23 24 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.256 $Y2=0.036
r72 18 23 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.252 $Y2=0.036
r73 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r74 16 50 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.405 $Y2=0.036
r75 16 28 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.36 $Y2=0.036
r76 14 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.198 $X2=0.378
+ $Y2=0.198
r77 11 14 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.216 $X2=0.376 $Y2=0.216
r78 10 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.198 $X2=0.27
+ $Y2=0.198
r79 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.216 $X2=0.27 $Y2=0.216
r80 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.216 $X2=0.27 $Y2=0.216
r81 5 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r82 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r83 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./AOI33xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt AOI33xp33_ASAP7_75t_L  VSS VDD A1 A2 A3 B1 B2 B3 Y
* 
* Y	Y
* B3	B3
* B2	B2
* B1	B1
* A3	A3
* A2	A2
* A1	A1
M0 noxref_11 N_A1_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_12 N_A2_M1_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_A3_M2_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_13 N_B1_M3_g N_Y_M3_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_14 N_B2_M4_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 VSS N_B3_M5_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_9 N_A1_M6_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M7 VDD N_A2_M7_g noxref_9 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M8 noxref_9 N_A3_M8_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M9 N_Y_M9_d N_B1_M9_g noxref_9 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M10 noxref_9 N_B2_M10_g N_Y_M10_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.189
M11 N_Y_M11_d N_B3_M11_g noxref_9 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341
+ $Y=0.189
*
* 
* .include "AOI33xp33_ASAP7_75t_L.pex.sp.AOI33XP33_ASAP7_75T_L.pxi"
* BEGIN of "./AOI33xp33_ASAP7_75t_L.pex.sp.AOI33XP33_ASAP7_75T_L.pxi"
* File: AOI33xp33_ASAP7_75t_L.pex.sp.AOI33XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:17:02 2017
* 
x_PM_AOI33XP33_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M6_g A1 N_A1_c_3_p
+ N_A1_c_4_p VSS PM_AOI33XP33_ASAP7_75T_L%A1
x_PM_AOI33XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_10_n N_A2_M7_g N_A2_c_20_p
+ N_A2_c_11_n N_A2_c_12_n N_A2_c_13_n N_A2_c_25_p N_A2_c_26_p N_A2_c_21_p
+ N_A2_c_14_n N_A2_c_19_p A2 VSS PM_AOI33XP33_ASAP7_75T_L%A2
x_PM_AOI33XP33_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_35_n N_A3_M8_g N_A3_c_36_n
+ N_A3_c_37_n A3 N_A3_c_39_n VSS PM_AOI33XP33_ASAP7_75T_L%A3
x_PM_AOI33XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_51_n N_B1_M9_g B1 VSS
+ PM_AOI33XP33_ASAP7_75T_L%B1
x_PM_AOI33XP33_ASAP7_75T_L%B2 N_B2_M4_g N_B2_c_64_n N_B2_M10_g B2 VSS
+ PM_AOI33XP33_ASAP7_75T_L%B2
x_PM_AOI33XP33_ASAP7_75T_L%B3 N_B3_M5_g N_B3_c_76_n N_B3_M11_g B3 VSS
+ PM_AOI33XP33_ASAP7_75T_L%B3
x_PM_AOI33XP33_ASAP7_75T_L%Y N_Y_M3_s N_Y_M2_d N_Y_M10_s N_Y_M9_d N_Y_c_98_n
+ N_Y_M11_d N_Y_c_101_n N_Y_c_83_n N_Y_c_84_n N_Y_c_88_n N_Y_c_107_p N_Y_c_89_n
+ N_Y_c_108_p N_Y_c_93_n N_Y_c_85_n N_Y_c_91_n N_Y_c_106_n N_Y_c_95_n N_Y_c_97_n
+ Y VSS PM_AOI33XP33_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00328721f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_10_n 6.89019e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p N_A2_c_11_n 0.0017332f $X=0.027 $Y=0.135 $X2=0.027 $Y2=0.198
cc_4 N_A1_c_4_p N_A2_c_12_n 0.0017332f $X=0.063 $Y=0.135 $X2=0.064 $Y2=0.198
cc_5 N_A1_M0_g N_A2_c_13_n 4.2257e-19 $X=0.081 $Y=0.0675 $X2=0.09 $Y2=0.198
cc_6 A1 N_A2_c_14_n 6.80848e-19 $X=0.027 $Y=0.08 $X2=0.135 $Y2=0.135
cc_7 N_A1_c_4_p N_A2_c_14_n 0.0036144f $X=0.063 $Y=0.135 $X2=0.135 $Y2=0.135
cc_8 N_A1_M0_g N_A3_M2_g 2.48122e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_9 N_A2_M1_g N_A3_M2_g 0.00312021f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_10 N_A2_c_10_n N_A3_c_35_n 6.52245e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_11 N_A2_c_14_n N_A3_c_36_n 0.00117226f $X=0.135 $Y=0.135 $X2=0.018 $Y2=0.08
cc_12 N_A2_c_19_p N_A3_c_37_n 0.00117226f $X=0.135 $Y=0.1665 $X2=0 $Y2=0
cc_13 N_A2_c_20_p A3 0.00117226f $X=0.126 $Y=0.198 $X2=0 $Y2=0
cc_14 N_A2_c_21_p N_A3_c_39_n 0.00117226f $X=0.135 $Y=0.189 $X2=0.027 $Y2=0.135
cc_15 N_A2_M1_g N_B1_M3_g 2.53865e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_A2_c_14_n B1 6.71971e-19 $X=0.135 $Y=0.135 $X2=0.018 $Y2=0.08
cc_17 VSS N_A2_c_20_p 0.00101017f $X=0.126 $Y=0.198 $X2=0.081 $Y2=0.135
cc_18 VSS N_A2_c_25_p 7.27109e-19 $X=0.099 $Y=0.198 $X2=0.081 $Y2=0.135
cc_19 VSS N_A2_c_26_p 0.00171909f $X=0.1125 $Y=0.198 $X2=0.081 $Y2=0.135
cc_20 VSS N_A2_M1_g 2.35623e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_21 VSS N_A2_c_26_p 0.00402668f $X=0.1125 $Y=0.198 $X2=0 $Y2=0
cc_22 VSS A2 6.90371e-19 $X=0.024 $Y=0.233 $X2=0 $Y2=0
cc_23 N_A2_c_14_n N_Y_c_83_n 9.2243e-19 $X=0.135 $Y=0.135 $X2=0.027 $Y2=0.135
cc_24 N_A2_c_14_n N_Y_c_84_n 0.00134497f $X=0.135 $Y=0.135 $X2=0.063 $Y2=0.135
cc_25 VSS N_A2_c_14_n 3.86632e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_26 N_A3_M2_g N_B1_M3_g 0.00353416f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_27 N_A3_c_35_n N_B1_c_51_n 6.52245e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_28 N_A3_c_36_n B1 0.00253315f $X=0.189 $Y=0.135 $X2=0.018 $Y2=0.08
cc_29 N_A3_M2_g N_B2_M4_g 2.88628e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_30 VSS A3 0.00226216f $X=0.186 $Y=0.198 $X2=0.018 $Y2=0.126
cc_31 VSS N_A3_M2_g 2.38942e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_32 VSS A3 0.004203f $X=0.186 $Y=0.198 $X2=0.081 $Y2=0.135
cc_33 A3 N_Y_c_85_n 8.35736e-19 $X=0.186 $Y=0.198 $X2=0 $Y2=0
cc_34 N_B1_M3_g N_B2_M4_g 0.00355599f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_35 N_B1_c_51_n N_B2_c_64_n 6.52245e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_36 B1 B2 0.00487337f $X=0.238 $Y=0.115 $X2=0.018 $Y2=0.225
cc_37 N_B1_M3_g N_B3_M5_g 2.88628e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_38 VSS N_B1_M3_g 3.50057e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_39 VSS B1 5.3295e-19 $X=0.238 $Y=0.115 $X2=0 $Y2=0
cc_40 B1 N_Y_c_83_n 0.00422873f $X=0.238 $Y=0.115 $X2=0 $Y2=0
cc_41 B1 N_Y_c_84_n 0.00318534f $X=0.238 $Y=0.115 $X2=0 $Y2=0
cc_42 N_B1_M3_g N_Y_c_88_n 2.35623e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_43 N_B2_M4_g N_B3_M5_g 0.00353416f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_44 N_B2_c_64_n N_B3_c_76_n 6.86053e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_45 B2 B3 0.00498824f $X=0.303 $Y=0.122 $X2=0.189 $Y2=0.135
cc_46 VSS N_B2_M4_g 2.38942e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_B2_M4_g N_Y_c_89_n 3.49568e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_48 B2 N_Y_c_89_n 0.00124849f $X=0.303 $Y=0.122 $X2=0 $Y2=0
cc_49 N_B2_M4_g N_Y_c_91_n 2.79215e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_50 B2 N_Y_c_91_n 0.00123647f $X=0.303 $Y=0.122 $X2=0 $Y2=0
cc_51 N_B3_M5_g N_Y_c_93_n 2.65232e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_52 B3 N_Y_c_93_n 0.00124849f $X=0.353 $Y=0.122 $X2=0 $Y2=0
cc_53 N_B3_M5_g N_Y_c_95_n 3.54918e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_54 B3 N_Y_c_95_n 0.00121958f $X=0.353 $Y=0.122 $X2=0 $Y2=0
cc_55 B3 N_Y_c_97_n 0.00401351f $X=0.353 $Y=0.122 $X2=0 $Y2=0
cc_56 VSS N_Y_c_98_n 0.00288888f $X=0.216 $Y=0.216 $X2=0.018 $Y2=0.225
cc_57 VSS N_Y_c_98_n 0.00299929f $X=0.324 $Y=0.216 $X2=0.018 $Y2=0.225
cc_58 VSS N_Y_c_98_n 0.00250965f $X=0.324 $Y=0.234 $X2=0.018 $Y2=0.225
cc_59 VSS N_Y_c_101_n 0.00270623f $X=0.324 $Y=0.216 $X2=0.09 $Y2=0.198
cc_60 VSS N_Y_c_101_n 3.09693e-19 $X=0.324 $Y=0.234 $X2=0.09 $Y2=0.198
cc_61 VSS N_Y_c_84_n 7.80071e-19 $X=0.216 $Y=0.216 $X2=0 $Y2=0
cc_62 VSS N_Y_c_85_n 2.52562e-19 $X=0.216 $Y=0.216 $X2=0 $Y2=0
cc_63 VSS N_Y_c_85_n 0.0070243f $X=0.324 $Y=0.234 $X2=0 $Y2=0
cc_64 VSS N_Y_c_106_n 0.00365671f $X=0.324 $Y=0.216 $X2=0 $Y2=0
cc_65 VSS N_Y_c_107_p 4.20159e-19 $X=0.288 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_66 VSS N_Y_c_108_p 4.51936e-19 $X=0.342 $Y=0.036 $X2=0.135 $Y2=0.0675

* END of "./AOI33xp33_ASAP7_75t_L.pex.sp.AOI33XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: A2O1A1Ixp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 11:57:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "A2O1A1Ixp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./A2O1A1Ixp33_ASAP7_75t_L.pex.sp.pex"
* File: A2O1A1Ixp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 11:57:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_A2O1A1IXP33_ASAP7_75T_L%A1 2 5 7 14 17 19 20 24 VSS
c19 24 VSS 0.00553658f $X=0.018 $Y=0.135
c20 20 VSS 1.29148e-19 $X=0.0635 $Y=0.135
c21 19 VSS 0.00104753f $X=0.046 $Y=0.135
c22 17 VSS 5.51854e-19 $X=0.081 $Y=0.135
c23 14 VSS 0.00487907f $X=0.018 $Y=0.187
c24 5 VSS 0.00263014f $X=0.081 $Y=0.135
c25 2 VSS 0.0632929f $X=0.081 $Y=0.0675
r26 19 20 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r27 17 20 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r28 15 24 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r29 15 19 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.046 $Y2=0.135
r30 11 24 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r31 11 14 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.187
r32 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r33 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r34 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_A2O1A1IXP33_ASAP7_75T_L%A2 2 5 7 12 17 19 VSS
c18 19 VSS 2.14622e-20 $X=0.135 $Y=0.148
c19 17 VSS 0.00320123f $X=0.132 $Y=0.152
c20 12 VSS 0.00309788f $X=0.135 $Y=0.136
c21 5 VSS 0.00107247f $X=0.135 $Y=0.136
c22 2 VSS 0.0588446f $X=0.135 $Y=0.0675
r23 18 19 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.148
r24 17 19 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.152 $X2=0.135 $Y2=0.148
r25 12 18 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.136 $X2=0.135 $Y2=0.144
r26 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.136 $X2=0.135
+ $Y2=0.136
r27 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.136 $X2=0.135 $Y2=0.2025
r28 2 5 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.136
.ends

.subckt PM_A2O1A1IXP33_ASAP7_75T_L%B 2 5 7 12 19 21 VSS
c19 21 VSS 0.00151874f $X=0.189 $Y=0.115
c20 12 VSS 0.00146933f $X=0.189 $Y=0.136
c21 5 VSS 0.00107335f $X=0.189 $Y=0.136
c22 2 VSS 0.0617009f $X=0.189 $Y=0.054
r23 19 21 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.187
+ $Y=0.115 $X2=0.189 $Y2=0.115
r24 9 21 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.124 $X2=0.189 $Y2=0.115
r25 9 12 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.124 $X2=0.189 $Y2=0.136
r26 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.136 $X2=0.189
+ $Y2=0.136
r27 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.136 $X2=0.189 $Y2=0.2025
r28 2 5 307.213 $w=2e-08 $l=8.2e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.136
.ends

.subckt PM_A2O1A1IXP33_ASAP7_75T_L%C 2 5 7 11 13 16 VSS
c13 16 VSS 4.92608e-21 $X=0.297 $Y=0.13
c14 13 VSS 8.06259e-19 $X=0.297 $Y=0.136
c15 11 VSS 0.00208843f $X=0.296 $Y=0.083
c16 5 VSS 0.00170008f $X=0.297 $Y=0.136
c17 2 VSS 0.0661183f $X=0.297 $Y=0.0675
r18 15 16 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.124 $X2=0.297 $Y2=0.13
r19 13 16 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.136 $X2=0.297 $Y2=0.13
r20 11 15 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.083 $X2=0.297 $Y2=0.124
r21 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.136 $X2=0.297
+ $Y2=0.136
r22 5 7 299.72 $w=2e-08 $l=8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.136 $X2=0.297 $Y2=0.216
r23 2 5 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.136
.ends

.subckt PM_A2O1A1IXP33_ASAP7_75T_L%8 1 4 6 7 10 12 18 20 22 VSS
c16 23 VSS 9.96927e-19 $X=0.153 $Y=0.234
c17 22 VSS 0.0042362f $X=0.144 $Y=0.234
c18 21 VSS 0.00244569f $X=0.107 $Y=0.234
c19 20 VSS 0.00369061f $X=0.095 $Y=0.234
c20 18 VSS 0.00478328f $X=0.162 $Y=0.234
c21 12 VSS 0.00186838f $X=0.054 $Y=0.234
c22 10 VSS 0.00764745f $X=0.162 $Y=0.2025
c23 6 VSS 5.38922e-19 $X=0.179 $Y=0.2025
c24 4 VSS 0.00609725f $X=0.056 $Y=0.2025
c25 1 VSS 3.33606e-19 $X=0.071 $Y=0.2025
r26 22 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.153 $Y2=0.234
r27 21 22 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.234 $X2=0.144 $Y2=0.234
r28 20 21 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.234 $X2=0.107 $Y2=0.234
r29 18 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.153 $Y2=0.234
r30 12 20 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.095 $Y2=0.234
r31 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r32 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r33 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r34 4 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r35 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
.ends

.subckt PM_A2O1A1IXP33_ASAP7_75T_L%Y 1 6 11 14 21 22 23 26 30 32 VSS
c16 34 VSS 3.79545e-19 $X=0.351 $Y=0.2145
c17 33 VSS 3.69599e-19 $X=0.351 $Y=0.207
c18 32 VSS 0.00583981f $X=0.351 $Y=0.2
c19 31 VSS 8.85605e-19 $X=0.351 $Y=0.063
c20 30 VSS 5.0606e-19 $X=0.352 $Y=0.222
c21 26 VSS 0.00320547f $X=0.324 $Y=0.036
c22 23 VSS 0.00958109f $X=0.342 $Y=0.036
c23 22 VSS 0.00146498f $X=0.306 $Y=0.234
c24 21 VSS 0.00385745f $X=0.288 $Y=0.234
c25 16 VSS 0.00877172f $X=0.342 $Y=0.234
c26 14 VSS 0.0213714f $X=0.272 $Y=0.216
c27 11 VSS 2.6657e-19 $X=0.287 $Y=0.216
c28 9 VSS 4.25082e-19 $X=0.214 $Y=0.2025
c29 4 VSS 2.69461e-19 $X=0.322 $Y=0.0675
r30 33 34 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.207 $X2=0.351 $Y2=0.2145
r31 32 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.2 $X2=0.351 $Y2=0.207
r32 31 32 9.30247 $w=1.8e-08 $l=1.37e-07 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.063 $X2=0.351 $Y2=0.2
r33 30 34 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.222 $X2=0.351 $Y2=0.2145
r34 28 30 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.222
r35 27 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.063
r36 25 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r37 23 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.036 $X2=0.351 $Y2=0.045
r38 23 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.324 $Y2=0.036
r39 21 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r40 18 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.288 $Y2=0.234
r41 16 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.234 $X2=0.351 $Y2=0.225
r42 16 22 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.306 $Y2=0.234
r43 14 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r44 11 14 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.216 $X2=0.272 $Y2=0.216
r45 9 14 14.321 $w=8.1e-08 $l=5.6e-08 $layer=LISD $thickness=2.8e-08 $X=0.214
+ $Y=0.2025 $X2=0.27 $Y2=0.2025
r46 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.2025 $X2=0.214 $Y2=0.2025
r47 4 26 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r48 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends


* END of "./A2O1A1Ixp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt A2O1A1Ixp33_ASAP7_75t_L  VSS VDD A1 A2 B C Y
* 
* Y	Y
* C	C
* B	B
* A2	A2
* A1	A1
M0 noxref_10 N_A1_M0_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_A2_M1_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_7 N_B_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_C_M3_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M4 VDD N_A1_M4_g N_8_M4_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 N_8_M5_d N_A2_M5_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 N_Y_M6_d N_B_M6_g N_8_M6_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M7 VDD N_C_M7_g N_Y_M7_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287 $Y=0.189
*
* 
* .include "A2O1A1Ixp33_ASAP7_75t_L.pex.sp.A2O1A1IXP33_ASAP7_75T_L.pxi"
* BEGIN of "./A2O1A1Ixp33_ASAP7_75t_L.pex.sp.A2O1A1IXP33_ASAP7_75T_L.pxi"
* File: A2O1A1Ixp33_ASAP7_75t_L.pex.sp.A2O1A1IXP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 11:57:55 2017
* 
x_PM_A2O1A1IXP33_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M4_g A1 N_A1_c_3_p
+ N_A1_c_8_p N_A1_c_9_p N_A1_c_4_p VSS PM_A2O1A1IXP33_ASAP7_75T_L%A1
x_PM_A2O1A1IXP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_21_n N_A2_M5_g N_A2_c_22_n A2
+ N_A2_c_25_n VSS PM_A2O1A1IXP33_ASAP7_75T_L%A2
x_PM_A2O1A1IXP33_ASAP7_75T_L%B N_B_M2_g N_B_c_40_n N_B_M6_g N_B_c_41_n B
+ N_B_c_44_n VSS PM_A2O1A1IXP33_ASAP7_75T_L%B
x_PM_A2O1A1IXP33_ASAP7_75T_L%C N_C_M3_g N_C_c_58_n N_C_M7_g C N_C_c_62_p
+ N_C_c_60_n VSS PM_A2O1A1IXP33_ASAP7_75T_L%C
x_PM_A2O1A1IXP33_ASAP7_75T_L%8 N_8_M4_s N_8_c_70_n N_8_M6_s N_8_M5_d N_8_c_76_n
+ N_8_c_71_n N_8_c_80_n N_8_c_74_n N_8_c_77_n VSS PM_A2O1A1IXP33_ASAP7_75T_L%8
x_PM_A2O1A1IXP33_ASAP7_75T_L%Y N_Y_M3_d N_Y_M6_d N_Y_M7_s N_Y_c_86_n N_Y_c_101_n
+ N_Y_c_88_n N_Y_c_90_n N_Y_c_92_n Y N_Y_c_93_n VSS PM_A2O1A1IXP33_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00304756f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_21_n 0.00118189f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.136
cc_3 N_A1_c_3_p N_A2_c_22_n 8.78098e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.136
cc_4 N_A1_c_4_p N_A2_c_22_n 8.8451e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.136
cc_5 A1 A2 3.12618e-19 $X=0.018 $Y=0.187 $X2=0.132 $Y2=0.152
cc_6 A1 N_A2_c_25_n 4.6296e-19 $X=0.018 $Y=0.187 $X2=0.135 $Y2=0.148
cc_7 N_A1_M0_g N_B_M2_g 2.13359e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_8 VSS N_A1_c_8_p 3.04973e-19 $X=0.046 $Y=0.135 $X2=0.132 $Y2=0.152
cc_9 VSS N_A1_c_9_p 3.04973e-19 $X=0.0635 $Y=0.135 $X2=0.132 $Y2=0.152
cc_10 VSS N_A1_c_4_p 7.45434e-19 $X=0.018 $Y=0.135 $X2=0.132 $Y2=0.152
cc_11 VSS N_A1_c_4_p 0.0021283f $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.144
cc_12 VSS N_A1_M0_g 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_13 VSS N_A1_c_3_p 3.04973e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_14 A1 N_8_c_70_n 0.00201602f $X=0.018 $Y=0.187 $X2=0.135 $Y2=0.136
cc_15 A1 N_8_c_71_n 7.45434e-19 $X=0.018 $Y=0.187 $X2=0.135 $Y2=0.136
cc_16 N_A1_c_8_p N_8_c_71_n 3.04973e-19 $X=0.046 $Y=0.135 $X2=0.135 $Y2=0.136
cc_17 N_A1_c_9_p N_8_c_71_n 3.04973e-19 $X=0.0635 $Y=0.135 $X2=0.135 $Y2=0.136
cc_18 N_A1_M0_g N_8_c_74_n 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_19 N_A1_c_3_p N_8_c_74_n 3.04973e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_20 N_A2_M1_g N_B_M2_g 0.00304756f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_21 N_A2_c_21_n N_B_c_40_n 9.35653e-19 $X=0.135 $Y=0.136 $X2=0.081 $Y2=0.135
cc_22 N_A2_c_22_n N_B_c_41_n 0.00101107f $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_23 A2 N_B_c_41_n 0.00101107f $X=0.132 $Y=0.152 $X2=0 $Y2=0
cc_24 N_A2_c_25_n N_B_c_41_n 0.00101107f $X=0.135 $Y=0.148 $X2=0 $Y2=0
cc_25 N_A2_c_22_n N_B_c_44_n 0.00165689f $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_26 VSS N_A2_c_22_n 6.85004e-19 $X=0.135 $Y=0.136 $X2=0.081 $Y2=0.135
cc_27 VSS N_A2_M1_g 2.38524e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_28 VSS N_A2_c_22_n 0.00415914f $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_29 A2 N_8_c_76_n 0.00135883f $X=0.132 $Y=0.152 $X2=0 $Y2=0
cc_30 N_A2_M1_g N_8_c_77_n 2.34767e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_31 A2 N_8_c_77_n 0.00375078f $X=0.132 $Y=0.152 $X2=0 $Y2=0
cc_32 N_B_M2_g N_C_M3_g 2.82885e-19 $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.0675
cc_33 N_B_c_40_n N_C_c_58_n 5.73908e-19 $X=0.189 $Y=0.136 $X2=0.081 $Y2=0.135
cc_34 N_B_c_44_n C 0.00169053f $X=0.189 $Y=0.115 $X2=0.018 $Y2=0.144
cc_35 N_B_c_41_n N_C_c_60_n 7.59063e-19 $X=0.189 $Y=0.136 $X2=0.081 $Y2=0.135
cc_36 VSS N_B_c_44_n 0.00343225f $X=0.189 $Y=0.115 $X2=0.018 $Y2=0.187
cc_37 VSS N_B_c_44_n 0.00113066f $X=0.189 $Y=0.115 $X2=0 $Y2=0
cc_38 VSS N_B_M2_g 3.58121e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_39 VSS N_B_c_44_n 7.70781e-19 $X=0.189 $Y=0.115 $X2=0 $Y2=0
cc_40 N_B_c_41_n N_8_c_76_n 0.00135201f $X=0.189 $Y=0.136 $X2=0 $Y2=0
cc_41 N_B_M2_g N_8_c_80_n 2.58023e-19 $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.135
cc_42 N_B_c_41_n N_8_c_80_n 0.00231231f $X=0.189 $Y=0.136 $X2=0.081 $Y2=0.135
cc_43 N_B_c_41_n N_Y_c_86_n 0.00280707f $X=0.189 $Y=0.136 $X2=0.018 $Y2=0.187
cc_44 VSS C 0.00357219f $X=0.296 $Y=0.083 $X2=0 $Y2=0
cc_45 N_C_c_62_p N_Y_c_86_n 0.00137619f $X=0.297 $Y=0.136 $X2=0 $Y2=0
cc_46 N_C_M3_g N_Y_c_88_n 2.63936e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_C_c_62_p N_Y_c_88_n 0.0012541f $X=0.297 $Y=0.136 $X2=0 $Y2=0
cc_48 N_C_M3_g N_Y_c_90_n 2.37171e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_49 C N_Y_c_90_n 0.00264064f $X=0.296 $Y=0.083 $X2=0 $Y2=0
cc_50 C N_Y_c_92_n 0.00134376f $X=0.296 $Y=0.083 $X2=0 $Y2=0
cc_51 N_C_c_58_n N_Y_c_93_n 3.26679e-19 $X=0.297 $Y=0.136 $X2=0 $Y2=0
cc_52 C N_Y_c_93_n 0.00564195f $X=0.296 $Y=0.083 $X2=0 $Y2=0
cc_53 VSS N_8_c_70_n 0.00107739f $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.135
cc_54 VSS N_Y_c_86_n 0.00325693f $X=0.272 $Y=0.0675 $X2=0.018 $Y2=0.187
cc_55 VSS N_Y_c_90_n 0.00111196f $X=0.272 $Y=0.0675 $X2=0 $Y2=0
cc_56 VSS N_Y_c_90_n 5.50102e-19 $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_57 VSS N_Y_c_92_n 0.00408029f $X=0.272 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_8_c_76_n N_Y_c_86_n 0.00366257f $X=0.162 $Y=0.2025 $X2=0.018 $Y2=0.187
cc_59 N_8_c_80_n N_Y_c_86_n 5.63911e-19 $X=0.162 $Y=0.234 $X2=0.018 $Y2=0.187
cc_60 N_8_c_80_n N_Y_c_101_n 3.85189e-19 $X=0.162 $Y=0.234 $X2=0 $Y2=0

* END of "./A2O1A1Ixp33_ASAP7_75t_L.pex.sp.A2O1A1IXP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: A2O1A1O1Ixp25_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 11:58:20 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "A2O1A1O1Ixp25_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./A2O1A1O1Ixp25_ASAP7_75t_L.pex.sp.pex"
* File: A2O1A1O1Ixp25_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 11:58:20 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_A2O1A1O1IXP25_ASAP7_75T_L%A2 2 5 7 12 17 19 20 24 VSS
c19 24 VSS 0.00563078f $X=0.018 $Y=0.135
c20 20 VSS 1.29148e-19 $X=0.0635 $Y=0.135
c21 19 VSS 0.00104753f $X=0.046 $Y=0.135
c22 17 VSS 5.58361e-19 $X=0.081 $Y=0.135
c23 12 VSS 0.00487476f $X=0.018 $Y=0.082
c24 5 VSS 0.00271507f $X=0.081 $Y=0.135
c25 2 VSS 0.0632929f $X=0.081 $Y=0.0675
r26 19 20 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r27 17 20 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r28 15 24 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r29 15 19 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.046 $Y2=0.135
r30 10 24 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.135
r31 10 12 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.082
r32 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r33 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r34 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_A2O1A1O1IXP25_ASAP7_75T_L%A1 2 5 7 12 17 19 VSS
c17 19 VSS 3.26314e-19 $X=0.135 $Y=0.166
c18 17 VSS 0.00311793f $X=0.136 $Y=0.188
c19 12 VSS 0.00360143f $X=0.135 $Y=0.135
c20 5 VSS 0.00112843f $X=0.135 $Y=0.135
c21 2 VSS 0.0581466f $X=0.135 $Y=0.0675
r22 18 19 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.166
r23 17 19 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.188 $X2=0.135 $Y2=0.166
r24 12 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r25 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_A2O1A1O1IXP25_ASAP7_75T_L%B 2 5 7 10 14 VSS
c11 10 VSS 0.00104703f $X=0.189 $Y=0.135
c12 5 VSS 0.00119297f $X=0.189 $Y=0.135
c13 2 VSS 0.0579003f $X=0.189 $Y=0.0675
r14 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.154
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_A2O1A1O1IXP25_ASAP7_75T_L%C 2 5 7 10 15 VSS
c11 15 VSS 4.54256e-19 $X=0.243 $Y=0.135
c12 10 VSS 0.00240263f $X=0.242 $Y=0.119
c13 5 VSS 0.00222303f $X=0.243 $Y=0.135
c14 2 VSS 0.0616768f $X=0.243 $Y=0.0675
r15 10 15 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.119 $X2=0.243 $Y2=0.135
r16 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_A2O1A1O1IXP25_ASAP7_75T_L%D 2 7 17 19 20 30 VSS
c17 30 VSS 0.00545897f $X=0.35 $Y=0.136
c18 20 VSS 1.95978e-19 $X=0.392 $Y=0.136
c19 19 VSS 7.88734e-19 $X=0.386 $Y=0.136
c20 17 VSS 3.41901e-19 $X=0.405 $Y=0.136
c21 5 VSS 0.00387112f $X=0.405 $Y=0.135
c22 2 VSS 0.0673057f $X=0.405 $Y=0.0675
r23 19 20 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.386
+ $Y=0.136 $X2=0.392 $Y2=0.136
r24 17 20 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.136 $X2=0.392 $Y2=0.136
r25 15 30 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.136 $X2=0.351 $Y2=0.136
r26 15 19 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.136 $X2=0.386 $Y2=0.136
r27 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.136 $X2=0.405
+ $Y2=0.136
r28 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r29 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_A2O1A1O1IXP25_ASAP7_75T_L%Y 1 6 11 14 19 23 24 25 26 27 31 33 35 36
+ 37 43 VSS
c20 43 VSS 0.0016534f $X=0.45 $Y=0.19
c21 42 VSS 0.00154763f $X=0.459 $Y=0.19
c22 37 VSS 7.68871e-19 $X=0.459 $Y=0.145
c23 36 VSS 0.00263815f $X=0.459 $Y=0.127
c24 35 VSS 8.60367e-19 $X=0.459 $Y=0.081
c25 34 VSS 0.00108941f $X=0.459 $Y=0.063
c26 33 VSS 0.00336356f $X=0.46 $Y=0.045
c27 31 VSS 0.00160863f $X=0.459 $Y=0.181
c28 29 VSS 0.00222592f $X=0.4365 $Y=0.036
c29 28 VSS 0.00144627f $X=0.423 $Y=0.036
c30 27 VSS 0.00236097f $X=0.414 $Y=0.036
c31 26 VSS 0.00368782f $X=0.386 $Y=0.036
c32 25 VSS 0.00361856f $X=0.342 $Y=0.036
c33 24 VSS 0.00640137f $X=0.311 $Y=0.036
c34 23 VSS 0.00647799f $X=0.378 $Y=0.036
c35 19 VSS 0.00379642f $X=0.27 $Y=0.036
c36 16 VSS 0.00206701f $X=0.45 $Y=0.036
c37 14 VSS 0.00292697f $X=0.43 $Y=0.2025
c38 6 VSS 5.34579e-19 $X=0.395 $Y=0.0675
c39 4 VSS 3.25039e-19 $X=0.268 $Y=0.0675
r40 43 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.19 $X2=0.4545 $Y2=0.19
r41 42 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.19 $X2=0.4545 $Y2=0.19
r42 39 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.19 $X2=0.45 $Y2=0.19
r43 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.127 $X2=0.459 $Y2=0.145
r44 35 36 3.12346 $w=1.8e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.127
r45 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.063 $X2=0.459 $Y2=0.081
r46 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.063
r47 31 42 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.181 $X2=0.459 $Y2=0.19
r48 31 37 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.181 $X2=0.459 $Y2=0.145
r49 28 29 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.423
+ $Y=0.036 $X2=0.4365 $Y2=0.036
r50 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.423 $Y2=0.036
r51 26 27 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.386
+ $Y=0.036 $X2=0.414 $Y2=0.036
r52 24 25 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.036 $X2=0.342 $Y2=0.036
r53 22 26 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.386 $Y2=0.036
r54 22 25 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.342 $Y2=0.036
r55 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r56 18 24 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.311 $Y2=0.036
r57 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r58 16 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.459 $Y2=0.036
r59 16 29 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4365 $Y2=0.036
r60 14 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.19 $X2=0.432
+ $Y2=0.19
r61 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.43 $Y2=0.2025
r62 9 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r63 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r64 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r65 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.268 $Y2=0.0675
.ends


* END of "./A2O1A1O1Ixp25_ASAP7_75t_L.pex.sp.pex"
* 
.subckt A2O1A1O1Ixp25_ASAP7_75t_L  VSS VDD A2 A1 B C D Y
* 
* Y	Y
* D	D
* C	C
* B	B
* A1	A1
* A2	A2
M0 noxref_12 N_A2_M0_g noxref_8 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_A1_M1_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_8 N_B_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_C_M3_g noxref_8 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 VSS N_D_M4_g N_Y_M4_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M5 VDD N_A2_M5_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M6 noxref_9 N_A1_M6_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 noxref_10 N_B_M7_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M8 VDD N_C_M8_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M9 N_Y_M9_d N_D_M9_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
*
* 
* .include "A2O1A1O1Ixp25_ASAP7_75t_L.pex.sp.A2O1A1O1IXP25_ASAP7_75T_L.pxi"
* BEGIN of "./A2O1A1O1Ixp25_ASAP7_75t_L.pex.sp.A2O1A1O1IXP25_ASAP7_75T_L.pxi"
* File: A2O1A1O1Ixp25_ASAP7_75t_L.pex.sp.A2O1A1O1IXP25_ASAP7_75T_L.pxi
* Created: Tue Sep  5 11:58:20 2017
* 
x_PM_A2O1A1O1IXP25_ASAP7_75T_L%A2 N_A2_M0_g N_A2_c_2_p N_A2_M5_g A2 N_A2_c_4_p
+ N_A2_c_9_p N_A2_c_10_p N_A2_c_5_p VSS PM_A2O1A1O1IXP25_ASAP7_75T_L%A2
x_PM_A2O1A1O1IXP25_ASAP7_75T_L%A1 N_A1_M1_g N_A1_c_21_n N_A1_M6_g N_A1_c_22_n A1
+ N_A1_c_25_n VSS PM_A2O1A1O1IXP25_ASAP7_75T_L%A1
x_PM_A2O1A1O1IXP25_ASAP7_75T_L%B N_B_M2_g N_B_c_39_n N_B_M7_g N_B_c_40_n B VSS
+ PM_A2O1A1O1IXP25_ASAP7_75T_L%B
x_PM_A2O1A1O1IXP25_ASAP7_75T_L%C N_C_M3_g N_C_c_50_n N_C_M8_g C N_C_c_53_p VSS
+ PM_A2O1A1O1IXP25_ASAP7_75T_L%C
x_PM_A2O1A1O1IXP25_ASAP7_75T_L%D N_D_M4_g N_D_M9_g N_D_c_74_p N_D_c_62_p
+ N_D_c_70_p D VSS PM_A2O1A1O1IXP25_ASAP7_75T_L%D
x_PM_A2O1A1O1IXP25_ASAP7_75T_L%Y N_Y_M3_d N_Y_M4_s N_Y_M9_d N_Y_c_91_n
+ N_Y_c_76_n N_Y_c_78_n N_Y_c_90_n N_Y_c_79_n N_Y_c_80_n N_Y_c_82_n N_Y_c_84_n Y
+ N_Y_c_85_n N_Y_c_86_n N_Y_c_87_n N_Y_c_88_n VSS PM_A2O1A1O1IXP25_ASAP7_75T_L%Y
cc_1 N_A2_M0_g N_A1_M1_g 0.00304756f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A2_c_2_p N_A1_c_21_n 0.00120928f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A2 N_A1_c_22_n 8.7742e-19 $X=0.018 $Y=0.082 $X2=0.135 $Y2=0.135
cc_4 N_A2_c_4_p N_A1_c_22_n 8.78098e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_5 N_A2_c_5_p A1 3.41226e-19 $X=0.018 $Y=0.135 $X2=0.136 $Y2=0.188
cc_6 N_A2_c_5_p N_A1_c_25_n 4.69126e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.166
cc_7 N_A2_M0_g N_B_M2_g 2.13359e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_8 VSS A2 7.45434e-19 $X=0.018 $Y=0.082 $X2=0.135 $Y2=0.135
cc_9 VSS N_A2_c_9_p 3.04973e-19 $X=0.046 $Y=0.135 $X2=0.135 $Y2=0.135
cc_10 VSS N_A2_c_10_p 3.04973e-19 $X=0.0635 $Y=0.135 $X2=0.135 $Y2=0.135
cc_11 VSS A2 0.0021283f $X=0.018 $Y=0.082 $X2=0.135 $Y2=0.135
cc_12 VSS N_A2_M0_g 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_13 VSS N_A2_c_4_p 3.04973e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_14 VSS N_A2_c_5_p 0.00201307f $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.135
cc_15 VSS N_A2_c_9_p 3.04973e-19 $X=0.046 $Y=0.135 $X2=0.135 $Y2=0.135
cc_16 VSS N_A2_c_10_p 3.04973e-19 $X=0.0635 $Y=0.135 $X2=0.135 $Y2=0.135
cc_17 VSS N_A2_c_5_p 7.45434e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.135
cc_18 VSS N_A2_M0_g 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_19 VSS N_A2_c_4_p 3.04973e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_20 N_A1_M1_g N_B_M2_g 0.00299674f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_21 N_A1_c_21_n N_B_c_39_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 N_A1_c_22_n N_B_c_40_n 0.00378938f $X=0.135 $Y=0.135 $X2=0.018 $Y2=0.126
cc_23 N_A1_M1_g N_C_M3_g 2.42379e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_24 VSS N_A1_c_22_n 6.85228e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_25 VSS A1 2.06869e-19 $X=0.136 $Y=0.188 $X2=0 $Y2=0
cc_26 VSS N_A1_M1_g 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_27 VSS N_A1_c_22_n 0.0042365f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_28 VSS N_A1_c_25_n 0.00138171f $X=0.135 $Y=0.166 $X2=0.018 $Y2=0.126
cc_29 VSS N_A1_M1_g 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_30 VSS A1 0.00406043f $X=0.136 $Y=0.188 $X2=0 $Y2=0
cc_31 N_B_M2_g N_C_M3_g 0.00335986f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_32 N_B_c_39_n N_C_c_50_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_33 N_B_c_40_n C 0.00388834f $X=0.189 $Y=0.135 $X2=0.018 $Y2=0.126
cc_34 VSS N_B_M2_g 3.47199e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_35 VSS N_B_c_40_n 5.30079e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_36 VSS N_B_c_40_n 0.00114532f $X=0.189 $Y=0.135 $X2=0.018 $Y2=0.126
cc_37 VSS N_B_c_40_n 0.00114532f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_38 C D 0.00158134f $X=0.242 $Y=0.119 $X2=0 $Y2=0
cc_39 N_C_c_53_p D 2.9478e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_40 VSS C 0.00129165f $X=0.242 $Y=0.119 $X2=0.135 $Y2=0.166
cc_41 VSS C 0.00113861f $X=0.242 $Y=0.119 $X2=0.135 $Y2=0.135
cc_42 VSS N_C_M3_g 2.56935e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_43 VSS N_C_c_53_p 0.00123604f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_44 C N_Y_c_76_n 0.00130873f $X=0.242 $Y=0.119 $X2=0.135 $Y2=0.166
cc_45 VSS D 0.00163356f $X=0.35 $Y=0.136 $X2=0 $Y2=0
cc_46 VSS N_D_c_62_p 6.59338e-19 $X=0.386 $Y=0.136 $X2=0.135 $Y2=0.188
cc_47 VSS D 0.00468336f $X=0.35 $Y=0.136 $X2=0 $Y2=0
cc_48 D N_Y_c_76_n 7.11362e-19 $X=0.35 $Y=0.136 $X2=0.135 $Y2=0.166
cc_49 D N_Y_c_78_n 0.00258211f $X=0.35 $Y=0.136 $X2=0 $Y2=0
cc_50 D N_Y_c_79_n 4.50315e-19 $X=0.35 $Y=0.136 $X2=0 $Y2=0
cc_51 N_D_c_62_p N_Y_c_80_n 2.80503e-19 $X=0.386 $Y=0.136 $X2=0 $Y2=0
cc_52 D N_Y_c_80_n 0.0042362f $X=0.35 $Y=0.136 $X2=0 $Y2=0
cc_53 N_D_M4_g N_Y_c_82_n 4.08393e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_54 N_D_c_70_p N_Y_c_82_n 2.80503e-19 $X=0.392 $Y=0.136 $X2=0 $Y2=0
cc_55 D N_Y_c_84_n 4.50945e-19 $X=0.35 $Y=0.136 $X2=0 $Y2=0
cc_56 D N_Y_c_85_n 2.3791e-19 $X=0.35 $Y=0.136 $X2=0 $Y2=0
cc_57 D N_Y_c_86_n 5.24172e-19 $X=0.35 $Y=0.136 $X2=0 $Y2=0
cc_58 N_D_c_74_p N_Y_c_87_n 7.35052e-19 $X=0.405 $Y=0.136 $X2=0 $Y2=0
cc_59 D N_Y_c_88_n 2.47164e-19 $X=0.35 $Y=0.136 $X2=0 $Y2=0
cc_60 VSS N_Y_c_76_n 0.00286928f $X=0.216 $Y=0.036 $X2=0.046 $Y2=0.135
cc_61 VSS N_Y_c_90_n 7.1482e-19 $X=0.216 $Y=0.036 $X2=0.018 $Y2=0.135
cc_62 VSS N_Y_c_91_n 0.00378962f $X=0.38 $Y=0.2025 $X2=0.185 $Y2=0.154
cc_63 VSS N_Y_c_91_n 3.09692e-19 $X=0.378 $Y=0.234 $X2=0.185 $Y2=0.154
cc_64 VSS N_Y_c_78_n 0.00125584f $X=0.38 $Y=0.2025 $X2=0 $Y2=0
cc_65 VSS N_Y_c_90_n 2.60604e-19 $X=0.311 $Y=0.234 $X2=0 $Y2=0
cc_66 VSS N_Y_c_79_n 2.60604e-19 $X=0.36 $Y=0.234 $X2=0 $Y2=0

* END of "./A2O1A1O1Ixp25_ASAP7_75t_L.pex.sp.A2O1A1O1IXP25_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

