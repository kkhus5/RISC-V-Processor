* File: OA211x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:47:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA211x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA211x2_ASAP7_75t_L.pex.sp.pex"
* File: OA211x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:47:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA211X2_ASAP7_75T_L%A2 2 5 7 11 16 21 24 26 VSS
c14 26 VSS 0.00509824f $X=0.018 $Y=0.135
c15 24 VSS 2.25698e-19 $X=0.046 $Y=0.135
c16 23 VSS 0.00101227f $X=0.04 $Y=0.135
c17 21 VSS 4.44824e-19 $X=0.081 $Y=0.135
c18 16 VSS 5.51618e-19 $X=0.018 $Y=0.116
c19 11 VSS 0.00245719f $X=0.018 $Y=0.083
c20 9 VSS 5.16126e-19 $X=0.018 $Y=0.126
c21 5 VSS 0.00258444f $X=0.081 $Y=0.135
c22 2 VSS 0.0662757f $X=0.081 $Y=0.0675
r23 23 24 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.135 $X2=0.046 $Y2=0.135
r24 21 24 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.046 $Y2=0.135
r25 19 26 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r26 19 23 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.04 $Y2=0.135
r27 15 16 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.106 $X2=0.018 $Y2=0.116
r28 11 15 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.083 $X2=0.018 $Y2=0.106
r29 9 26 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.135
r30 9 16 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.116
r31 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r32 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r33 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA211X2_ASAP7_75T_L%A1 2 5 7 10 16 18 VSS
c17 18 VSS 2.03296e-19 $X=0.135 $Y=0.171
c18 16 VSS 6.5677e-19 $X=0.134 $Y=0.187
c19 10 VSS 4.62526e-19 $X=0.135 $Y=0.135
c20 5 VSS 0.00118075f $X=0.135 $Y=0.135
c21 2 VSS 0.0602081f $X=0.135 $Y=0.0675
r22 17 18 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.171
r23 16 18 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.187 $X2=0.135 $Y2=0.171
r24 10 17 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r25 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r26 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OA211X2_ASAP7_75T_L%B 2 5 7 10 14 VSS
c15 14 VSS 8.28011e-19 $X=0.188 $Y=0.148
c16 10 VSS 4.80806e-19 $X=0.189 $Y=0.135
c17 5 VSS 0.00110856f $X=0.189 $Y=0.135
c18 2 VSS 0.0589701f $X=0.189 $Y=0.0675
r19 10 14 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.148
r20 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r21 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2295
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA211X2_ASAP7_75T_L%C 2 5 7 10 VSS
c11 10 VSS 4.32501e-19 $X=0.241 $Y=0.123
c12 5 VSS 0.00107228f $X=0.243 $Y=0.135
c13 2 VSS 0.0581648f $X=0.243 $Y=0.0675
r14 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.123 $X2=0.243 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r16 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2295
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OA211X2_ASAP7_75T_L%7 2 7 10 13 15 17 18 21 22 25 27 28 32 34 42 45
+ 47 48 53 54 55 57 58 59 63 64 68 71 VSS
c46 73 VSS 3.58896e-19 $X=0.297 $Y=0.1765
c47 71 VSS 1.68016e-19 $X=0.297 $Y=0.12
c48 70 VSS 3.26038e-19 $X=0.297 $Y=0.106
c49 68 VSS 2.92217e-19 $X=0.297 $Y=0.134
c50 64 VSS 4.15825e-19 $X=0.252 $Y=0.198
c51 63 VSS 0.00375332f $X=0.288 $Y=0.198
c52 62 VSS 0.00111524f $X=0.243 $Y=0.225
c53 60 VSS 0.00381525f $X=0.286 $Y=0.072
c54 59 VSS 5.17397e-19 $X=0.252 $Y=0.072
c55 58 VSS 0.00176262f $X=0.234 $Y=0.072
c56 57 VSS 5.17397e-19 $X=0.198 $Y=0.072
c57 56 VSS 2.28963e-19 $X=0.18 $Y=0.072
c58 55 VSS 4.67884e-19 $X=0.176 $Y=0.072
c59 54 VSS 8.46035e-21 $X=0.144 $Y=0.072
c60 53 VSS 6.951e-19 $X=0.126 $Y=0.072
c61 48 VSS 5.71206e-20 $X=0.288 $Y=0.072
c62 47 VSS 0.00146362f $X=0.198 $Y=0.234
c63 46 VSS 0.00577713f $X=0.18 $Y=0.234
c64 45 VSS 0.00146362f $X=0.144 $Y=0.234
c65 44 VSS 0.00257933f $X=0.126 $Y=0.234
c66 43 VSS 9.36518e-19 $X=0.099 $Y=0.234
c67 42 VSS 0.00329977f $X=0.09 $Y=0.234
c68 34 VSS 0.00189006f $X=0.054 $Y=0.234
c69 32 VSS 0.00639545f $X=0.234 $Y=0.234
c70 31 VSS 0.00587039f $X=0.216 $Y=0.2295
c71 27 VSS 5.34547e-19 $X=0.233 $Y=0.2295
c72 25 VSS 0.00356808f $X=0.056 $Y=0.216
c73 22 VSS 2.6657e-19 $X=0.071 $Y=0.216
c74 21 VSS 0.00210789f $X=0.108 $Y=0.0675
c75 17 VSS 6.64001e-19 $X=0.125 $Y=0.0675
c76 13 VSS 0.00381033f $X=0.351 $Y=0.134
c77 10 VSS 0.0632947f $X=0.351 $Y=0.0675
c78 2 VSS 0.0597618f $X=0.297 $Y=0.0675
r79 72 73 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.164 $X2=0.297 $Y2=0.1765
r80 70 71 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.12
r81 68 72 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.134 $X2=0.297 $Y2=0.164
r82 68 71 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.134 $X2=0.297 $Y2=0.12
r83 66 73 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.1765
r84 65 70 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.081 $X2=0.297 $Y2=0.106
r85 63 66 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.198 $X2=0.297 $Y2=0.189
r86 63 64 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.252 $Y2=0.198
r87 61 64 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.243 $Y=0.207 $X2=0.252 $Y2=0.198
r88 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.207 $X2=0.243 $Y2=0.225
r89 59 60 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.072 $X2=0.286 $Y2=0.072
r90 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.252 $Y2=0.072
r91 57 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.072 $X2=0.234 $Y2=0.072
r92 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.072 $X2=0.198 $Y2=0.072
r93 55 56 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.072 $X2=0.18 $Y2=0.072
r94 54 55 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.176 $Y2=0.072
r95 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.144 $Y2=0.072
r96 50 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.126 $Y2=0.072
r97 48 65 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.072 $X2=0.297 $Y2=0.081
r98 48 60 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.286 $Y2=0.072
r99 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r100 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.18 $Y2=0.234
r101 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r102 43 44 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.234 $X2=0.126 $Y2=0.234
r103 42 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.099 $Y2=0.234
r104 40 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.198 $Y2=0.234
r105 34 42 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.09 $Y2=0.234
r106 32 62 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r107 32 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r108 31 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r109 28 31 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2295 $X2=0.216 $Y2=0.2295
r110 27 31 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2295 $X2=0.216 $Y2=0.2295
r111 25 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r112 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r113 21 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072
+ $X2=0.108 $Y2=0.072
r114 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r115 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r116 13 15 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.134 $X2=0.351 $Y2=0.2025
r117 10 13 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.134
r118 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.134 $X2=0.351 $Y2=0.134
r119 5 68 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.134 $X2=0.297
+ $Y2=0.134
r120 5 7 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.134 $X2=0.297 $Y2=0.2025
r121 2 5 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.134
.ends

.subckt PM_OA211X2_ASAP7_75T_L%Y 1 2 6 7 10 11 13 14 18 20 28 30 VSS
c18 30 VSS 0.0076332f $X=0.405 $Y=0.207
c19 29 VSS 8.85605e-19 $X=0.405 $Y=0.063
c20 28 VSS 8.85605e-19 $X=0.405 $Y=0.223
c21 20 VSS 0.00261875f $X=0.324 $Y=0.234
c22 18 VSS 0.0131443f $X=0.396 $Y=0.234
c23 14 VSS 0.0103019f $X=0.324 $Y=0.036
c24 13 VSS 0.0037985f $X=0.324 $Y=0.036
c25 11 VSS 0.013133f $X=0.396 $Y=0.036
c26 10 VSS 0.0103073f $X=0.324 $Y=0.2025
c27 6 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c28 1 VSS 5.38922e-19 $X=0.341 $Y=0.0675
r29 29 30 9.77778 $w=1.8e-08 $l=1.44e-07 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.063 $X2=0.405 $Y2=0.207
r30 28 30 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.223 $X2=0.405 $Y2=0.207
r31 26 28 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.223
r32 25 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.063
r33 18 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r34 18 20 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.324 $Y2=0.234
r35 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r36 11 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r37 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.324 $Y2=0.036
r38 10 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r39 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r40 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r41 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r42 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.324 $Y2=0.0675
r43 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.0675 $X2=0.324 $Y2=0.0675
.ends


* END of "./OA211x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA211x2_ASAP7_75t_L  VSS VDD A2 A1 B C Y
* 
* Y	Y
* C	C
* B	B
* A1	A1
* A2	A2
M0 N_7_M0_d N_A2_M0_g noxref_8 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_8 N_A1_M1_g N_7_M1_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_10 N_B_M2_g noxref_8 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_C_M3_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_7_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_7_M5_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 noxref_11 N_A2_M6_g N_7_M6_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M7 VDD N_A1_M7_g noxref_11 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M8 N_7_M8_d N_B_M8_g VDD VDD PMOS_LVT L=2e-08 W=2.7e-08 NFIN=1 $X=0.179 $Y=0.216
M9 VDD N_C_M9_g N_7_M9_s VDD PMOS_LVT L=2e-08 W=2.7e-08 NFIN=1 $X=0.233 $Y=0.216
M10 N_Y_M10_d N_7_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_Y_M11_d N_7_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "OA211x2_ASAP7_75t_L.pex.sp.OA211X2_ASAP7_75T_L.pxi"
* BEGIN of "./OA211x2_ASAP7_75t_L.pex.sp.OA211X2_ASAP7_75T_L.pxi"
* File: OA211x2_ASAP7_75t_L.pex.sp.OA211X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:47:18 2017
* 
x_PM_OA211X2_ASAP7_75T_L%A2 N_A2_M0_g N_A2_c_2_p N_A2_M6_g A2 N_A2_c_3_p
+ N_A2_c_4_p N_A2_c_9_p N_A2_c_5_p VSS PM_OA211X2_ASAP7_75T_L%A2
x_PM_OA211X2_ASAP7_75T_L%A1 N_A1_M1_g N_A1_c_16_n N_A1_M7_g N_A1_c_17_n A1
+ N_A1_c_20_n VSS PM_OA211X2_ASAP7_75T_L%A1
x_PM_OA211X2_ASAP7_75T_L%B N_B_M2_g N_B_c_34_n N_B_M8_g N_B_c_35_n B VSS
+ PM_OA211X2_ASAP7_75T_L%B
x_PM_OA211X2_ASAP7_75T_L%C N_C_M3_g N_C_c_49_n N_C_M9_g C VSS
+ PM_OA211X2_ASAP7_75T_L%C
x_PM_OA211X2_ASAP7_75T_L%7 N_7_M4_g N_7_M10_g N_7_M5_g N_7_c_74_n N_7_M11_g
+ N_7_M1_s N_7_M0_d N_7_c_79_p N_7_M6_s N_7_c_80_p N_7_M9_s N_7_M8_d N_7_c_99_p
+ N_7_c_58_n N_7_c_61_n N_7_c_62_n N_7_c_67_n N_7_c_93_p N_7_c_82_p N_7_c_64_n
+ N_7_c_84_p N_7_c_69_n N_7_c_103_p N_7_c_75_n N_7_c_100_p N_7_c_71_n N_7_c_89_p
+ N_7_c_78_n VSS PM_OA211X2_ASAP7_75T_L%7
x_PM_OA211X2_ASAP7_75T_L%Y N_Y_M5_d N_Y_M4_d N_Y_M11_d N_Y_M10_d N_Y_c_106_n
+ N_Y_c_108_n N_Y_c_109_n N_Y_c_112_n N_Y_c_114_n N_Y_c_115_n Y N_Y_c_119_n VSS
+ PM_OA211X2_ASAP7_75T_L%Y
cc_1 N_A2_M0_g N_A1_M1_g 0.00364065f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A2_c_2_p N_A1_c_16_n 9.88642e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A2_c_3_p N_A1_c_17_n 3.70126e-19 $X=0.018 $Y=0.116 $X2=0.135 $Y2=0.135
cc_4 N_A2_c_4_p N_A1_c_17_n 6.0497e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_5 N_A2_c_5_p A1 4.47736e-19 $X=0.018 $Y=0.135 $X2=0.134 $Y2=0.187
cc_6 N_A2_c_5_p N_A1_c_20_n 4.7353e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.171
cc_7 N_A2_M0_g N_B_M2_g 2.6588e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_8 N_A2_c_4_p N_7_c_58_n 4.05923e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_A2_c_9_p N_7_c_58_n 4.05923e-19 $X=0.046 $Y=0.135 $X2=0 $Y2=0
cc_10 N_A2_c_5_p N_7_c_58_n 3.17673e-19 $X=0.018 $Y=0.135 $X2=0 $Y2=0
cc_11 N_A2_M0_g N_7_c_61_n 4.01862e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_12 VSS A2 0.00146526f $X=0.018 $Y=0.083 $X2=0 $Y2=0
cc_13 VSS N_A2_M0_g 4.01862e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.171
cc_14 VSS N_A2_c_9_p 9.66105e-19 $X=0.046 $Y=0.135 $X2=0.135 $Y2=0.171
cc_15 N_A1_M1_g N_B_M2_g 0.0032267f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_A1_c_16_n N_B_c_34_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_17 N_A1_c_17_n N_B_c_35_n 0.00150681f $X=0.135 $Y=0.135 $X2=0.018 $Y2=0.083
cc_18 N_A1_c_17_n B 0.00150681f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_19 A1 B 0.00150681f $X=0.134 $Y=0.187 $X2=0 $Y2=0
cc_20 N_A1_M1_g N_C_M3_g 2.60137e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_21 N_A1_M1_g N_7_c_62_n 2.64276e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_22 A1 N_7_c_62_n 0.00124805f $X=0.134 $Y=0.187 $X2=0 $Y2=0
cc_23 N_A1_M1_g N_7_c_64_n 2.76185e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_24 N_A1_c_17_n N_7_c_64_n 0.0012322f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_25 VSS N_A1_M1_g 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0.018 $Y2=0.116
cc_26 N_B_M2_g N_C_M3_g 0.0033937f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_27 N_B_c_34_n N_C_c_49_n 8.88902e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_28 N_B_c_35_n C 0.00299705f $X=0.189 $Y=0.135 $X2=0.018 $Y2=0.083
cc_29 N_B_M2_g N_7_M4_g 2.25374e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_30 N_B_M2_g N_7_c_67_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_31 B N_7_c_67_n 0.00124805f $X=0.188 $Y=0.148 $X2=0 $Y2=0
cc_32 N_B_M2_g N_7_c_69_n 3.51973e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_33 N_B_c_35_n N_7_c_69_n 0.00121543f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_34 B N_7_c_71_n 6.96907e-19 $X=0.188 $Y=0.148 $X2=0 $Y2=0
cc_35 N_C_M3_g N_7_M4_g 0.00279092f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_36 N_C_M3_g N_7_M5_g 2.25374e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_37 N_C_c_49_n N_7_c_74_n 9.17673e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_38 N_C_M3_g N_7_c_75_n 3.51973e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_39 C N_7_c_75_n 0.00120437f $X=0.241 $Y=0.123 $X2=0 $Y2=0
cc_40 C N_7_c_71_n 0.00130733f $X=0.241 $Y=0.123 $X2=0 $Y2=0
cc_41 C N_7_c_78_n 0.00273632f $X=0.241 $Y=0.123 $X2=0 $Y2=0
cc_42 VSS N_7_c_79_p 0.00335635f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_43 VSS N_7_c_80_p 8.32391e-19 $X=0.056 $Y=0.216 $X2=0 $Y2=0
cc_44 VSS N_7_c_79_p 0.00189275f $X=0.108 $Y=0.0675 $X2=0.018 $Y2=0.116
cc_45 VSS N_7_c_82_p 0.00666759f $X=0.126 $Y=0.072 $X2=0.018 $Y2=0.116
cc_46 VSS N_7_c_79_p 0.00359732f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_47 VSS N_7_c_84_p 0.00262229f $X=0.176 $Y=0.072 $X2=0 $Y2=0
cc_48 VSS N_7_c_79_p 6.35113e-19 $X=0.108 $Y=0.0675 $X2=0.027 $Y2=0.135
cc_49 N_7_c_74_n N_Y_M5_d 3.87022e-19 $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.0675
cc_50 N_7_c_74_n N_Y_M11_d 3.7444e-19 $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.216
cc_51 N_7_c_74_n N_Y_c_106_n 7.60428e-19 $X=0.351 $Y=0.134 $X2=0.018 $Y2=0.083
cc_52 N_7_c_89_p N_Y_c_106_n 0.00160113f $X=0.297 $Y=0.134 $X2=0.018 $Y2=0.083
cc_53 N_7_M5_g N_Y_c_108_n 4.56718e-19 $X=0.351 $Y=0.0675 $X2=0.018 $Y2=0.083
cc_54 N_7_M4_g N_Y_c_109_n 2.34767e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_55 N_7_c_74_n N_Y_c_109_n 5.97402e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_56 N_7_c_93_p N_Y_c_109_n 0.00214292f $X=0.288 $Y=0.072 $X2=0 $Y2=0
cc_57 N_7_c_74_n N_Y_c_112_n 8.43851e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_58 N_7_c_93_p N_Y_c_112_n 0.00161003f $X=0.288 $Y=0.072 $X2=0 $Y2=0
cc_59 N_7_M5_g N_Y_c_114_n 4.61823e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_60 N_7_M4_g N_Y_c_115_n 2.63162e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_61 N_7_c_74_n N_Y_c_115_n 5.97991e-19 $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.135
cc_62 N_7_c_99_p N_Y_c_115_n 5.28228e-19 $X=0.234 $Y=0.234 $X2=0.081 $Y2=0.135
cc_63 N_7_c_100_p N_Y_c_115_n 9.14711e-19 $X=0.288 $Y=0.198 $X2=0.081 $Y2=0.135
cc_64 N_7_c_74_n N_Y_c_119_n 4.01182e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_65 N_7_c_93_p N_Y_c_119_n 0.00158346f $X=0.288 $Y=0.072 $X2=0 $Y2=0
cc_66 VSS N_7_c_103_p 4.30621e-19 $X=0.234 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_67 VSS N_Y_c_109_n 2.04426e-19 $X=0.162 $Y=0.036 $X2=0 $Y2=0

* END of "./OA211x2_ASAP7_75t_L.pex.sp.OA211X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA21x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:47:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA21x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA21x2_ASAP7_75t_L.pex.sp.pex"
* File: OA21x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:47:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA21X2_ASAP7_75T_L%A1 2 5 7 12 16 VSS
c15 16 VSS 0.00930798f $X=0.064 $Y=0.135
c16 12 VSS 0.0058019f $X=0.065 $Y=0.115
c17 5 VSS 0.00611424f $X=0.081 $Y=0.135
c18 2 VSS 0.06629f $X=0.081 $Y=0.0675
r19 16 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r20 12 16 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.115 $X2=0.064 $Y2=0.135
r21 5 17 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA21X2_ASAP7_75T_L%A2 2 5 7 10 13 VSS
c13 13 VSS 6.67386e-19 $X=0.135 $Y=0.135
c14 10 VSS 4.4801e-19 $X=0.134 $Y=0.121
c15 5 VSS 0.00124291f $X=0.135 $Y=0.135
c16 2 VSS 0.0614068f $X=0.135 $Y=0.0675
r17 10 13 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.121 $X2=0.135 $Y2=0.135
r18 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r19 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r20 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OA21X2_ASAP7_75T_L%B 2 5 7 11 14 VSS
c19 14 VSS 0.00229205f $X=0.189 $Y=0.135
c20 11 VSS 5.45659e-19 $X=0.193 $Y=0.115
c21 5 VSS 0.00155304f $X=0.189 $Y=0.135
c22 2 VSS 0.059622f $X=0.189 $Y=0.0675
r23 11 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r24 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r25 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r26 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA21X2_ASAP7_75T_L%6 2 7 10 13 15 17 18 21 22 23 26 27 32 33 35 37 38
+ 40 45 46 49 50 56 59 61 VSS
c47 61 VSS 3.5347e-19 $X=0.297 $Y=0.171
c48 59 VSS 1.94103e-19 $X=0.297 $Y=0.1205
c49 58 VSS 9.7335e-19 $X=0.297 $Y=0.106
c50 56 VSS 1.67689e-19 $X=0.297 $Y=0.135
c51 54 VSS 5.63105e-19 $X=0.297 $Y=0.189
c52 52 VSS 6.07985e-19 $X=0.256 $Y=0.198
c53 51 VSS 0.00110427f $X=0.239 $Y=0.198
c54 50 VSS 0.00119368f $X=0.224 $Y=0.198
c55 49 VSS 8.49048e-19 $X=0.288 $Y=0.198
c56 48 VSS 8.92485e-19 $X=0.215 $Y=0.225
c57 46 VSS 0.00105706f $X=0.193 $Y=0.234
c58 45 VSS 0.00364928f $X=0.18 $Y=0.234
c59 40 VSS 0.00475705f $X=0.206 $Y=0.234
c60 39 VSS 6.07985e-19 $X=0.256 $Y=0.072
c61 38 VSS 0.00370219f $X=0.239 $Y=0.072
c62 37 VSS 5.31938e-19 $X=0.198 $Y=0.072
c63 36 VSS 2.03739e-19 $X=0.18 $Y=0.072
c64 35 VSS 2.44387e-19 $X=0.176 $Y=0.072
c65 34 VSS 1.23838e-19 $X=0.148 $Y=0.072
c66 33 VSS 8.46035e-21 $X=0.144 $Y=0.072
c67 32 VSS 7.45119e-19 $X=0.126 $Y=0.072
c68 27 VSS 8.53644e-19 $X=0.288 $Y=0.072
c69 26 VSS 0.00746522f $X=0.162 $Y=0.2025
c70 22 VSS 6.48401e-19 $X=0.179 $Y=0.2025
c71 21 VSS 0.00241637f $X=0.108 $Y=0.0675
c72 17 VSS 6.411e-19 $X=0.125 $Y=0.0675
c73 13 VSS 0.00355466f $X=0.297 $Y=0.135
c74 10 VSS 0.0641602f $X=0.297 $Y=0.0675
c75 2 VSS 0.0615618f $X=0.243 $Y=0.0675
r76 60 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.153 $X2=0.297 $Y2=0.171
r77 58 59 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.1205
r78 56 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.153
r79 56 59 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.1205
r80 54 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.171
r81 53 58 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.081 $X2=0.297 $Y2=0.106
r82 51 52 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.239
+ $Y=0.198 $X2=0.256 $Y2=0.198
r83 50 51 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.224
+ $Y=0.198 $X2=0.239 $Y2=0.198
r84 49 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.198 $X2=0.297 $Y2=0.189
r85 49 52 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.256 $Y2=0.198
r86 47 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.215 $Y=0.207 $X2=0.224 $Y2=0.198
r87 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.215
+ $Y=0.207 $X2=0.215 $Y2=0.225
r88 45 46 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.193 $Y2=0.234
r89 42 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r90 40 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.206 $Y=0.234 $X2=0.215 $Y2=0.225
r91 40 46 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.206
+ $Y=0.234 $X2=0.193 $Y2=0.234
r92 38 39 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.239
+ $Y=0.072 $X2=0.256 $Y2=0.072
r93 37 38 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.072 $X2=0.239 $Y2=0.072
r94 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.072 $X2=0.198 $Y2=0.072
r95 35 36 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.072 $X2=0.18 $Y2=0.072
r96 34 35 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.072 $X2=0.176 $Y2=0.072
r97 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.148 $Y2=0.072
r98 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.144 $Y2=0.072
r99 29 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.126 $Y2=0.072
r100 27 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.072 $X2=0.297 $Y2=0.081
r101 27 39 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.256 $Y2=0.072
r102 26 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r103 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r104 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r105 21 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072
+ $X2=0.108 $Y2=0.072
r106 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r107 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r108 13 56 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r109 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.135 $X2=0.297 $Y2=0.2025
r110 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.0675 $X2=0.297 $Y2=0.135
r111 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r112 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r113 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OA21X2_ASAP7_75T_L%Y 1 2 6 7 10 14 16 23 28 30 VSS
c18 32 VSS 4.55454e-19 $X=0.351 $Y=0.216
c19 30 VSS 0.00177815f $X=0.351 $Y=0.102
c20 29 VSS 8.85605e-19 $X=0.351 $Y=0.063
c21 28 VSS 0.00474802f $X=0.352 $Y=0.141
c22 26 VSS 4.30151e-19 $X=0.351 $Y=0.225
c23 24 VSS 0.00305433f $X=0.324 $Y=0.234
c24 23 VSS 0.00474145f $X=0.306 $Y=0.234
c25 18 VSS 0.00620931f $X=0.342 $Y=0.234
c26 17 VSS 0.00305433f $X=0.324 $Y=0.036
c27 16 VSS 0.00496237f $X=0.306 $Y=0.036
c28 14 VSS 0.0104266f $X=0.27 $Y=0.036
c29 11 VSS 0.00620931f $X=0.342 $Y=0.036
c30 10 VSS 0.0101216f $X=0.27 $Y=0.2025
c31 6 VSS 6.41856e-19 $X=0.287 $Y=0.2025
c32 1 VSS 6.41856e-19 $X=0.287 $Y=0.0675
r33 31 32 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.207 $X2=0.351 $Y2=0.216
r34 29 30 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.063 $X2=0.351 $Y2=0.102
r35 28 31 4.48148 $w=1.8e-08 $l=6.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.141 $X2=0.351 $Y2=0.207
r36 28 30 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.141 $X2=0.351 $Y2=0.102
r37 26 32 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.216
r38 25 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.063
r39 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.324 $Y2=0.234
r40 20 23 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.306 $Y2=0.234
r41 18 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.234 $X2=0.351 $Y2=0.225
r42 18 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.324 $Y2=0.234
r43 16 17 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.324 $Y2=0.036
r44 13 16 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.306 $Y2=0.036
r45 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r46 11 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.036 $X2=0.351 $Y2=0.045
r47 11 17 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.324 $Y2=0.036
r48 10 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r49 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r50 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r51 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r52 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
r53 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends


* END of "./OA21x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA21x2_ASAP7_75t_L  VSS VDD A1 A2 B Y
* 
* Y	Y
* B	B
* A2	A2
* A1	A1
M0 N_6_M0_d N_A1_M0_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_7 N_A2_M1_g N_6_M1_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_B_M2_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_6_M3_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_6_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 noxref_9 N_A1_M5_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M6 N_6_M6_d N_A2_M6_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 VDD N_B_M7_g N_6_M7_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M8 N_Y_M8_d N_6_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M9 N_Y_M9_d N_6_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
*
* 
* .include "OA21x2_ASAP7_75t_L.pex.sp.OA21X2_ASAP7_75T_L.pxi"
* BEGIN of "./OA21x2_ASAP7_75t_L.pex.sp.OA21X2_ASAP7_75T_L.pxi"
* File: OA21x2_ASAP7_75t_L.pex.sp.OA21X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:47:41 2017
* 
x_PM_OA21X2_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M5_g A1 N_A1_c_9_p VSS
+ PM_OA21X2_ASAP7_75T_L%A1
x_PM_OA21X2_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_17_n N_A2_M6_g A2 N_A2_c_19_n VSS
+ PM_OA21X2_ASAP7_75T_L%A2
x_PM_OA21X2_ASAP7_75T_L%B N_B_M2_g N_B_c_31_n N_B_M7_g B N_B_c_34_p VSS
+ PM_OA21X2_ASAP7_75T_L%B
x_PM_OA21X2_ASAP7_75T_L%6 N_6_M3_g N_6_M8_g N_6_M4_g N_6_c_60_n N_6_M9_g
+ N_6_M1_s N_6_M0_d N_6_c_48_n N_6_M7_s N_6_M6_d N_6_c_49_n N_6_c_86_p
+ N_6_c_50_n N_6_c_54_n N_6_c_76_p N_6_c_62_n N_6_c_64_n N_6_c_65_n N_6_c_51_n
+ N_6_c_66_n N_6_c_83_p N_6_c_56_n N_6_c_93_p N_6_c_69_n N_6_c_70_n VSS
+ PM_OA21X2_ASAP7_75T_L%6
x_PM_OA21X2_ASAP7_75T_L%Y N_Y_M4_d N_Y_M3_d N_Y_M9_d N_Y_M8_d N_Y_c_95_n
+ N_Y_c_102_n N_Y_c_104_n N_Y_c_106_n Y N_Y_c_111_n VSS PM_OA21X2_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00361888f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_17_n 0.00106637f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A1 A2 0.00149415f $X=0.065 $Y=0.115 $X2=0.134 $Y2=0.121
cc_4 A1 N_A2_c_19_n 0.00149415f $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.135
cc_5 N_A1_M0_g N_B_M2_g 2.98169e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 A1 N_6_c_48_n 7.0658e-19 $X=0.065 $Y=0.115 $X2=0 $Y2=0
cc_7 A1 N_6_c_49_n 3.89749e-19 $X=0.065 $Y=0.115 $X2=0 $Y2=0
cc_8 A1 N_6_c_50_n 0.00129829f $X=0.065 $Y=0.115 $X2=0 $Y2=0
cc_9 N_A1_c_9_p N_6_c_51_n 5.30907e-19 $X=0.064 $Y=0.135 $X2=0 $Y2=0
cc_10 VSS A1 2.11432e-19 $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_11 VSS N_A1_c_2_p 4.0003e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_12 VSS A1 0.00353122f $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.135
cc_13 VSS A1 0.00324399f $X=0.065 $Y=0.115 $X2=0 $Y2=0
cc_14 VSS N_A1_M0_g 2.39633e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_15 VSS N_A1_c_2_p 3.09341e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_16 N_A2_M1_g N_B_M2_g 0.00354623f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 N_A2_c_17_n N_B_c_31_n 9.06722e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_18 A2 B 0.00309704f $X=0.134 $Y=0.121 $X2=0.064 $Y2=0.115
cc_19 N_A2_M1_g N_6_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_20 A2 N_6_c_49_n 0.00145684f $X=0.134 $Y=0.121 $X2=0.081 $Y2=0.135
cc_21 N_A2_M1_g N_6_c_54_n 2.76185e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_22 A2 N_6_c_54_n 0.0012322f $X=0.134 $Y=0.121 $X2=0 $Y2=0
cc_23 N_A2_c_19_n N_6_c_56_n 2.02524e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_24 VSS N_A2_M1_g 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0.064 $Y2=0.135
cc_25 N_B_M2_g N_6_M3_g 0.00287079f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_26 N_B_c_34_p N_6_M3_g 2.98947e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_27 N_B_M2_g N_6_M4_g 2.34385e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_28 N_B_c_31_n N_6_c_60_n 0.00122083f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_29 N_B_c_34_p N_6_c_49_n 2.79734e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_30 N_B_M2_g N_6_c_62_n 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_31 B N_6_c_62_n 0.00122403f $X=0.193 $Y=0.115 $X2=0 $Y2=0
cc_32 N_B_c_34_p N_6_c_64_n 8.51968e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_33 N_B_c_34_p N_6_c_65_n 4.77538e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_34 N_B_M2_g N_6_c_66_n 2.4825e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_B_c_34_p N_6_c_66_n 4.77538e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_36 N_B_c_34_p N_6_c_56_n 0.00293653f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_37 B N_6_c_69_n 6.8968e-19 $X=0.193 $Y=0.115 $X2=0 $Y2=0
cc_38 N_B_c_34_p N_6_c_70_n 5.51828e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_39 N_B_c_34_p N_Y_c_95_n 2.19213e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_40 VSS N_6_c_48_n 0.00391978f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_41 VSS N_6_c_48_n 0.00189275f $X=0.108 $Y=0.0675 $X2=0.064 $Y2=0.135
cc_42 VSS N_6_c_50_n 0.00666757f $X=0.126 $Y=0.072 $X2=0.064 $Y2=0.135
cc_43 VSS N_6_c_48_n 0.00352055f $X=0.108 $Y=0.0675 $X2=0.064 $Y2=0.135
cc_44 VSS N_6_c_49_n 0.00138157f $X=0.162 $Y=0.2025 $X2=0.064 $Y2=0.135
cc_45 VSS N_6_c_76_p 0.00233206f $X=0.176 $Y=0.072 $X2=0.064 $Y2=0.135
cc_46 VSS N_6_M1_s 2.09551e-19 $X=0.125 $Y=0.0675 $X2=0 $Y2=0
cc_47 VSS N_6_c_48_n 6.2062e-19 $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_48 N_6_c_60_n N_Y_M4_d 3.80246e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_49 N_6_c_60_n N_Y_M9_d 3.80246e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_50 N_6_c_60_n N_Y_c_95_n 8.00061e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_51 N_6_c_49_n N_Y_c_95_n 2.03108e-19 $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_52 N_6_c_83_p N_Y_c_95_n 0.00193825f $X=0.288 $Y=0.198 $X2=0 $Y2=0
cc_53 N_6_c_70_n N_Y_c_95_n 2.93295e-19 $X=0.297 $Y=0.171 $X2=0 $Y2=0
cc_54 N_6_c_60_n N_Y_c_102_n 8.00061e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_55 N_6_c_86_p N_Y_c_102_n 0.00193825f $X=0.288 $Y=0.072 $X2=0 $Y2=0
cc_56 N_6_M4_g N_Y_c_104_n 2.34993e-19 $X=0.297 $Y=0.0675 $X2=0.064 $Y2=0.135
cc_57 N_6_c_86_p N_Y_c_104_n 0.00444012f $X=0.288 $Y=0.072 $X2=0.064 $Y2=0.135
cc_58 N_6_M4_g N_Y_c_106_n 2.34993e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_59 N_6_c_65_n N_Y_c_106_n 8.87186e-19 $X=0.206 $Y=0.234 $X2=0 $Y2=0
cc_60 N_6_c_83_p N_Y_c_106_n 0.00410725f $X=0.288 $Y=0.198 $X2=0 $Y2=0
cc_61 N_6_c_60_n Y 3.32221e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_62 N_6_c_93_p Y 0.00274805f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_63 N_6_c_86_p N_Y_c_111_n 0.00274805f $X=0.288 $Y=0.072 $X2=0 $Y2=0
cc_64 VSS N_Y_c_104_n 2.88175e-19 $X=0.162 $Y=0.036 $X2=0.064 $Y2=0.135

* END of "./OA21x2_ASAP7_75t_L.pex.sp.OA21X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA221x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:48:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA221x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA221x2_ASAP7_75t_L.pex.sp.pex"
* File: OA221x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:48:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA221X2_ASAP7_75T_L%3 1 2 6 11 14 17 19 21 22 25 26 29 31 34 36 39 42
+ 43 44 46 50 51 52 53 54 55 56 57 61 62 63 65 66 72 73 77 78 79 81 86 VSS
c87 87 VSS 4.63222e-19 $X=0.144 $Y=0.135
c88 86 VSS 9.66734e-19 $X=0.153 $Y=0.135
c89 81 VSS 3.27401e-19 $X=0.135 $Y=0.135
c90 79 VSS 8.14173e-19 $X=0.837 $Y=0.207
c91 78 VSS 0.00356595f $X=0.837 $Y=0.189
c92 77 VSS 7.61702e-19 $X=0.837 $Y=0.117
c93 76 VSS 8.85605e-19 $X=0.837 $Y=0.099
c94 75 VSS 9.23055e-19 $X=0.837 $Y=0.225
c95 73 VSS 5.93175e-19 $X=0.824 $Y=0.072
c96 67 VSS 0.00220535f $X=0.828 $Y=0.072
c97 66 VSS 0.00319915f $X=0.7925 $Y=0.234
c98 65 VSS 0.00287092f $X=0.757 $Y=0.234
c99 64 VSS 0.00842861f $X=0.72 $Y=0.234
c100 63 VSS 0.00622549f $X=0.668 $Y=0.234
c101 62 VSS 0.00313021f $X=0.63 $Y=0.234
c102 61 VSS 0.00560798f $X=0.593 $Y=0.234
c103 57 VSS 8.6677e-19 $X=0.531 $Y=0.234
c104 56 VSS 0.00301945f $X=0.522 $Y=0.234
c105 55 VSS 0.010266f $X=0.485 $Y=0.234
c106 54 VSS 0.00301945f $X=0.379 $Y=0.234
c107 53 VSS 0.00832583f $X=0.342 $Y=0.234
c108 52 VSS 0.00278303f $X=0.252 $Y=0.234
c109 51 VSS 0.00112093f $X=0.215 $Y=0.234
c110 50 VSS 0.00445798f $X=0.202 $Y=0.234
c111 46 VSS 0.00270205f $X=0.162 $Y=0.234
c112 45 VSS 0.00687786f $X=0.828 $Y=0.234
c113 44 VSS 5.01276e-19 $X=0.153 $Y=0.207
c114 43 VSS 0.00158716f $X=0.153 $Y=0.189
c115 42 VSS 0.00126427f $X=0.153 $Y=0.225
c116 39 VSS 0.0062255f $X=0.754 $Y=0.216
c117 34 VSS 0.00361472f $X=0.542 $Y=0.2025
c118 31 VSS 4.59792e-19 $X=0.557 $Y=0.2025
c119 29 VSS 0.0031663f $X=0.322 $Y=0.2025
c120 25 VSS 0.0027496f $X=0.756 $Y=0.0675
c121 21 VSS 5.95149e-19 $X=0.773 $Y=0.0675
c122 17 VSS 0.00441776f $X=0.135 $Y=0.135
c123 14 VSS 0.0590374f $X=0.135 $Y=0.0675
c124 6 VSS 0.06187f $X=0.081 $Y=0.0675
c125 2 VSS 1.98976e-19 $X=0.336 $Y=0.174
c126 1 VSS 0.158442f $X=0.528 $Y=0.174
r127 87 88 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.1485 $Y2=0.135
r128 86 88 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.135 $X2=0.1485 $Y2=0.135
r129 81 87 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.144 $Y2=0.135
r130 78 79 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.189 $X2=0.837 $Y2=0.207
r131 77 78 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.117 $X2=0.837 $Y2=0.189
r132 76 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.117
r133 75 79 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.207
r134 74 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.081 $X2=0.837 $Y2=0.099
r135 72 73 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.757
+ $Y=0.072 $X2=0.824 $Y2=0.072
r136 69 72 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.072 $X2=0.757 $Y2=0.072
r137 67 74 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.072 $X2=0.837 $Y2=0.081
r138 67 73 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.072 $X2=0.824 $Y2=0.072
r139 65 66 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.757
+ $Y=0.234 $X2=0.7925 $Y2=0.234
r140 63 64 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.668
+ $Y=0.234 $X2=0.72 $Y2=0.234
r141 62 63 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.234 $X2=0.668 $Y2=0.234
r142 61 62 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.593
+ $Y=0.234 $X2=0.63 $Y2=0.234
r143 59 65 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.757 $Y2=0.234
r144 59 64 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.72 $Y2=0.234
r145 56 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.234 $X2=0.531 $Y2=0.234
r146 55 56 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.485
+ $Y=0.234 $X2=0.522 $Y2=0.234
r147 54 55 7.19753 $w=1.8e-08 $l=1.06e-07 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.234 $X2=0.485 $Y2=0.234
r148 53 54 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.379 $Y2=0.234
r149 52 53 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.342 $Y2=0.234
r150 51 52 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.215
+ $Y=0.234 $X2=0.252 $Y2=0.234
r151 50 51 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.234 $X2=0.215 $Y2=0.234
r152 48 61 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.593 $Y2=0.234
r153 48 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.531 $Y2=0.234
r154 46 50 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.202 $Y2=0.234
r155 45 75 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r156 45 66 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.7925 $Y2=0.234
r157 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.189 $X2=0.153 $Y2=0.207
r158 42 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.153 $Y=0.225 $X2=0.162 $Y2=0.234
r159 42 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.225 $X2=0.153 $Y2=0.207
r160 41 86 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.144 $X2=0.153 $Y2=0.135
r161 41 43 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.144 $X2=0.153 $Y2=0.189
r162 39 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234
+ $X2=0.756 $Y2=0.234
r163 36 39 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.216 $X2=0.754 $Y2=0.216
r164 34 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r165 31 34 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.542 $Y2=0.2025
r166 26 29 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.322 $Y2=0.2025
r167 25 69 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.072
+ $X2=0.756 $Y2=0.072
r168 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.756 $Y2=0.0675
r169 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.756 $Y2=0.0675
r170 17 81 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r171 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r172 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r173 9 17 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r174 9 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r175 6 9 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
r176 4 34 14.2411 $w=2.4e-08 $l=1.65e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.186 $X2=0.54 $Y2=0.2025
r177 3 29 14.2411 $w=2.4e-08 $l=1.65e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.186 $X2=0.324 $Y2=0.2025
r178 2 3 11.5737 $w=2.4e-08 $l=1.69706e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.336 $Y=0.174 $X2=0.324 $Y2=0.186
r179 1 4 11.5737 $w=2.4e-08 $l=1.69706e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.528 $Y=0.174 $X2=0.54 $Y2=0.186
r180 1 2 165.714 $w=2.4e-08 $l=1.92e-07 $layer=LISD $thickness=2.8e-08 $X=0.528
+ $Y=0.174 $X2=0.336 $Y2=0.174
.ends

.subckt PM_OA221X2_ASAP7_75T_L%A1 2 7 10 13 18 23 VSS
c25 23 VSS 4.55298e-19 $X=0.248 $Y=0.149
c26 18 VSS 0.00219659f $X=0.243 $Y=0.135
c27 13 VSS 0.00348524f $X=0.243 $Y=0.135
c28 10 VSS 0.0594912f $X=0.243 $Y=0.0675
c29 2 VSS 0.0587296f $X=0.189 $Y=0.0675
r30 18 23 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.149
r31 13 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r32 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r33 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r34 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r35 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA221X2_ASAP7_75T_L%A2 2 7 10 13 18 21 VSS
c24 21 VSS 5.91336e-19 $X=0.353 $Y=0.151
c25 18 VSS 0.00222665f $X=0.351 $Y=0.135
c26 13 VSS 0.00437597f $X=0.351 $Y=0.135
c27 10 VSS 0.0630057f $X=0.351 $Y=0.0675
c28 2 VSS 0.0598587f $X=0.297 $Y=0.0675
r29 18 21 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.151
r30 13 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r31 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r32 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r33 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r34 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OA221X2_ASAP7_75T_L%B2 2 8 11 13 18 21 VSS
c27 21 VSS 5.91336e-19 $X=0.511 $Y=0.151
c28 18 VSS 0.00141245f $X=0.513 $Y=0.135
c29 11 VSS 0.00423146f $X=0.567 $Y=0.135
c30 8 VSS 0.0610308f $X=0.567 $Y=0.0675
c31 2 VSS 0.0644501f $X=0.513 $Y=0.0675
r32 18 21 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.151
r33 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r34 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r35 5 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r36 5 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r37 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OA221X2_ASAP7_75T_L%B1 2 7 10 13 18 21 VSS
c28 21 VSS 8.68036e-19 $X=0.622 $Y=0.151
c29 18 VSS 0.00209539f $X=0.621 $Y=0.135
c30 13 VSS 0.00674707f $X=0.675 $Y=0.135
c31 10 VSS 0.0641433f $X=0.675 $Y=0.0675
c32 2 VSS 0.060715f $X=0.621 $Y=0.0675
r33 18 21 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.151
r34 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0675 $X2=0.675 $Y2=0.135
r35 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621
+ $Y=0.135 $X2=0.675 $Y2=0.135
r36 5 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r37 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r38 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
.ends

.subckt PM_OA221X2_ASAP7_75T_L%C 2 7 10 13 18 21 VSS
c26 21 VSS 9.46463e-19 $X=0.733 $Y=0.151
c27 18 VSS 0.00121581f $X=0.729 $Y=0.135
c28 13 VSS 0.00381291f $X=0.783 $Y=0.135
c29 10 VSS 0.0656485f $X=0.783 $Y=0.0675
c30 2 VSS 0.0596856f $X=0.729 $Y=0.0675
r31 18 21 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.135 $X2=0.729 $Y2=0.151
r32 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0675 $X2=0.783 $Y2=0.135
r33 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.135 $X2=0.783 $Y2=0.135
r34 5 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.729 $Y=0.135 $X2=0.729
+ $Y2=0.135
r35 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.135 $X2=0.729 $Y2=0.216
r36 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0675 $X2=0.729 $Y2=0.135
.ends

.subckt PM_OA221X2_ASAP7_75T_L%Y 1 2 6 7 10 14 19 20 26 28 32 41 VSS
c16 41 VSS 0.00144832f $X=0.108 $Y=0.216
c17 35 VSS 0.00230208f $X=0.0805 $Y=0.234
c18 34 VSS 0.00605721f $X=0.062 $Y=0.234
c19 33 VSS 0.00319807f $X=0.027 $Y=0.234
c20 32 VSS 0.00368818f $X=0.099 $Y=0.234
c21 28 VSS 0.00277412f $X=0.085 $Y=0.036
c22 27 VSS 0.00605721f $X=0.062 $Y=0.036
c23 26 VSS 0.00922845f $X=0.108 $Y=0.036
c24 25 VSS 0.00446698f $X=0.108 $Y=0.036
c25 23 VSS 0.00320021f $X=0.027 $Y=0.036
c26 22 VSS 3.21881e-19 $X=0.018 $Y=0.216
c27 20 VSS 8.11473e-19 $X=0.018 $Y=0.144
c28 19 VSS 6.07641e-19 $X=0.018 $Y=0.126
c29 18 VSS 0.0012055f $X=0.018 $Y=0.117
c30 17 VSS 0.00119129f $X=0.018 $Y=0.099
c31 16 VSS 0.00101662f $X=0.018 $Y=0.081
c32 15 VSS 8.29409e-19 $X=0.018 $Y=0.063
c33 14 VSS 0.00323297f $X=0.018 $Y=0.189
c34 12 VSS 3.03999e-19 $X=0.018 $Y=0.225
c35 10 VSS 0.0106335f $X=0.108 $Y=0.2025
c36 6 VSS 5.945e-19 $X=0.125 $Y=0.2025
c37 1 VSS 5.58795e-19 $X=0.125 $Y=0.0675
r38 39 41 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.225 $X2=0.108 $Y2=0.216
r39 34 35 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.062
+ $Y=0.234 $X2=0.0805 $Y2=0.234
r40 33 34 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.062 $Y2=0.234
r41 32 39 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.099 $Y=0.234 $X2=0.108 $Y2=0.225
r42 32 35 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.234 $X2=0.0805 $Y2=0.234
r43 27 28 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.062
+ $Y=0.036 $X2=0.085 $Y2=0.036
r44 25 28 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.085 $Y2=0.036
r45 25 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r46 23 27 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.062 $Y2=0.036
r47 21 22 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.207 $X2=0.018 $Y2=0.216
r48 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.144
r49 18 19 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.117 $X2=0.018 $Y2=0.126
r50 17 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.099 $X2=0.018 $Y2=0.117
r51 16 17 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.099
r52 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.081
r53 14 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.207
r54 14 20 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.144
r55 12 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r56 12 22 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.216
r57 11 23 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r58 11 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r59 10 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.216 $X2=0.108
+ $Y2=0.216
r60 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r61 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r62 5 26 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r63 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r64 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OA221x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA221x2_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 C Y
* 
* Y	Y
* C	C
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_10 N_A1_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_10 N_A1_M3_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_10 N_A2_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_10 N_A2_M5_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_10 N_B2_M6_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M7 noxref_10 N_B2_M7_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M8 noxref_10 N_B1_M8_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M9 noxref_10 N_B1_M9_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M10 N_3_M10_d N_C_M10_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M11 N_3_M11_d N_C_M11_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.027
M12 N_Y_M12_d N_3_M12_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M13 N_Y_M13_d N_3_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M14 noxref_12 N_A1_M14_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M15 N_3_M15_d N_A2_M15_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M16 noxref_13 N_B2_M16_g N_3_M16_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M17 VDD N_B1_M17_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M18 N_3_M18_d N_C_M18_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.719
+ $Y=0.189
*
* 
* .include "OA221x2_ASAP7_75t_L.pex.sp.OA221X2_ASAP7_75T_L.pxi"
* BEGIN of "./OA221x2_ASAP7_75t_L.pex.sp.OA221X2_ASAP7_75T_L.pxi"
* File: OA221x2_ASAP7_75t_L.pex.sp.OA221X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:48:03 2017
* 
x_PM_OA221X2_ASAP7_75T_L%3 N_3_c_12_p N_3_c_14_p N_3_M0_g N_3_M12_g N_3_M1_g
+ N_3_c_5_p N_3_M13_g N_3_M11_d N_3_M10_d N_3_c_38_p N_3_M15_d N_3_c_17_p
+ N_3_M16_s N_3_c_26_p N_3_M18_d N_3_c_39_p N_3_c_63_p N_3_c_7_p N_3_c_9_p
+ N_3_c_60_p N_3_c_3_p N_3_c_67_p N_3_c_10_p N_3_c_11_p N_3_c_13_p N_3_c_69_p
+ N_3_c_21_p N_3_c_24_p N_3_c_22_p N_3_c_29_p N_3_c_30_p N_3_c_34_p N_3_c_35_p
+ N_3_c_44_p N_3_c_36_p N_3_c_45_p N_3_c_42_p N_3_c_49_p N_3_c_56_p N_3_c_8_p
+ VSS PM_OA221X2_ASAP7_75T_L%3
x_PM_OA221X2_ASAP7_75T_L%A1 N_A1_M2_g N_A1_M14_g N_A1_M3_g N_A1_c_92_n
+ N_A1_c_94_n A1 VSS PM_OA221X2_ASAP7_75T_L%A1
x_PM_OA221X2_ASAP7_75T_L%A2 N_A2_M4_g N_A2_M15_g N_A2_M5_g N_A2_c_116_n
+ N_A2_c_118_n A2 VSS PM_OA221X2_ASAP7_75T_L%A2
x_PM_OA221X2_ASAP7_75T_L%B2 N_B2_M6_g N_B2_M7_g N_B2_c_140_n N_B2_M16_g
+ N_B2_c_142_n B2 VSS PM_OA221X2_ASAP7_75T_L%B2
x_PM_OA221X2_ASAP7_75T_L%B1 N_B1_M8_g N_B1_M17_g N_B1_M9_g N_B1_c_165_n
+ N_B1_c_166_n B1 VSS PM_OA221X2_ASAP7_75T_L%B1
x_PM_OA221X2_ASAP7_75T_L%C N_C_M10_g N_C_M18_g N_C_M11_g N_C_c_195_n N_C_c_201_n
+ C VSS PM_OA221X2_ASAP7_75T_L%C
x_PM_OA221X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_M13_d N_Y_M12_d N_Y_c_220_n Y
+ N_Y_c_223_n N_Y_c_224_n N_Y_c_225_n N_Y_c_226_n N_Y_c_228_n N_Y_c_229_n VSS
+ PM_OA221X2_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A1_M2_g 2.13359e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_A1_M2_g 0.00268443f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_A1_M2_g 2.52946e-19 $X=0.202 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_4 N_3_M1_g N_A1_M3_g 2.13359e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_5 N_3_c_5_p N_A1_c_92_n 0.00118083f $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_6 N_3_c_3_p N_A1_c_92_n 4.56852e-19 $X=0.202 $Y=0.234 $X2=0.243 $Y2=0.135
cc_7 N_3_c_7_p N_A1_c_94_n 6.07186e-19 $X=0.153 $Y=0.189 $X2=0.243 $Y2=0.135
cc_8 N_3_c_8_p N_A1_c_94_n 6.07186e-19 $X=0.153 $Y=0.135 $X2=0.243 $Y2=0.135
cc_9 N_3_c_9_p A1 3.65184e-19 $X=0.153 $Y=0.207 $X2=0.248 $Y2=0.149
cc_10 N_3_c_10_p A1 0.00347072f $X=0.252 $Y=0.234 $X2=0.248 $Y2=0.149
cc_11 N_3_c_11_p N_A2_M4_g 4.62717e-19 $X=0.342 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_12 N_3_c_12_p N_A2_M5_g 0.00173898f $X=0.528 $Y=0.174 $X2=0.243 $Y2=0.0675
cc_13 N_3_c_13_p N_A2_M5_g 2.23802e-19 $X=0.379 $Y=0.234 $X2=0.243 $Y2=0.0675
cc_14 N_3_c_14_p N_A2_c_116_n 0.00309362f $X=0.336 $Y=0.174 $X2=0.243 $Y2=0.135
cc_15 N_3_c_11_p N_A2_c_116_n 5.30479e-19 $X=0.342 $Y=0.234 $X2=0.243 $Y2=0.135
cc_16 N_3_c_12_p N_A2_c_118_n 0.00284835f $X=0.528 $Y=0.174 $X2=0.243 $Y2=0.135
cc_17 N_3_c_17_p N_A2_c_118_n 7.27996e-19 $X=0.322 $Y=0.2025 $X2=0.243 $Y2=0.135
cc_18 N_3_c_12_p A2 8.14496e-19 $X=0.528 $Y=0.174 $X2=0 $Y2=0
cc_19 N_3_c_13_p A2 0.00363104f $X=0.379 $Y=0.234 $X2=0 $Y2=0
cc_20 N_3_c_12_p N_B2_M6_g 0.00173898f $X=0.528 $Y=0.174 $X2=0.189 $Y2=0.0675
cc_21 N_3_c_21_p N_B2_M6_g 2.23802e-19 $X=0.522 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_22 N_3_c_22_p N_B2_M7_g 4.62717e-19 $X=0.593 $Y=0.234 $X2=0 $Y2=0
cc_23 N_3_c_12_p N_B2_c_140_n 0.00309362f $X=0.528 $Y=0.174 $X2=0 $Y2=0
cc_24 N_3_c_24_p N_B2_c_140_n 5.14245e-19 $X=0.531 $Y=0.234 $X2=0 $Y2=0
cc_25 N_3_c_12_p N_B2_c_142_n 0.00284835f $X=0.528 $Y=0.174 $X2=0.243 $Y2=0.135
cc_26 N_3_c_26_p N_B2_c_142_n 7.3354e-19 $X=0.542 $Y=0.2025 $X2=0.243 $Y2=0.135
cc_27 N_3_c_12_p B2 8.14496e-19 $X=0.528 $Y=0.174 $X2=0 $Y2=0
cc_28 N_3_c_21_p B2 0.00363104f $X=0.522 $Y=0.234 $X2=0 $Y2=0
cc_29 N_3_c_29_p N_B1_M8_g 2.38303e-19 $X=0.63 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_30 N_3_c_30_p N_B1_c_165_n 7.50137e-19 $X=0.668 $Y=0.234 $X2=0.243 $Y2=0.135
cc_31 N_3_c_12_p N_B1_c_166_n 3.21078e-19 $X=0.528 $Y=0.174 $X2=0.243 $Y2=0.135
cc_32 N_3_c_26_p B1 3.76498e-19 $X=0.542 $Y=0.2025 $X2=0 $Y2=0
cc_33 N_3_c_29_p B1 0.00399719f $X=0.63 $Y=0.234 $X2=0 $Y2=0
cc_34 N_3_c_34_p N_C_M10_g 2.34993e-19 $X=0.757 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_35 N_3_c_35_p N_C_M11_g 4.48264e-19 $X=0.7925 $Y=0.234 $X2=0.243 $Y2=0.0675
cc_36 N_3_c_36_p N_C_M11_g 3.95625e-19 $X=0.824 $Y=0.072 $X2=0.243 $Y2=0.0675
cc_37 N_3_M11_d N_C_c_195_n 3.78279e-19 $X=0.773 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_38 N_3_c_38_p N_C_c_195_n 9.18375e-19 $X=0.756 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_39 N_3_c_39_p N_C_c_195_n 3.82299e-19 $X=0.754 $Y=0.216 $X2=0.243 $Y2=0.135
cc_40 N_3_c_35_p N_C_c_195_n 3.33534e-19 $X=0.7925 $Y=0.234 $X2=0.243 $Y2=0.135
cc_41 N_3_c_36_p N_C_c_195_n 6.23903e-19 $X=0.824 $Y=0.072 $X2=0.243 $Y2=0.135
cc_42 N_3_c_42_p N_C_c_195_n 4.19219e-19 $X=0.837 $Y=0.189 $X2=0.243 $Y2=0.135
cc_43 N_3_c_38_p N_C_c_201_n 9.73005e-19 $X=0.756 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_44 N_3_c_44_p N_C_c_201_n 0.00149047f $X=0.757 $Y=0.072 $X2=0.243 $Y2=0.135
cc_45 N_3_c_45_p N_C_c_201_n 3.69833e-19 $X=0.837 $Y=0.117 $X2=0.243 $Y2=0.135
cc_46 N_3_c_42_p N_C_c_201_n 0.00123821f $X=0.837 $Y=0.189 $X2=0.243 $Y2=0.135
cc_47 N_3_c_39_p C 0.00167024f $X=0.754 $Y=0.216 $X2=0 $Y2=0
cc_48 N_3_c_34_p C 0.00374043f $X=0.757 $Y=0.234 $X2=0 $Y2=0
cc_49 N_3_c_49_p C 3.6188e-19 $X=0.837 $Y=0.207 $X2=0 $Y2=0
cc_50 N_3_c_5_p N_Y_M1_d 3.80485e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_51 N_3_c_5_p N_Y_M13_d 3.80277e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_52 N_3_c_5_p N_Y_c_220_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_53 N_3_c_7_p N_Y_c_220_n 0.00142308f $X=0.153 $Y=0.189 $X2=0.243 $Y2=0.0675
cc_54 N_3_c_7_p Y 3.93135e-19 $X=0.153 $Y=0.189 $X2=0 $Y2=0
cc_55 N_3_c_5_p N_Y_c_223_n 3.93676e-19 $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_56 N_3_c_56_p N_Y_c_224_n 2.04685e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_57 N_3_c_5_p N_Y_c_225_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_58 N_3_M0_g N_Y_c_226_n 3.21831e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_59 N_3_c_5_p N_Y_c_226_n 5.30465e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_60 N_3_c_60_p N_Y_c_228_n 0.00111712f $X=0.162 $Y=0.234 $X2=0 $Y2=0
cc_61 N_3_M0_g N_Y_c_229_n 3.68592e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_62 N_3_c_5_p N_Y_c_229_n 7.80348e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_63 N_3_c_63_p N_Y_c_229_n 0.00111712f $X=0.153 $Y=0.225 $X2=0 $Y2=0
cc_64 N_3_c_9_p N_Y_c_229_n 0.00111712f $X=0.153 $Y=0.207 $X2=0 $Y2=0
cc_65 VSS N_3_c_14_p 0.00126357f $X=0.336 $Y=0.174 $X2=0.243 $Y2=0.0675
cc_66 VSS N_3_c_12_p 0.00126357f $X=0.528 $Y=0.174 $X2=0 $Y2=0
cc_67 VSS N_3_c_67_p 3.73938e-19 $X=0.215 $Y=0.234 $X2=0.243 $Y2=0.149
cc_68 VSS N_3_c_11_p 3.73938e-19 $X=0.342 $Y=0.234 $X2=0 $Y2=0
cc_69 VSS N_3_c_69_p 3.73938e-19 $X=0.485 $Y=0.234 $X2=0 $Y2=0
cc_70 VSS N_3_c_12_p 0.00158021f $X=0.528 $Y=0.174 $X2=0 $Y2=0
cc_71 VSS N_3_c_24_p 3.73938e-19 $X=0.531 $Y=0.234 $X2=0 $Y2=0
cc_72 VSS N_3_c_22_p 3.73938e-19 $X=0.593 $Y=0.234 $X2=0 $Y2=0
cc_73 VSS N_3_c_44_p 3.09983e-19 $X=0.757 $Y=0.072 $X2=0 $Y2=0
cc_74 VSS N_3_c_30_p 3.73938e-19 $X=0.668 $Y=0.234 $X2=0 $Y2=0
cc_75 VSS N_3_c_36_p 2.53396e-19 $X=0.824 $Y=0.072 $X2=0.243 $Y2=0.135
cc_76 VSS N_3_c_12_p 9.24871e-19 $X=0.528 $Y=0.174 $X2=0.248 $Y2=0.149
cc_77 VSS N_3_c_38_p 0.00342838f $X=0.756 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_78 VSS N_3_c_44_p 4.44103e-19 $X=0.757 $Y=0.072 $X2=0.243 $Y2=0.135
cc_79 VSS N_3_c_38_p 0.00255008f $X=0.756 $Y=0.0675 $X2=0 $Y2=0
cc_80 VSS N_3_c_44_p 0.00718543f $X=0.757 $Y=0.072 $X2=0 $Y2=0
cc_81 VSS N_3_c_38_p 0.00381356f $X=0.756 $Y=0.0675 $X2=0 $Y2=0
cc_82 VSS N_3_c_36_p 0.00263302f $X=0.824 $Y=0.072 $X2=0 $Y2=0
cc_83 VSS N_3_c_45_p 3.06659e-19 $X=0.837 $Y=0.117 $X2=0 $Y2=0
cc_84 VSS N_3_c_14_p 0.00540341f $X=0.336 $Y=0.174 $X2=0.243 $Y2=0.0675
cc_85 VSS N_3_c_67_p 0.00127469f $X=0.215 $Y=0.234 $X2=0.243 $Y2=0.0675
cc_86 VSS N_3_c_10_p 0.0022705f $X=0.252 $Y=0.234 $X2=0.243 $Y2=0.0675
cc_87 VSS N_3_c_11_p 0.00287843f $X=0.342 $Y=0.234 $X2=0.243 $Y2=0.0675
cc_88 N_A1_M2_g N_A2_M4_g 2.48122e-19 $X=0.189 $Y=0.0675 $X2=0.336 $Y2=0.174
cc_89 N_A1_M3_g N_A2_M4_g 0.00312021f $X=0.243 $Y=0.0675 $X2=0.336 $Y2=0.174
cc_90 N_A1_M3_g N_A2_M5_g 2.53865e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.2025
cc_91 N_A1_c_92_n N_A2_c_116_n 0.00136394f $X=0.243 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_92 N_A1_c_94_n N_A2_c_118_n 9.90273e-19 $X=0.243 $Y=0.135 $X2=0.135
+ $Y2=0.2025
cc_93 N_A1_c_94_n A2 4.95137e-19 $X=0.243 $Y=0.135 $X2=0.773 $Y2=0.0675
cc_94 VSS N_A1_c_92_n 3.78404e-19 $X=0.243 $Y=0.135 $X2=0.528 $Y2=0.174
cc_95 VSS N_A1_c_92_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_96 VSS N_A1_c_94_n 8.82763e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_97 VSS N_A1_M3_g 3.37536e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_98 VSS N_A1_c_94_n 0.00371264f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_99 VSS N_A1_M3_g 0.00382057f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_100 VSS N_A1_c_92_n 0.00312836f $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_101 VSS N_A1_c_94_n 0.00265784f $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_102 VSS A1 0.00289131f $X=0.248 $Y=0.149 $X2=0.081 $Y2=0.135
cc_103 N_A2_c_118_n N_B2_c_142_n 7.63935e-19 $X=0.351 $Y=0.135 $X2=0.135
+ $Y2=0.2025
cc_104 A2 B2 4.24115e-19 $X=0.353 $Y=0.151 $X2=0.773 $Y2=0.0675
cc_105 VSS N_A2_c_116_n 3.80246e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_106 VSS N_A2_c_116_n 8.0006e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_107 VSS N_A2_c_118_n 3.18961e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_108 VSS N_A2_c_116_n 9.0655e-19 $X=0.351 $Y=0.135 $X2=0.557 $Y2=0.2025
cc_109 VSS N_A2_M4_g 4.62282e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_110 VSS N_A2_M5_g 3.4229e-19 $X=0.351 $Y=0.0675 $X2=0.739 $Y2=0.216
cc_111 VSS N_A2_c_118_n 0.00376019f $X=0.351 $Y=0.135 $X2=0.739 $Y2=0.216
cc_112 N_B2_M6_g N_B1_M8_g 2.88628e-19 $X=0.513 $Y=0.0675 $X2=0.336 $Y2=0.174
cc_113 N_B2_M7_g N_B1_M8_g 0.00353416f $X=0.567 $Y=0.0675 $X2=0.336 $Y2=0.174
cc_114 N_B2_M7_g N_B1_M9_g 2.53865e-19 $X=0.567 $Y=0.0675 $X2=0.081 $Y2=0.2025
cc_115 N_B2_c_140_n N_B1_c_165_n 0.00133245f $X=0.567 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_116 N_B2_c_142_n N_B1_c_166_n 0.00146965f $X=0.513 $Y=0.135 $X2=0.135
+ $Y2=0.2025
cc_117 B2 B1 3.25705e-19 $X=0.511 $Y=0.151 $X2=0.773 $Y2=0.0675
cc_118 VSS N_B2_c_140_n 3.80246e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_119 VSS N_B2_c_140_n 8.0006e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_120 VSS N_B2_c_142_n 3.14208e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_121 VSS N_B2_M6_g 2.52885e-19 $X=0.513 $Y=0.0675 $X2=0.754 $Y2=0.216
cc_122 VSS N_B2_c_142_n 0.00373896f $X=0.513 $Y=0.135 $X2=0.754 $Y2=0.216
cc_123 VSS N_B2_c_140_n 8.82678e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_124 VSS N_B2_M7_g 3.97719e-19 $X=0.567 $Y=0.0675 $X2=0.153 $Y2=0.207
cc_125 VSS N_B2_c_142_n 0.0313993f $X=0.513 $Y=0.135 $X2=0.756 $Y2=0.0675
cc_126 VSS N_B2_M6_g 2.38303e-19 $X=0.513 $Y=0.0675 $X2=0.557 $Y2=0.2025
cc_127 VSS N_B2_M7_g 2.64781e-19 $X=0.567 $Y=0.0675 $X2=0.557 $Y2=0.2025
cc_128 N_B1_M8_g N_C_M10_g 2.4073e-19 $X=0.621 $Y=0.0675 $X2=0.336 $Y2=0.174
cc_129 N_B1_M9_g N_C_M10_g 0.00317103f $X=0.675 $Y=0.0675 $X2=0.336 $Y2=0.174
cc_130 N_B1_M9_g N_C_M11_g 2.53865e-19 $X=0.675 $Y=0.0675 $X2=0.081 $Y2=0.2025
cc_131 N_B1_c_165_n N_C_c_195_n 0.00133355f $X=0.675 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_132 N_B1_c_166_n N_C_c_201_n 9.28358e-19 $X=0.621 $Y=0.135 $X2=0.135
+ $Y2=0.2025
cc_133 B1 C 4.64179e-19 $X=0.622 $Y=0.151 $X2=0.773 $Y2=0.0675
cc_134 VSS N_B1_c_165_n 3.80246e-19 $X=0.675 $Y=0.135 $X2=0.135 $Y2=0.135
cc_135 VSS N_B1_c_165_n 8.0006e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_136 VSS N_B1_c_166_n 3.18961e-19 $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_137 VSS N_B1_M9_g 2.41848e-19 $X=0.675 $Y=0.0675 $X2=0.153 $Y2=0.225
cc_138 VSS N_B1_c_165_n 6.22411e-19 $X=0.675 $Y=0.135 $X2=0.153 $Y2=0.225
cc_139 VSS N_B1_M8_g 2.56447e-19 $X=0.621 $Y=0.0675 $X2=0.828 $Y2=0.234
cc_140 VSS N_B1_c_166_n 0.00376032f $X=0.621 $Y=0.135 $X2=0.828 $Y2=0.234
cc_141 VSS N_B1_c_166_n 0.0313424f $X=0.621 $Y=0.135 $X2=0.322 $Y2=0.2025
cc_142 VSS N_B1_M8_g 2.38303e-19 $X=0.621 $Y=0.0675 $X2=0.557 $Y2=0.2025
cc_143 VSS N_B1_M9_g 3.89858e-19 $X=0.675 $Y=0.0675 $X2=0.542 $Y2=0.2025
cc_144 VSS B1 2.98476e-19 $X=0.622 $Y=0.151 $X2=0.528 $Y2=0.174
cc_145 VSS N_C_c_201_n 3.18961e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_146 VSS N_C_M11_g 2.64781e-19 $X=0.783 $Y=0.0675 $X2=0.542 $Y2=0.2025
cc_147 VSS N_C_M10_g 3.43731e-19 $X=0.729 $Y=0.0675 $X2=0.754 $Y2=0.216
cc_148 VSS N_C_c_201_n 8.36793e-19 $X=0.729 $Y=0.135 $X2=0.754 $Y2=0.216
cc_149 VSS N_Y_c_220_n 3.54299e-19 $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135

* END of "./OA221x2_ASAP7_75t_L.pex.sp.OA221X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA222x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:48:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA222x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA222x2_ASAP7_75t_L.pex.sp.pex"
* File: OA222x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:48:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA222X2_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c11 10 VSS 5.09652e-19 $X=0.081 $Y=0.135
c12 5 VSS 0.00171842f $X=0.081 $Y=0.135
c13 2 VSS 0.066866f $X=0.081 $Y=0.0675
r14 10 14 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.147
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA222X2_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c11 10 VSS 0.00167719f $X=0.135 $Y=0.135
c12 5 VSS 0.00113686f $X=0.135 $Y=0.135
c13 2 VSS 0.062389f $X=0.135 $Y=0.0675
r14 10 14 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.147
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OA222X2_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c11 10 VSS 0.00167719f $X=0.189 $Y=0.135
c12 5 VSS 0.00113407f $X=0.189 $Y=0.135
c13 2 VSS 0.062389f $X=0.189 $Y=0.0675
r14 10 14 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.147
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA222X2_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c11 10 VSS 7.9511e-19 $X=0.243 $Y=0.135
c12 5 VSS 0.00220625f $X=0.243 $Y=0.135
c13 2 VSS 0.0662287f $X=0.243 $Y=0.0675
r14 10 14 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.147
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OA222X2_ASAP7_75T_L%C1 2 5 7 10 16 VSS
c12 10 VSS 0.00231526f $X=0.405 $Y=0.135
c13 5 VSS 0.00216395f $X=0.405 $Y=0.135
c14 2 VSS 0.0637934f $X=0.405 $Y=0.0675
r15 10 16 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.147
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OA222X2_ASAP7_75T_L%C2 2 5 7 10 16 VSS
c14 10 VSS 0.00234157f $X=0.459 $Y=0.135
c15 5 VSS 0.00115457f $X=0.459 $Y=0.135
c16 2 VSS 0.0591635f $X=0.459 $Y=0.0675
r17 10 16 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.147
r18 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r19 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r20 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OA222X2_ASAP7_75T_L%9 2 7 10 13 15 17 18 21 22 25 27 30 32 35 39 40
+ 43 46 47 50 59 60 62 64 66 67 71 72 73 74 75 76 78 79 80 81 83 86 VSS
c58 86 VSS 4.68643e-20 $X=0.531 $Y=0.135
c59 85 VSS 6.11899e-19 $X=0.526 $Y=0.135
c60 83 VSS 5.23673e-20 $X=0.54 $Y=0.135
c61 81 VSS 9.96284e-19 $X=0.504 $Y=0.135
c62 80 VSS 2.58269e-19 $X=0.495 $Y=0.2
c63 79 VSS 0.00118967f $X=0.495 $Y=0.189
c64 78 VSS 0.00176136f $X=0.495 $Y=0.225
c65 76 VSS 0.00146362f $X=0.468 $Y=0.234
c66 75 VSS 0.00346383f $X=0.45 $Y=0.234
c67 74 VSS 0.00146362f $X=0.414 $Y=0.234
c68 73 VSS 0.00271257f $X=0.396 $Y=0.234
c69 72 VSS 9.85989e-19 $X=0.369 $Y=0.234
c70 71 VSS 0.0127088f $X=0.36 $Y=0.234
c71 67 VSS 0.00146362f $X=0.252 $Y=0.234
c72 66 VSS 0.00302652f $X=0.234 $Y=0.234
c73 65 VSS 4.63288e-19 $X=0.202 $Y=0.234
c74 64 VSS 0.00142296f $X=0.198 $Y=0.234
c75 63 VSS 0.00660983f $X=0.18 $Y=0.234
c76 62 VSS 0.00142296f $X=0.144 $Y=0.234
c77 61 VSS 4.63288e-19 $X=0.126 $Y=0.234
c78 60 VSS 0.00287317f $X=0.122 $Y=0.234
c79 59 VSS 0.00146362f $X=0.09 $Y=0.234
c80 58 VSS 0.00454946f $X=0.072 $Y=0.234
c81 51 VSS 0.00326963f $X=0.027 $Y=0.234
c82 50 VSS 0.00556194f $X=0.486 $Y=0.234
c83 48 VSS 1.45514e-19 $X=0.099 $Y=0.072
c84 47 VSS 8.46035e-21 $X=0.09 $Y=0.072
c85 46 VSS 3.8564e-19 $X=0.072 $Y=0.072
c86 45 VSS 0.00112964f $X=0.04 $Y=0.072
c87 43 VSS 3.25827e-19 $X=0.108 $Y=0.072
c88 41 VSS 0.00191981f $X=0.027 $Y=0.072
c89 40 VSS 0.00432139f $X=0.018 $Y=0.2
c90 39 VSS 0.00107066f $X=0.018 $Y=0.106
c91 38 VSS 9.39296e-19 $X=0.018 $Y=0.225
c92 35 VSS 0.00470811f $X=0.38 $Y=0.2025
c93 32 VSS 2.69461e-19 $X=0.395 $Y=0.2025
c94 30 VSS 0.00392489f $X=0.268 $Y=0.2025
c95 25 VSS 0.00358217f $X=0.056 $Y=0.2025
c96 22 VSS 2.69461e-19 $X=0.071 $Y=0.2025
c97 21 VSS 0.0023085f $X=0.108 $Y=0.0675
c98 17 VSS 5.76042e-19 $X=0.125 $Y=0.0675
c99 13 VSS 0.00418741f $X=0.567 $Y=0.135
c100 10 VSS 0.0645347f $X=0.567 $Y=0.0675
c101 2 VSS 0.0618812f $X=0.513 $Y=0.0675
r102 85 86 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.526
+ $Y=0.135 $X2=0.531 $Y2=0.135
r103 83 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.135 $X2=0.531 $Y2=0.135
r104 83 84 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.54 $Y=0.135 $X2=0.54
+ $Y2=0.135
r105 81 85 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.135 $X2=0.526 $Y2=0.135
r106 79 80 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.189 $X2=0.495 $Y2=0.2
r107 78 80 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.225 $X2=0.495 $Y2=0.2
r108 77 81 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.495 $Y=0.144 $X2=0.504 $Y2=0.135
r109 77 79 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.144 $X2=0.495 $Y2=0.189
r110 75 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r111 74 75 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.45 $Y2=0.234
r112 73 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r113 71 72 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.369 $Y2=0.234
r114 69 73 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r115 69 72 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.369 $Y2=0.234
r116 66 67 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r117 65 66 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.234 $X2=0.234 $Y2=0.234
r118 64 65 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.202 $Y2=0.234
r119 63 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r120 62 63 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.18 $Y2=0.234
r121 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r122 60 61 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.122
+ $Y=0.234 $X2=0.126 $Y2=0.234
r123 59 60 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.122 $Y2=0.234
r124 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r125 56 71 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.36 $Y2=0.234
r126 56 67 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.252 $Y2=0.234
r127 53 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.072 $Y2=0.234
r128 51 53 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.054 $Y2=0.234
r129 50 78 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.486 $Y=0.234 $X2=0.495 $Y2=0.225
r130 50 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.468 $Y2=0.234
r131 47 48 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.099 $Y2=0.072
r132 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.072 $X2=0.09 $Y2=0.072
r133 45 46 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.072 $X2=0.072 $Y2=0.072
r134 43 48 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.099 $Y2=0.072
r135 41 45 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.072 $X2=0.04 $Y2=0.072
r136 39 40 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.106 $X2=0.018 $Y2=0.2
r137 38 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r138 38 40 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2
r139 37 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.081 $X2=0.027 $Y2=0.072
r140 37 39 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.106
r141 35 69 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r142 32 35 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.38 $Y2=0.2025
r143 30 56 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r144 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.268 $Y2=0.2025
r145 25 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r146 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r147 21 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072
+ $X2=0.108 $Y2=0.072
r148 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r149 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r150 13 84 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.567
+ $Y=0.135 $X2=0.54 $Y2=0.135
r151 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.135 $X2=0.567 $Y2=0.2025
r152 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.0675 $X2=0.567 $Y2=0.135
r153 5 84 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.54 $Y2=0.135
r154 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r155 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OA222X2_ASAP7_75T_L%Y 1 2 6 7 10 14 16 17 21 27 28 33 35 36 37 VSS
c19 39 VSS 7.27544e-19 $X=0.621 $Y=0.207
c20 37 VSS 6.80214e-20 $X=0.621 $Y=0.1455
c21 36 VSS 7.60733e-19 $X=0.621 $Y=0.144
c22 35 VSS 0.00342139f $X=0.621 $Y=0.126
c23 34 VSS 0.00131846f $X=0.621 $Y=0.07
c24 33 VSS 0.00245372f $X=0.624 $Y=0.147
c25 31 VSS 6.50936e-19 $X=0.621 $Y=0.225
c26 29 VSS 0.00215218f $X=0.599 $Y=0.234
c27 28 VSS 0.00361204f $X=0.586 $Y=0.234
c28 27 VSS 0.0020117f $X=0.549 $Y=0.234
c29 26 VSS 0.00537021f $X=0.612 $Y=0.234
c30 21 VSS 0.00131996f $X=0.54 $Y=0.216
c31 17 VSS 0.00354758f $X=0.586 $Y=0.036
c32 16 VSS 0.00311271f $X=0.554 $Y=0.036
c33 14 VSS 0.00901311f $X=0.54 $Y=0.036
c34 11 VSS 0.0075137f $X=0.612 $Y=0.036
c35 10 VSS 0.010507f $X=0.54 $Y=0.2025
c36 6 VSS 5.945e-19 $X=0.557 $Y=0.2025
c37 1 VSS 5.58795e-19 $X=0.557 $Y=0.0675
r38 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.189 $X2=0.621 $Y2=0.207
r39 36 37 0.101852 $w=1.8e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.144 $X2=0.621 $Y2=0.1455
r40 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.126 $X2=0.621 $Y2=0.144
r41 34 35 3.80247 $w=1.8e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.07 $X2=0.621 $Y2=0.126
r42 33 38 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.147 $X2=0.621 $Y2=0.189
r43 33 37 0.101852 $w=1.8e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.147 $X2=0.621 $Y2=0.1455
r44 31 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.207
r45 30 34 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.07
r46 28 29 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.586
+ $Y=0.234 $X2=0.599 $Y2=0.234
r47 27 28 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.549
+ $Y=0.234 $X2=0.586 $Y2=0.234
r48 26 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r49 26 29 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.599 $Y2=0.234
r50 19 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.54 $Y=0.225 $X2=0.549 $Y2=0.234
r51 19 21 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.225 $X2=0.54 $Y2=0.216
r52 16 17 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.554
+ $Y=0.036 $X2=0.586 $Y2=0.036
r53 13 16 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.554 $Y2=0.036
r54 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r55 11 30 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r56 11 17 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.586 $Y2=0.036
r57 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.216 $X2=0.54
+ $Y2=0.216
r58 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r59 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r60 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r61 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.523
+ $Y=0.0675 $X2=0.54 $Y2=0.0675
r62 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.557
+ $Y=0.0675 $X2=0.54 $Y2=0.0675
.ends


* END of "./OA222x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA222x2_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 C1 C2 Y
* 
* Y	Y
* C2	C2
* C1	C1
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 N_9_M0_d N_A1_M0_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_10 N_A2_M1_g N_9_M1_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_11 N_B2_M2_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_10 N_B1_M3_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_11 N_C1_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 VSS N_C2_M5_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 N_Y_M6_d N_9_M6_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M7 N_Y_M7_d N_9_M7_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M8 noxref_13 N_A1_M8_g N_9_M8_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M9 VDD N_A2_M9_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M10 noxref_14 N_B2_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M11 N_9_M11_d N_B1_M11_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M12 noxref_15 N_C1_M12_g N_9_M12_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M13 VDD N_C2_M13_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M14 N_Y_M14_d N_9_M14_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M15 N_Y_M15_d N_9_M15_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
*
* 
* .include "OA222x2_ASAP7_75t_L.pex.sp.OA222X2_ASAP7_75T_L.pxi"
* BEGIN of "./OA222x2_ASAP7_75t_L.pex.sp.OA222X2_ASAP7_75T_L.pxi"
* File: OA222x2_ASAP7_75t_L.pex.sp.OA222X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:48:26 2017
* 
x_PM_OA222X2_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M8_g N_A1_c_3_p A1 VSS
+ PM_OA222X2_ASAP7_75T_L%A1
x_PM_OA222X2_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_13_n N_A2_M9_g N_A2_c_14_n A2 VSS
+ PM_OA222X2_ASAP7_75T_L%A2
x_PM_OA222X2_ASAP7_75T_L%B2 N_B2_M2_g N_B2_c_25_n N_B2_M10_g N_B2_c_26_n B2 VSS
+ PM_OA222X2_ASAP7_75T_L%B2
x_PM_OA222X2_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_36_n N_B1_M11_g N_B1_c_37_n B1 VSS
+ PM_OA222X2_ASAP7_75T_L%B1
x_PM_OA222X2_ASAP7_75T_L%C1 N_C1_M4_g N_C1_c_47_p N_C1_M12_g N_C1_c_45_n C1 VSS
+ PM_OA222X2_ASAP7_75T_L%C1
x_PM_OA222X2_ASAP7_75T_L%C2 N_C2_M5_g N_C2_c_58_n N_C2_M13_g N_C2_c_59_n C2 VSS
+ PM_OA222X2_ASAP7_75T_L%C2
x_PM_OA222X2_ASAP7_75T_L%9 N_9_M6_g N_9_M14_g N_9_M7_g N_9_c_90_n N_9_M15_g
+ N_9_M1_s N_9_M0_d N_9_c_96_p N_9_M8_s N_9_c_71_n N_9_M11_d N_9_c_81_n
+ N_9_M12_s N_9_c_85_n N_9_c_98_p N_9_c_72_n N_9_c_101_p N_9_c_95_p N_9_c_73_n
+ N_9_c_121_p N_9_c_75_n N_9_c_126_p N_9_c_77_n N_9_c_79_n N_9_c_106_p
+ N_9_c_82_n N_9_c_107_p N_9_c_109_p N_9_c_108_p N_9_c_86_n N_9_c_128_p
+ N_9_c_91_n N_9_c_118_p N_9_c_93_n N_9_c_119_p N_9_c_94_n N_9_c_120_p
+ N_9_c_114_p VSS PM_OA222X2_ASAP7_75T_L%9
x_PM_OA222X2_ASAP7_75T_L%Y N_Y_M7_d N_Y_M6_d N_Y_M15_d N_Y_M14_d N_Y_c_132_n
+ N_Y_c_146_n N_Y_c_133_n N_Y_c_135_n N_Y_c_136_n N_Y_c_141_n N_Y_c_142_n Y
+ N_Y_c_129_n N_Y_c_144_n N_Y_c_145_n VSS PM_OA222X2_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00372052f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_13_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p N_A2_c_14_n 0.00477924f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A1_M0_g N_B2_M2_g 2.74891e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 N_A1_c_3_p N_9_c_71_n 0.00141058f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_6 N_A1_c_3_p N_9_c_72_n 0.00311007f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_7 N_A1_M0_g N_9_c_73_n 2.68514e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_8 N_A1_c_3_p N_9_c_73_n 0.00121543f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_A1_M0_g N_9_c_75_n 2.64276e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_10 N_A1_c_3_p N_9_c_75_n 0.00124805f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 VSS N_A1_M0_g 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_12 N_A2_M1_g N_B2_M2_g 0.00335739f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_13 N_A2_c_13_n N_B2_c_25_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 N_A2_c_14_n N_B2_c_26_n 0.00406615f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 N_A2_M1_g N_B1_M3_g 2.74891e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_A2_M1_g N_9_c_77_n 2.56935e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_17 N_A2_c_14_n N_9_c_77_n 0.00123064f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_18 VSS N_A2_M1_g 3.47199e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 VSS N_A2_c_14_n 5.30079e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_20 N_B2_M2_g N_B1_M3_g 0.00372052f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_21 N_B2_c_25_n N_B1_c_36_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 N_B2_c_26_n N_B1_c_37_n 0.00477924f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 N_B2_M2_g N_9_c_79_n 2.56935e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 N_B2_c_26_n N_9_c_79_n 0.00123064f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_25 VSS N_B2_M2_g 3.57119e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 VSS N_B2_c_26_n 5.37372e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_27 N_B1_c_37_n N_C1_c_45_n 5.27113e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_28 N_B1_c_37_n N_9_c_81_n 0.00153032f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_29 N_B1_M3_g N_9_c_82_n 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_B1_c_37_n N_9_c_82_n 0.00124805f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 VSS N_B1_M3_g 2.08515e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_32 VSS N_B1_M3_g 2.76185e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_33 VSS N_B1_c_37_n 0.0012322f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_34 N_C1_M4_g N_C2_M5_g 0.00347357f $X=0.405 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_35 N_C1_c_47_p N_C2_c_58_n 9.33263e-19 $X=0.405 $Y=0.135 $X2=0.243 $Y2=0.135
cc_36 N_C1_c_45_n N_C2_c_59_n 0.00575765f $X=0.405 $Y=0.135 $X2=0.243 $Y2=0.135
cc_37 N_C1_M4_g N_9_M6_g 2.34385e-19 $X=0.405 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_38 N_C1_c_45_n N_9_c_85_n 0.00153032f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_39 N_C1_M4_g N_9_c_86_n 2.64276e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_40 N_C1_c_45_n N_9_c_86_n 0.00125352f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_41 VSS N_C1_c_45_n 4.64783e-19 $X=0.405 $Y=0.135 $X2=0.243 $Y2=0.135
cc_42 VSS N_C1_c_45_n 0.0011319f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_43 VSS N_C1_M4_g 2.64276e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_44 VSS N_C1_c_45_n 0.00125352f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_45 N_C2_M5_g N_9_M6_g 0.00287079f $X=0.459 $Y=0.0675 $X2=0.405 $Y2=0.0675
cc_46 N_C2_M5_g N_9_M7_g 2.34385e-19 $X=0.459 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_47 N_C2_c_58_n N_9_c_90_n 0.00109069f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_48 N_C2_M5_g N_9_c_91_n 2.64276e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_49 N_C2_c_59_n N_9_c_91_n 0.00125352f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_50 N_C2_c_59_n N_9_c_93_n 0.00306679f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_51 N_C2_c_59_n N_9_c_94_n 0.00306679f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_52 VSS N_C2_M5_g 2.87532e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_53 VSS N_C2_c_59_n 0.00125352f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_54 VSS N_C2_c_59_n 0.00114532f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_55 N_C2_c_59_n N_Y_c_129_n 3.09931e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_56 VSS N_9_c_95_p 2.63376e-19 $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_57 VSS N_9_c_96_p 0.00359992f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_58 VSS N_9_c_71_n 0.00138157f $X=0.056 $Y=0.2025 $X2=0 $Y2=0
cc_59 VSS N_9_c_98_p 3.56073e-19 $X=0.018 $Y=0.106 $X2=0 $Y2=0
cc_60 VSS N_9_c_95_p 0.00256253f $X=0.072 $Y=0.072 $X2=0 $Y2=0
cc_61 VSS N_9_c_96_p 0.00333673f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_62 VSS N_9_c_101_p 4.46493e-19 $X=0.108 $Y=0.072 $X2=0 $Y2=0
cc_63 VSS N_9_c_96_p 0.00250965f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_64 VSS N_9_c_95_p 0.00707171f $X=0.072 $Y=0.072 $X2=0 $Y2=0
cc_65 VSS N_9_c_81_n 0.00138157f $X=0.268 $Y=0.2025 $X2=0 $Y2=0
cc_66 VSS N_9_c_101_p 2.90501e-19 $X=0.108 $Y=0.072 $X2=0 $Y2=0
cc_67 VSS N_9_c_106_p 8.02788e-19 $X=0.234 $Y=0.234 $X2=0 $Y2=0
cc_68 VSS N_9_c_107_p 8.02788e-19 $X=0.36 $Y=0.234 $X2=0 $Y2=0
cc_69 VSS N_9_c_108_p 2.14558e-19 $X=0.396 $Y=0.234 $X2=0 $Y2=0
cc_70 VSS N_9_c_109_p 2.14558e-19 $X=0.369 $Y=0.234 $X2=0 $Y2=0
cc_71 N_9_c_90_n N_Y_M7_d 3.80351e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_72 N_9_c_90_n N_Y_M15_d 3.80315e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_73 N_9_c_93_n N_Y_c_132_n 0.00141371f $X=0.495 $Y=0.189 $X2=0.081 $Y2=0.135
cc_74 N_9_c_90_n N_Y_c_133_n 3.2373e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_75 N_9_c_114_p N_Y_c_133_n 3.16052e-19 $X=0.531 $Y=0.135 $X2=0 $Y2=0
cc_76 N_9_M7_g N_Y_c_135_n 4.59758e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_77 N_9_M7_g N_Y_c_136_n 3.68592e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_78 N_9_c_90_n N_Y_c_136_n 4.61714e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_79 N_9_c_118_p N_Y_c_136_n 0.00111326f $X=0.495 $Y=0.225 $X2=0 $Y2=0
cc_80 N_9_c_119_p N_Y_c_136_n 0.00111326f $X=0.495 $Y=0.2 $X2=0 $Y2=0
cc_81 N_9_c_120_p N_Y_c_136_n 6.29344e-19 $X=0.54 $Y=0.135 $X2=0 $Y2=0
cc_82 N_9_c_121_p N_Y_c_141_n 0.00111326f $X=0.486 $Y=0.234 $X2=0 $Y2=0
cc_83 N_9_M7_g N_Y_c_142_n 2.35972e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_84 N_9_c_90_n N_Y_c_129_n 4.54439e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_85 N_9_c_120_p N_Y_c_144_n 4.01628e-19 $X=0.54 $Y=0.135 $X2=0 $Y2=0
cc_86 N_9_c_93_n N_Y_c_145_n 4.32146e-19 $X=0.495 $Y=0.189 $X2=0 $Y2=0
cc_87 VSS N_9_c_126_p 3.16424e-19 $X=0.122 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_88 VSS N_9_c_106_p 3.16424e-19 $X=0.234 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_89 VSS N_9_c_128_p 3.56327e-19 $X=0.45 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_90 VSS N_Y_c_146_n 2.23372e-19 $X=0.432 $Y=0.036 $X2=0.189 $Y2=0.147
cc_91 VSS N_Y_c_133_n 3.94427e-19 $X=0.432 $Y=0.036 $X2=0 $Y2=0

* END of "./OA222x2_ASAP7_75t_L.pex.sp.OA222X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA22x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:48:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA22x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA22x2_ASAP7_75t_L.pex.sp.pex"
* File: OA22x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:48:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA22X2_ASAP7_75T_L%3 2 7 10 15 17 18 21 22 23 26 27 30 33 35 38 39 40
+ 42 46 47 48 49 51 53 56 57 58 VSS
c44 61 VSS 2.87023e-19 $X=0.189 $Y=0.135
c45 58 VSS 0.0018889f $X=0.342 $Y=0.234
c46 57 VSS 0.00314389f $X=0.321 $Y=0.234
c47 56 VSS 0.0076088f $X=0.289 $Y=0.234
c48 55 VSS 0.00473092f $X=0.239 $Y=0.234
c49 53 VSS 0.00471375f $X=0.378 $Y=0.234
c50 51 VSS 0.00344625f $X=0.198 $Y=0.234
c51 48 VSS 2.17889e-19 $X=0.321 $Y=0.072
c52 47 VSS 5.42127e-20 $X=0.289 $Y=0.072
c53 46 VSS 5.67855e-19 $X=0.256 $Y=0.072
c54 45 VSS 5.01107e-19 $X=0.244 $Y=0.072
c55 44 VSS 0.00292248f $X=0.239 $Y=0.072
c56 40 VSS 0.0022257f $X=0.198 $Y=0.072
c57 39 VSS 9.51753e-19 $X=0.189 $Y=0.203
c58 38 VSS 0.00196644f $X=0.189 $Y=0.185
c59 37 VSS 0.0012698f $X=0.189 $Y=0.225
c60 35 VSS 5.39386e-19 $X=0.189 $Y=0.121
c61 34 VSS 0.00123725f $X=0.189 $Y=0.103
c62 33 VSS 1.73808e-19 $X=0.189 $Y=0.126
c63 30 VSS 0.0130223f $X=0.151 $Y=0.135
c64 27 VSS 0.00194598f $X=0.18 $Y=0.135
c65 26 VSS 0.00498479f $X=0.378 $Y=0.2025
c66 22 VSS 6.13748e-19 $X=0.395 $Y=0.2025
c67 21 VSS 0.0024706f $X=0.324 $Y=0.0675
c68 17 VSS 7.42562e-19 $X=0.341 $Y=0.0675
c69 10 VSS 0.0655916f $X=0.135 $Y=0.0675
c70 2 VSS 0.0651466f $X=0.081 $Y=0.0675
r71 57 58 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.321
+ $Y=0.234 $X2=0.342 $Y2=0.234
r72 56 57 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.289
+ $Y=0.234 $X2=0.321 $Y2=0.234
r73 55 56 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.239
+ $Y=0.234 $X2=0.289 $Y2=0.234
r74 53 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.342 $Y2=0.234
r75 51 55 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.239 $Y2=0.234
r76 48 49 0.101852 $w=1.8e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.321
+ $Y=0.072 $X2=0.3225 $Y2=0.072
r77 47 48 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.289
+ $Y=0.072 $X2=0.321 $Y2=0.072
r78 46 47 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.072 $X2=0.289 $Y2=0.072
r79 45 46 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.244
+ $Y=0.072 $X2=0.256 $Y2=0.072
r80 44 45 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.239
+ $Y=0.072 $X2=0.244 $Y2=0.072
r81 42 49 0.101852 $w=1.8e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.072 $X2=0.3225 $Y2=0.072
r82 40 44 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.072 $X2=0.239 $Y2=0.072
r83 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.185 $X2=0.189 $Y2=0.203
r84 37 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.225 $X2=0.198 $Y2=0.234
r85 37 39 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.203
r86 36 61 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.135
r87 36 38 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.185
r88 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.103 $X2=0.189 $Y2=0.121
r89 33 61 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.135
r90 33 35 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.121
r91 32 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.081 $X2=0.198 $Y2=0.072
r92 32 34 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.081 $X2=0.189 $Y2=0.103
r93 29 30 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.151 $Y=0.135 $X2=0.151
+ $Y2=0.135
r94 27 61 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.189 $Y2=0.135
r95 27 29 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.151 $Y2=0.135
r96 26 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r97 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r98 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r99 21 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.072 $X2=0.324
+ $Y2=0.072
r100 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r101 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r102 13 30 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.151 $Y2=0.135
r103 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r104 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r105 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r106 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r107 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA22X2_ASAP7_75T_L%A1 2 5 7 14 VSS
c16 14 VSS 0.0050469f $X=0.281 $Y=0.14
c17 5 VSS 0.00473147f $X=0.297 $Y=0.135
c18 2 VSS 0.0650113f $X=0.297 $Y=0.0675
r19 13 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.28 $Y=0.135 $X2=0.28
+ $Y2=0.135
r20 5 13 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.28 $Y2=0.135
r21 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OA22X2_ASAP7_75T_L%A2 2 5 7 14 VSS
c16 14 VSS 0.00178683f $X=0.35 $Y=0.137
c17 5 VSS 0.00106707f $X=0.351 $Y=0.135
c18 2 VSS 0.0620629f $X=0.351 $Y=0.0675
r19 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r20 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r21 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OA22X2_ASAP7_75T_L%B2 2 5 7 15 VSS
c11 15 VSS 0.00352205f $X=0.405 $Y=0.138
c12 5 VSS 0.00119707f $X=0.405 $Y=0.135
c13 2 VSS 0.0615465f $X=0.405 $Y=0.0675
r14 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OA22X2_ASAP7_75T_L%B1 2 5 7 14 VSS
c9 14 VSS 0.0119976f $X=0.458 $Y=0.138
c10 5 VSS 0.00227588f $X=0.459 $Y=0.135
c11 2 VSS 0.064914f $X=0.459 $Y=0.0675
r12 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OA22X2_ASAP7_75T_L%Y 1 2 6 7 10 12 14 16 18 22 23 25 30 33 VSS
c18 33 VSS 6.97033e-19 $X=0.0995 $Y=0.234
c19 32 VSS 0.00317685f $X=0.091 $Y=0.234
c20 30 VSS 0.00287243f $X=0.108 $Y=0.234
c21 25 VSS 6.97033e-19 $X=0.0995 $Y=0.036
c22 24 VSS 0.00317685f $X=0.091 $Y=0.036
c23 23 VSS 0.0104531f $X=0.108 $Y=0.036
c24 22 VSS 0.00306745f $X=0.108 $Y=0.036
c25 18 VSS 9.31565e-19 $X=0.081 $Y=0.1845
c26 16 VSS 0.00161393f $X=0.081 $Y=0.126
c27 15 VSS 6.07644e-19 $X=0.081 $Y=0.063
c28 14 VSS 2.54708e-19 $X=0.081 $Y=0.141
c29 12 VSS 0.0012131f $X=0.081 $Y=0.225
c30 10 VSS 0.0104516f $X=0.108 $Y=0.2025
c31 6 VSS 5.58795e-19 $X=0.125 $Y=0.2025
c32 1 VSS 5.58795e-19 $X=0.125 $Y=0.0675
r33 32 33 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.091
+ $Y=0.234 $X2=0.0995 $Y2=0.234
r34 30 33 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.0995 $Y2=0.234
r35 27 32 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.234 $X2=0.091 $Y2=0.234
r36 24 25 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.091
+ $Y=0.036 $X2=0.0995 $Y2=0.036
r37 22 25 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.0995 $Y2=0.036
r38 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r39 19 24 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.036 $X2=0.091 $Y2=0.036
r40 17 18 2.4125 $w=2e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.144 $X2=0.081 $Y2=0.1845
r41 15 16 3.75278 $w=2e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.063 $X2=0.081 $Y2=0.126
r42 14 17 0.178704 $w=2e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.141 $X2=0.081 $Y2=0.144
r43 14 16 0.893519 $w=2e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.141 $X2=0.081 $Y2=0.126
r44 12 27 0.00634181 $w=2e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.225 $X2=0.081 $Y2=0.234
r45 12 18 2.4125 $w=2e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.225 $X2=0.081 $Y2=0.1845
r46 11 19 0.00634181 $w=2e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.045 $X2=0.081 $Y2=0.036
r47 11 15 1.07222 $w=2e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.045 $X2=0.081 $Y2=0.063
r48 10 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r49 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r50 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r51 5 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r52 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r53 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OA22x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA22x2_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 Y
* 
* Y	Y
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_3_M2_d N_A1_M2_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 noxref_9 N_A2_M3_g N_3_M3_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 VSS N_B2_M4_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 noxref_9 N_B1_M5_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 N_Y_M6_d N_3_M6_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M7 N_Y_M7_d N_3_M7_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M8 noxref_10 N_A1_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M9 N_3_M9_d N_A2_M9_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M10 noxref_11 N_B2_M10_g N_3_M10_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M11 VDD N_B1_M11_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "OA22x2_ASAP7_75t_L.pex.sp.OA22X2_ASAP7_75T_L.pxi"
* BEGIN of "./OA22x2_ASAP7_75t_L.pex.sp.OA22X2_ASAP7_75T_L.pxi"
* File: OA22x2_ASAP7_75t_L.pex.sp.OA22X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:48:48 2017
* 
x_PM_OA22X2_ASAP7_75T_L%3 N_3_M0_g N_3_M6_g N_3_M1_g N_3_M7_g N_3_M3_s N_3_M2_d
+ N_3_c_11_p N_3_M10_s N_3_M9_d N_3_c_12_p N_3_c_24_p N_3_c_3_p N_3_c_5_p
+ N_3_c_6_p N_3_c_31_p N_3_c_7_p N_3_c_28_p N_3_c_16_p N_3_c_8_p N_3_c_36_p
+ N_3_c_1_p N_3_c_13_p N_3_c_34_p N_3_c_10_p N_3_c_9_p N_3_c_2_p N_3_c_15_p VSS
+ PM_OA22X2_ASAP7_75T_L%3
x_PM_OA22X2_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_47_n N_A1_M8_g A1 VSS
+ PM_OA22X2_ASAP7_75T_L%A1
x_PM_OA22X2_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_68_n N_A2_M9_g A2 VSS
+ PM_OA22X2_ASAP7_75T_L%A2
x_PM_OA22X2_ASAP7_75T_L%B2 N_B2_M4_g N_B2_c_80_n N_B2_M10_g B2 VSS
+ PM_OA22X2_ASAP7_75T_L%B2
x_PM_OA22X2_ASAP7_75T_L%B1 N_B1_M5_g N_B1_c_93_n N_B1_M11_g B1 VSS
+ PM_OA22X2_ASAP7_75T_L%B1
x_PM_OA22X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_M7_d N_Y_M6_d N_Y_c_99_n
+ N_Y_c_100_n Y N_Y_c_104_n N_Y_c_107_n N_Y_c_114_p N_Y_c_110_n N_Y_c_111_n
+ N_Y_c_112_n N_Y_c_113_n VSS PM_OA22X2_ASAP7_75T_L%Y
cc_1 N_3_c_1_p N_A1_M2_g 3.51117e-19 $X=0.321 $Y=0.072 $X2=0.297 $Y2=0.0675
cc_2 N_3_c_2_p N_A1_M2_g 4.08036e-19 $X=0.321 $Y=0.234 $X2=0.297 $Y2=0.0675
cc_3 N_3_c_3_p N_A1_c_47_n 2.94734e-19 $X=0.151 $Y=0.135 $X2=0.297 $Y2=0.135
cc_4 N_3_c_1_p N_A1_c_47_n 2.72188e-19 $X=0.321 $Y=0.072 $X2=0.297 $Y2=0.135
cc_5 N_3_c_5_p A1 0.00126571f $X=0.189 $Y=0.126 $X2=0.281 $Y2=0.14
cc_6 N_3_c_6_p A1 7.07604e-19 $X=0.189 $Y=0.121 $X2=0.281 $Y2=0.14
cc_7 N_3_c_7_p A1 7.65941e-19 $X=0.189 $Y=0.203 $X2=0.281 $Y2=0.14
cc_8 N_3_c_8_p A1 0.00355645f $X=0.256 $Y=0.072 $X2=0.281 $Y2=0.14
cc_9 N_3_c_9_p A1 0.00394919f $X=0.289 $Y=0.234 $X2=0.281 $Y2=0.14
cc_10 N_3_c_10_p N_A2_M3_g 2.49978e-19 $X=0.378 $Y=0.234 $X2=0.297 $Y2=0.0675
cc_11 N_3_c_11_p A2 0.0348811f $X=0.324 $Y=0.0675 $X2=0.281 $Y2=0.14
cc_12 N_3_c_12_p A2 0.00247061f $X=0.378 $Y=0.2025 $X2=0.281 $Y2=0.14
cc_13 N_3_c_13_p A2 9.80889e-19 $X=0.3225 $Y=0.072 $X2=0.281 $Y2=0.14
cc_14 N_3_c_10_p A2 0.00336649f $X=0.378 $Y=0.234 $X2=0.281 $Y2=0.14
cc_15 N_3_c_15_p A2 3.783e-19 $X=0.342 $Y=0.234 $X2=0.281 $Y2=0.14
cc_16 N_3_c_16_p B2 7.04392e-19 $X=0.324 $Y=0.072 $X2=0 $Y2=0
cc_17 N_3_c_12_p B1 7.81587e-19 $X=0.378 $Y=0.2025 $X2=0.281 $Y2=0.14
cc_18 N_3_c_10_p B1 7.11117e-19 $X=0.378 $Y=0.234 $X2=0.281 $Y2=0.14
cc_19 N_3_c_3_p N_Y_M1_d 3.80663e-19 $X=0.151 $Y=0.135 $X2=0.297 $Y2=0.0675
cc_20 N_3_c_3_p N_Y_M7_d 3.80663e-19 $X=0.151 $Y=0.135 $X2=0.297 $Y2=0.2025
cc_21 N_3_c_3_p N_Y_c_99_n 8.00061e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_22 N_3_M0_g N_Y_c_100_n 4.84388e-19 $X=0.081 $Y=0.0675 $X2=0.28 $Y2=0.135
cc_23 N_3_c_7_p N_Y_c_100_n 3.95568e-19 $X=0.189 $Y=0.203 $X2=0.28 $Y2=0.135
cc_24 N_3_c_24_p Y 5.48227e-19 $X=0.18 $Y=0.135 $X2=0.281 $Y2=0.14
cc_25 N_3_c_3_p Y 0.00174918f $X=0.151 $Y=0.135 $X2=0.281 $Y2=0.14
cc_26 N_3_M0_g N_Y_c_104_n 0.00127573f $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_3_c_3_p N_Y_c_104_n 5.42937e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_28 N_3_c_28_p N_Y_c_104_n 6.68816e-19 $X=0.198 $Y=0.072 $X2=0 $Y2=0
cc_29 N_3_M0_g N_Y_c_107_n 9.43594e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_3_c_3_p N_Y_c_107_n 5.42937e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_31 N_3_c_31_p N_Y_c_107_n 3.95568e-19 $X=0.189 $Y=0.185 $X2=0 $Y2=0
cc_32 N_3_c_3_p N_Y_c_110_n 8.00061e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_33 N_3_c_3_p N_Y_c_111_n 3.2443e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_34 N_3_c_34_p N_Y_c_112_n 3.79805e-19 $X=0.198 $Y=0.234 $X2=0 $Y2=0
cc_35 N_3_c_3_p N_Y_c_113_n 3.2443e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_36 VSS N_3_c_36_p 3.3868e-19 $X=0.289 $Y=0.072 $X2=0.297 $Y2=0.0675
cc_37 VSS N_3_c_11_p 0.00373659f $X=0.324 $Y=0.0675 $X2=0 $Y2=0
cc_38 VSS N_3_c_36_p 0.00274491f $X=0.289 $Y=0.072 $X2=0 $Y2=0
cc_39 VSS N_3_c_11_p 0.0036864f $X=0.324 $Y=0.0675 $X2=0 $Y2=0
cc_40 VSS N_3_c_12_p 0.00158654f $X=0.378 $Y=0.2025 $X2=0 $Y2=0
cc_41 VSS N_3_c_11_p 0.0019294f $X=0.324 $Y=0.0675 $X2=0 $Y2=0
cc_42 VSS N_3_c_36_p 0.0066952f $X=0.289 $Y=0.072 $X2=0 $Y2=0
cc_43 VSS N_3_c_11_p 6.04418e-19 $X=0.324 $Y=0.0675 $X2=0 $Y2=0
cc_44 VSS N_3_c_15_p 2.5707e-19 $X=0.342 $Y=0.234 $X2=0.297 $Y2=0.0675
cc_45 N_A1_M2_g N_A2_M3_g 0.0036697f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_46 N_A1_c_47_n N_A2_c_68_n 0.00104216f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_47 A1 A2 0.00369736f $X=0.281 $Y=0.14 $X2=0.135 $Y2=0.2025
cc_48 N_A1_M2_g N_B2_M4_g 3.03912e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_49 VSS N_A1_c_47_n 4.0003e-19 $X=0.297 $Y=0.135 $X2=0.307 $Y2=0.0675
cc_50 VSS A1 0.00129736f $X=0.281 $Y=0.14 $X2=0.307 $Y2=0.0675
cc_51 VSS N_A1_M2_g 2.64781e-19 $X=0.297 $Y=0.0675 $X2=0.361 $Y2=0.2025
cc_52 N_A2_M3_g N_B2_M4_g 0.00361888f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_53 N_A2_c_68_n N_B2_c_80_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_54 A2 B2 0.00260149f $X=0.35 $Y=0.137 $X2=0.135 $Y2=0.2025
cc_55 N_A2_M3_g N_B1_M5_g 2.69148e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_56 A2 B1 3.68434e-19 $X=0.35 $Y=0.137 $X2=0.135 $Y2=0.2025
cc_57 VSS N_A2_M3_g 3.51619e-19 $X=0.351 $Y=0.0675 $X2=0.378 $Y2=0.2025
cc_58 VSS A2 9.28179e-19 $X=0.35 $Y=0.137 $X2=0.378 $Y2=0.2025
cc_59 N_B2_M4_g N_B1_M5_g 0.00323392f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_60 N_B2_c_80_n N_B1_c_93_n 9.33263e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_61 B2 B1 0.00297914f $X=0.405 $Y=0.138 $X2=0.135 $Y2=0.2025
cc_62 VSS B2 0.00238347f $X=0.405 $Y=0.138 $X2=0.395 $Y2=0.2025
cc_63 VSS B2 0.00451214f $X=0.405 $Y=0.138 $X2=0.378 $Y2=0.2025
cc_64 VSS N_B2_M4_g 2.34993e-19 $X=0.405 $Y=0.0675 $X2=0.151 $Y2=0.135
cc_65 VSS N_B1_M5_g 3.41852e-19 $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.081
cc_66 VSS B1 5.62514e-19 $X=0.458 $Y=0.138 $X2=0.189 $Y2=0.081
cc_67 VSS N_Y_c_114_p 2.40824e-19 $X=0.108 $Y=0.036 $X2=0.361 $Y2=0.2025

* END of "./OA22x2_ASAP7_75t_L.pex.sp.OA22X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA31x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:49:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA31x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA31x2_ASAP7_75t_L.pex.sp.pex"
* File: OA31x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:49:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA31X2_ASAP7_75T_L%A1 2 7 10 13 18 21 VSS
c24 21 VSS 0.00102095f $X=0.083 $Y=0.152
c25 18 VSS 0.00241334f $X=0.081 $Y=0.135
c26 10 VSS 0.0721423f $X=0.135 $Y=0.135
c27 2 VSS 0.0686416f $X=0.081 $Y=0.0675
r28 18 21 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.152
r29 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r30 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r31 5 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r32 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r33 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA31X2_ASAP7_75T_L%A2 2 5 8 11 13 18 19 20 21 25 VSS
c31 26 VSS 1.3589e-19 $X=0.176 $Y=0.135
c32 25 VSS 4.16237e-19 $X=0.163 $Y=0.135
c33 23 VSS 2.25678e-19 $X=0.189 $Y=0.135
c34 21 VSS 5.32335e-19 $X=0.144 $Y=0.135
c35 20 VSS 3.6486e-19 $X=0.135 $Y=0.1755
c36 19 VSS 5.97707e-19 $X=0.135 $Y=0.164
c37 18 VSS 0.0013246f $X=0.135 $Y=0.187
c38 11 VSS 0.00426697f $X=0.243 $Y=0.135
c39 8 VSS 0.0687639f $X=0.243 $Y=0.0675
c40 2 VSS 0.0641408f $X=0.189 $Y=0.135
r41 25 26 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.163
+ $Y=0.135 $X2=0.176 $Y2=0.135
r42 23 26 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.176 $Y2=0.135
r43 21 25 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.163 $Y2=0.135
r44 19 20 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.164 $X2=0.135 $Y2=0.1755
r45 18 20 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.187 $X2=0.135 $Y2=0.1755
r46 15 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.144 $X2=0.144 $Y2=0.135
r47 15 19 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.164
r48 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r49 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r50 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r51 2 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r52 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
.ends

.subckt PM_OA31X2_ASAP7_75T_L%A3 2 5 8 11 13 16 17 18 19 23 24 27 VSS
c28 27 VSS 6.76746e-19 $X=0.351 $Y=0.08
c29 24 VSS 1.01268e-19 $X=0.387 $Y=0.135
c30 23 VSS 5.53318e-19 $X=0.369 $Y=0.135
c31 21 VSS 3.59555e-19 $X=0.405 $Y=0.135
c32 19 VSS 0.00216903f $X=0.36 $Y=0.135
c33 18 VSS 9.9711e-20 $X=0.351 $Y=0.106
c34 17 VSS 3.57166e-19 $X=0.351 $Y=0.099
c35 16 VSS 9.08616e-19 $X=0.351 $Y=0.126
c36 11 VSS 0.00464802f $X=0.459 $Y=0.135
c37 8 VSS 0.0638058f $X=0.459 $Y=0.0675
c38 2 VSS 0.0690393f $X=0.405 $Y=0.135
r39 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.369
+ $Y=0.135 $X2=0.387 $Y2=0.135
r40 21 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.387 $Y2=0.135
r41 19 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.135 $X2=0.369 $Y2=0.135
r42 17 18 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.099 $X2=0.351 $Y2=0.106
r43 16 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.351 $Y=0.126 $X2=0.36 $Y2=0.135
r44 16 18 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.106
r45 15 27 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.072
r46 15 17 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.099
r47 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r48 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r49 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r50 2 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r51 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
.ends

.subckt PM_OA31X2_ASAP7_75T_L%B1 2 5 7 11 VSS
c15 11 VSS 0.0018203f $X=0.515 $Y=0.129
c16 5 VSS 0.00153111f $X=0.513 $Y=0.135
c17 2 VSS 0.0635225f $X=0.513 $Y=0.0675
r18 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r19 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.216
r20 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OA31X2_ASAP7_75T_L%7 1 2 6 11 14 17 19 21 24 26 29 31 34 36 39 42 43
+ 49 57 59 60 61 62 63 64 74 75 76 77 78 85 86 88 90 92 94 100 VSS
c86 100 VSS 1.91207e-19 $X=0.567 $Y=0.135
c87 97 VSS 0.00623377f $X=0.658 $Y=0.135
c88 94 VSS 0.00136805f $X=0.567 $Y=0.189
c89 92 VSS 4.94726e-19 $X=0.567 $Y=0.116
c90 91 VSS 0.00107686f $X=0.567 $Y=0.106
c91 90 VSS 3.57084e-19 $X=0.567 $Y=0.126
c92 88 VSS 5.31938e-19 $X=0.522 $Y=0.072
c93 87 VSS 1.63228e-19 $X=0.504 $Y=0.072
c94 86 VSS 6.49027e-20 $X=0.5 $Y=0.072
c95 85 VSS 6.60306e-19 $X=0.485 $Y=0.072
c96 80 VSS 0.00575401f $X=0.558 $Y=0.072
c97 79 VSS 0.00254755f $X=0.54 $Y=0.198
c98 78 VSS 0.00112812f $X=0.522 $Y=0.198
c99 77 VSS 0.00157938f $X=0.485 $Y=0.198
c100 76 VSS 1.67719e-19 $X=0.446 $Y=0.198
c101 75 VSS 1.10658e-19 $X=0.418 $Y=0.198
c102 74 VSS 7.12916e-20 $X=0.414 $Y=0.198
c103 66 VSS 0.0041777f $X=0.558 $Y=0.198
c104 64 VSS 3.3307e-19 $X=0.2365 $Y=0.072
c105 63 VSS 7.67329e-19 $X=0.203 $Y=0.072
c106 61 VSS 3.85413e-19 $X=0.126 $Y=0.072
c107 60 VSS 1.62371e-19 $X=0.094 $Y=0.072
c108 59 VSS 0.0010945f $X=0.09 $Y=0.072
c109 57 VSS 7.01881e-19 $X=0.27 $Y=0.072
c110 51 VSS 0.00171742f $X=0.054 $Y=0.072
c111 49 VSS 0.00357911f $X=0.486 $Y=0.2025
c112 44 VSS 6.64591e-19 $X=0.486 $Y=0.2245
c113 39 VSS 0.00311767f $X=0.38 $Y=0.2025
c114 36 VSS 3.2378e-19 $X=0.395 $Y=0.2025
c115 34 VSS 0.00289631f $X=0.434 $Y=0.0675
c116 31 VSS 4.59584e-19 $X=0.449 $Y=0.0675
c117 29 VSS 0.00310983f $X=0.268 $Y=0.0675
c118 24 VSS 9.0472e-19 $X=0.056 $Y=0.0675
c119 21 VSS 3.98338e-19 $X=0.071 $Y=0.0675
c120 17 VSS 0.00761819f $X=0.729 $Y=0.135
c121 14 VSS 0.0647446f $X=0.729 $Y=0.0675
c122 6 VSS 0.0657438f $X=0.675 $Y=0.0675
c123 2 VSS 1.751e-19 $X=0.282 $Y=0.096
c124 1 VSS 0.116569f $X=0.42 $Y=0.096
r125 97 98 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.658 $Y=0.135 $X2=0.658
+ $Y2=0.135
r126 95 100 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.135 $X2=0.567 $Y2=0.135
r127 95 97 5.5679 $w=1.8e-08 $l=8.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.135 $X2=0.658 $Y2=0.135
r128 93 100 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.144 $X2=0.567 $Y2=0.135
r129 93 94 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.144 $X2=0.567 $Y2=0.189
r130 91 92 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.106 $X2=0.567 $Y2=0.116
r131 90 100 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.126 $X2=0.567 $Y2=0.135
r132 90 92 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.126 $X2=0.567 $Y2=0.116
r133 89 91 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.567 $Y2=0.106
r134 87 88 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.072 $X2=0.522 $Y2=0.072
r135 86 87 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.5
+ $Y=0.072 $X2=0.504 $Y2=0.072
r136 85 86 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.485
+ $Y=0.072 $X2=0.5 $Y2=0.072
r137 82 85 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.072 $X2=0.485 $Y2=0.072
r138 80 89 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.072 $X2=0.567 $Y2=0.081
r139 80 88 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.072 $X2=0.522 $Y2=0.072
r140 78 79 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.198 $X2=0.54 $Y2=0.198
r141 76 77 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.446
+ $Y=0.198 $X2=0.485 $Y2=0.198
r142 75 76 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.198 $X2=0.446 $Y2=0.198
r143 74 75 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.418 $Y2=0.198
r144 72 78 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.198 $X2=0.522 $Y2=0.198
r145 72 77 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.198 $X2=0.485 $Y2=0.198
r146 68 74 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.198 $X2=0.414 $Y2=0.198
r147 66 94 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.198 $X2=0.567 $Y2=0.189
r148 66 79 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.198 $X2=0.54 $Y2=0.198
r149 63 64 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.203
+ $Y=0.072 $X2=0.2365 $Y2=0.072
r150 62 63 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.203 $Y2=0.072
r151 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.144 $Y2=0.072
r152 60 61 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.072 $X2=0.126 $Y2=0.072
r153 59 60 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.094 $Y2=0.072
r154 57 64 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.072 $X2=0.2365 $Y2=0.072
r155 51 59 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.072 $X2=0.09 $Y2=0.072
r156 49 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.198
+ $X2=0.486 $Y2=0.198
r157 43 44 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2245 $X2=0.486 $Y2=0.2245
r158 42 44 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.2245 $X2=0.486 $Y2=0.2245
r159 41 49 3.12934 $w=6.1e-08 $l=5.18073e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.486 $Y=0.206 $X2=0.469 $Y2=0.162
r160 41 44 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.486 $Y=0.206 $X2=0.486 $Y2=0.2245
r161 39 68 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.198
+ $X2=0.378 $Y2=0.198
r162 36 39 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.38 $Y2=0.2025
r163 34 82 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.072
+ $X2=0.432 $Y2=0.072
r164 31 34 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.434 $Y2=0.0675
r165 29 57 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.072 $X2=0.27
+ $Y2=0.072
r166 26 29 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.268 $Y2=0.0675
r167 24 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.072
+ $X2=0.054 $Y2=0.072
r168 21 24 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r169 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.135 $X2=0.729 $Y2=0.2025
r170 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.135
r171 9 17 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.729 $Y2=0.135
r172 9 98 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.658 $Y2=0.135
r173 9 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.2025
r174 6 9 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0675 $X2=0.675 $Y2=0.135
r175 4 34 14.2411 $w=2.4e-08 $l=1.65e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.084 $X2=0.432 $Y2=0.0675
r176 3 29 14.2411 $w=2.4e-08 $l=1.65e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.084 $X2=0.27 $Y2=0.0675
r177 2 3 11.5737 $w=2.4e-08 $l=1.69706e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.282 $Y=0.096 $X2=0.27 $Y2=0.084
r178 1 4 11.5737 $w=2.4e-08 $l=1.69706e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.42 $Y=0.096 $X2=0.432 $Y2=0.084
r179 1 2 119.107 $w=2.4e-08 $l=1.38e-07 $layer=LISD $thickness=2.8e-08 $X=0.42
+ $Y=0.096 $X2=0.282 $Y2=0.096
.ends

.subckt PM_OA31X2_ASAP7_75T_L%Y 1 2 6 7 10 11 14 16 24 29 VSS
c10 30 VSS 4.55454e-19 $X=0.783 $Y=0.216
c11 29 VSS 0.00406188f $X=0.783 $Y=0.207
c12 28 VSS 9.66845e-19 $X=0.783 $Y=0.144
c13 26 VSS 0.00207169f $X=0.783 $Y=0.09325
c14 25 VSS 8.85605e-19 $X=0.783 $Y=0.063
c15 24 VSS 0.00220141f $X=0.787 $Y=0.1235
c16 22 VSS 4.30151e-19 $X=0.783 $Y=0.225
c17 16 VSS 0.0141498f $X=0.774 $Y=0.234
c18 14 VSS 0.00966802f $X=0.702 $Y=0.036
c19 11 VSS 0.0139611f $X=0.774 $Y=0.036
c20 10 VSS 0.0095999f $X=0.702 $Y=0.2025
c21 6 VSS 5.945e-19 $X=0.719 $Y=0.2025
c22 1 VSS 5.945e-19 $X=0.719 $Y=0.0675
r23 29 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.207 $X2=0.783 $Y2=0.216
r24 28 29 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.144 $X2=0.783 $Y2=0.207
r25 27 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.126 $X2=0.783 $Y2=0.144
r26 25 26 2.05401 $w=1.8e-08 $l=3.025e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.063 $X2=0.783 $Y2=0.09325
r27 24 27 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.1235 $X2=0.783 $Y2=0.126
r28 24 26 2.05401 $w=1.8e-08 $l=3.025e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.1235 $X2=0.783 $Y2=0.09325
r29 22 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.225 $X2=0.783 $Y2=0.216
r30 21 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.063
r31 16 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.774 $Y=0.234 $X2=0.783 $Y2=0.225
r32 16 18 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.234 $X2=0.702 $Y2=0.234
r33 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.036 $X2=0.702
+ $Y2=0.036
r34 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.774 $Y=0.036 $X2=0.783 $Y2=0.045
r35 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.036 $X2=0.702 $Y2=0.036
r36 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.234 $X2=0.702
+ $Y2=0.234
r37 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2025 $X2=0.702 $Y2=0.2025
r38 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2025 $X2=0.702 $Y2=0.2025
r39 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.702
+ $Y=0.0675 $X2=0.702 $Y2=0.036
r40 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.685
+ $Y=0.0675 $X2=0.702 $Y2=0.0675
r41 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0675 $X2=0.702 $Y2=0.0675
.ends


* END of "./OA31x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA31x2_ASAP7_75t_L  VSS VDD A1 A2 A3 B1 Y
* 
* Y	Y
* B1	B1
* A3	A3
* A2	A2
* A1	A1
M0 noxref_9 N_A1_M0_g N_7_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_7_M1_d N_A2_M1_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M2 noxref_9 N_A3_M2_g N_7_M2_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M3 VSS N_B1_M3_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M4 N_Y_M4_d N_7_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665 $Y=0.027
M5 N_Y_M5_d N_7_M5_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M6 VDD N_A1_M6_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 VDD N_A1_M7_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 noxref_10 N_A2_M8_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 noxref_10 N_A2_M9_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 noxref_10 N_A3_M10_g N_7_M10_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M11 noxref_10 N_A3_M11_g N_7_M11_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M12 VDD N_B1_M12_g N_7_M12_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.503
+ $Y=0.189
M13 N_Y_M13_d N_7_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
M14 N_Y_M14_d N_7_M14_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
*
* 
* .include "OA31x2_ASAP7_75t_L.pex.sp.OA31X2_ASAP7_75T_L.pxi"
* BEGIN of "./OA31x2_ASAP7_75t_L.pex.sp.OA31X2_ASAP7_75T_L.pxi"
* File: OA31x2_ASAP7_75t_L.pex.sp.OA31X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:49:11 2017
* 
x_PM_OA31X2_ASAP7_75T_L%A1 N_A1_M0_g N_A1_M6_g N_A1_c_2_p N_A1_M7_g N_A1_c_7_p
+ A1 VSS PM_OA31X2_ASAP7_75T_L%A1
x_PM_OA31X2_ASAP7_75T_L%A2 N_A2_c_25_n N_A2_M8_g N_A2_M1_g N_A2_c_28_n N_A2_M9_g
+ A2 N_A2_c_30_n N_A2_c_32_n N_A2_c_33_n N_A2_c_35_n VSS
+ PM_OA31X2_ASAP7_75T_L%A2
x_PM_OA31X2_ASAP7_75T_L%A3 N_A3_c_56_p N_A3_M10_g N_A3_M2_g N_A3_c_58_p
+ N_A3_M11_g N_A3_c_59_p N_A3_c_63_p N_A3_c_64_p N_A3_c_82_p N_A3_c_65_p
+ N_A3_c_70_p A3 VSS PM_OA31X2_ASAP7_75T_L%A3
x_PM_OA31X2_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_86_n N_B1_M12_g B1 VSS
+ PM_OA31X2_ASAP7_75T_L%B1
x_PM_OA31X2_ASAP7_75T_L%7 N_7_c_109_n N_7_c_136_p N_7_M4_g N_7_M13_g N_7_M5_g
+ N_7_c_124_n N_7_M14_g N_7_M0_s N_7_c_99_n N_7_M1_d N_7_c_142_p N_7_M2_s
+ N_7_c_145_p N_7_M10_s N_7_c_137_p N_7_M12_s N_7_M11_s N_7_c_125_n N_7_c_104_n
+ N_7_c_100_n N_7_c_102_n N_7_c_138_p N_7_c_103_n N_7_c_106_n N_7_c_139_p
+ N_7_c_117_n N_7_c_170_p N_7_c_162_p N_7_c_120_n N_7_c_126_n N_7_c_121_n
+ N_7_c_128_n N_7_c_129_n N_7_c_131_n N_7_c_132_n N_7_c_133_n N_7_c_134_n VSS
+ PM_OA31X2_ASAP7_75T_L%7
x_PM_OA31X2_ASAP7_75T_L%Y N_Y_M5_d N_Y_M4_d N_Y_M14_d N_Y_M13_d N_Y_c_187_n
+ N_Y_c_188_n N_Y_c_190_n N_Y_c_191_n Y N_Y_c_194_n VSS PM_OA31X2_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_c_25_n 2.74891e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_2 N_A1_c_2_p N_A2_c_25_n 0.00372052f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_3 N_A1_c_2_p N_A2_M1_g 3.09654e-19 $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_4 N_A1_c_2_p N_A2_c_28_n 0.00153175f $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_5 A1 A2 0.0010886f $X=0.083 $Y=0.152 $X2=0.135 $Y2=0.187
cc_6 N_A1_c_2_p N_A2_c_30_n 4.68709e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.164
cc_7 N_A1_c_7_p N_A2_c_30_n 0.0010886f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.164
cc_8 N_A1_c_7_p N_A2_c_32_n 0.0010886f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.1755
cc_9 N_A1_c_2_p N_A2_c_33_n 0.0018007f $X=0.135 $Y=0.135 $X2=0.144 $Y2=0.135
cc_10 N_A1_c_7_p N_A2_c_33_n 0.0010886f $X=0.081 $Y=0.135 $X2=0.144 $Y2=0.135
cc_11 N_A1_c_2_p N_A2_c_35_n 4.61613e-19 $X=0.135 $Y=0.135 $X2=0.163 $Y2=0.135
cc_12 N_A1_c_7_p N_7_c_99_n 0.00117083f $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_13 N_A1_M0_g N_7_c_100_n 3.37536e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_14 N_A1_c_7_p N_7_c_100_n 0.00371968f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_15 N_A1_c_2_p N_7_c_102_n 5.39927e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_16 N_A1_c_2_p N_7_c_103_n 2.76185e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_17 VSS N_A1_c_7_p 4.92442e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_18 VSS A1 0.00179861f $X=0.083 $Y=0.152 $X2=0.189 $Y2=0.2025
cc_19 VSS N_A1_M0_g 2.34993e-19 $X=0.081 $Y=0.0675 $X2=0.163 $Y2=0.135
cc_20 VSS A1 0.00372137f $X=0.083 $Y=0.152 $X2=0.163 $Y2=0.135
cc_21 VSS N_A1_c_2_p 5.90915e-19 $X=0.135 $Y=0.135 $X2=0.176 $Y2=0.135
cc_22 VSS N_A1_c_2_p 2.34993e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_23 VSS N_A1_c_2_p 8.0006e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.187
cc_24 VSS N_A1_c_2_p 2.38303e-19 $X=0.135 $Y=0.135 $X2=0.176 $Y2=0.135
cc_25 N_A2_M1_g N_7_c_104_n 3.09722e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_A2_c_33_n N_7_c_103_n 0.00123353f $X=0.144 $Y=0.135 $X2=0 $Y2=0
cc_27 N_A2_c_25_n N_7_c_106_n 3.31725e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_28 N_A2_c_28_n N_7_c_106_n 7.60145e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_29 N_A2_c_35_n N_7_c_106_n 0.00209283f $X=0.163 $Y=0.135 $X2=0 $Y2=0
cc_30 VSS A2 0.00109041f $X=0.135 $Y=0.187 $X2=0.135 $Y2=0.135
cc_31 VSS N_A2_c_30_n 5.14282e-19 $X=0.135 $Y=0.164 $X2=0.135 $Y2=0.135
cc_32 VSS N_A2_M1_g 2.64781e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_33 VSS A2 0.00373885f $X=0.135 $Y=0.187 $X2=0.135 $Y2=0.135
cc_34 VSS N_A2_c_25_n 4.28653e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_35 VSS N_A2_c_35_n 7.32095e-19 $X=0.163 $Y=0.135 $X2=0 $Y2=0
cc_36 VSS N_A2_c_28_n 8.0006e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_37 VSS N_A2_c_25_n 2.64781e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_38 VSS N_A2_M1_g 2.64781e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_39 VSS N_A2_c_35_n 2.51638e-19 $X=0.163 $Y=0.135 $X2=0 $Y2=0
cc_40 VSS N_A2_c_28_n 3.8028e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_41 VSS N_A2_c_28_n 8.0006e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_42 VSS N_A2_c_28_n 6.91613e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_43 VSS A2 6.78462e-19 $X=0.135 $Y=0.187 $X2=0.135 $Y2=0.2025
cc_44 VSS N_A2_M1_g 3.99641e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_45 N_A3_c_56_p N_B1_M3_g 3.03912e-19 $X=0.405 $Y=0.135 $X2=0.189 $Y2=0.135
cc_46 N_A3_M2_g N_B1_M3_g 0.00359705f $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_47 N_A3_c_58_p N_B1_c_86_n 0.00130224f $X=0.459 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_48 N_A3_c_59_p B1 2.06743e-19 $X=0.351 $Y=0.126 $X2=0.243 $Y2=0.135
cc_49 N_A3_c_56_p N_7_c_109_n 0.00265807f $X=0.405 $Y=0.135 $X2=0.189 $Y2=0.135
cc_50 N_A3_c_58_p N_7_c_109_n 0.00132216f $X=0.459 $Y=0.135 $X2=0.189 $Y2=0.135
cc_51 N_A3_c_59_p N_7_c_109_n 7.47901e-19 $X=0.351 $Y=0.126 $X2=0.189 $Y2=0.135
cc_52 N_A3_c_63_p N_7_c_109_n 0.00117454f $X=0.351 $Y=0.099 $X2=0.189 $Y2=0.135
cc_53 N_A3_c_64_p N_7_c_109_n 5.47014e-19 $X=0.351 $Y=0.106 $X2=0.189 $Y2=0.135
cc_54 N_A3_c_65_p N_7_c_109_n 5.91517e-19 $X=0.369 $Y=0.135 $X2=0.189 $Y2=0.135
cc_55 A3 N_7_c_109_n 8.77807e-19 $X=0.351 $Y=0.08 $X2=0.189 $Y2=0.135
cc_56 A3 N_7_c_104_n 9.31566e-19 $X=0.351 $Y=0.08 $X2=0 $Y2=0
cc_57 N_A3_c_56_p N_7_c_117_n 3.19976e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_58 N_A3_c_58_p N_7_c_117_n 8.65402e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_59 N_A3_c_70_p N_7_c_117_n 0.00144344f $X=0.387 $Y=0.135 $X2=0 $Y2=0
cc_60 N_A3_M2_g N_7_c_120_n 4.89074e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_61 N_A3_M2_g N_7_c_121_n 3.93692e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_62 N_A3_c_58_p N_7_c_121_n 6.97968e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_63 A3 N_7_c_121_n 6.15281e-19 $X=0.351 $Y=0.08 $X2=0 $Y2=0
cc_64 VSS N_A3_M2_g 2.21754e-19 $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_65 VSS A3 0.00360338f $X=0.351 $Y=0.08 $X2=0 $Y2=0
cc_66 VSS N_A3_c_56_p 3.58882e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_67 VSS N_A3_c_65_p 9.39365e-19 $X=0.369 $Y=0.135 $X2=0 $Y2=0
cc_68 VSS N_A3_c_58_p 3.80246e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_69 VSS N_A3_c_58_p 8.0006e-19 $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.135
cc_70 VSS A3 2.80639e-19 $X=0.351 $Y=0.08 $X2=0.243 $Y2=0.135
cc_71 VSS N_A3_c_82_p 5.57567e-19 $X=0.36 $Y=0.135 $X2=0 $Y2=0
cc_72 VSS N_A3_c_65_p 2.35337e-19 $X=0.369 $Y=0.135 $X2=0 $Y2=0
cc_73 N_B1_c_86_n N_7_c_124_n 2.02195e-19 $X=0.513 $Y=0.135 $X2=0.351 $Y2=0.099
cc_74 B1 N_7_c_125_n 9.02364e-19 $X=0.515 $Y=0.129 $X2=0 $Y2=0
cc_75 N_B1_M3_g N_7_c_126_n 3.37536e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_76 B1 N_7_c_126_n 0.00373829f $X=0.515 $Y=0.129 $X2=0 $Y2=0
cc_77 B1 N_7_c_128_n 4.10939e-19 $X=0.515 $Y=0.129 $X2=0 $Y2=0
cc_78 N_B1_M3_g N_7_c_129_n 3.62029e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_79 B1 N_7_c_129_n 0.00122403f $X=0.515 $Y=0.129 $X2=0 $Y2=0
cc_80 B1 N_7_c_131_n 8.14929e-19 $X=0.515 $Y=0.129 $X2=0 $Y2=0
cc_81 B1 N_7_c_132_n 8.14929e-19 $X=0.515 $Y=0.129 $X2=0 $Y2=0
cc_82 B1 N_7_c_133_n 8.14929e-19 $X=0.515 $Y=0.129 $X2=0 $Y2=0
cc_83 B1 N_7_c_134_n 8.14929e-19 $X=0.515 $Y=0.129 $X2=0 $Y2=0
cc_84 VSS N_7_c_99_n 0.00134615f $X=0.056 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_85 VSS N_7_c_136_p 0.00151902f $X=0.282 $Y=0.096 $X2=0 $Y2=0
cc_86 VSS N_7_c_137_p 0.00138889f $X=0.38 $Y=0.2025 $X2=0 $Y2=0
cc_87 VSS N_7_c_138_p 3.00265e-19 $X=0.126 $Y=0.072 $X2=0.081 $Y2=0.135
cc_88 VSS N_7_c_139_p 3.29233e-19 $X=0.2365 $Y=0.072 $X2=0.081 $Y2=0.2025
cc_89 VSS N_7_c_99_n 0.00343094f $X=0.056 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_90 VSS N_7_c_138_p 0.00262229f $X=0.126 $Y=0.072 $X2=0.081 $Y2=0.135
cc_91 VSS N_7_c_142_p 0.00355213f $X=0.268 $Y=0.0675 $X2=0 $Y2=0
cc_92 VSS N_7_c_139_p 0.00255088f $X=0.2365 $Y=0.072 $X2=0 $Y2=0
cc_93 VSS N_7_c_128_n 0.00353488f $X=0.5 $Y=0.072 $X2=0 $Y2=0
cc_94 VSS N_7_c_145_p 0.00359031f $X=0.434 $Y=0.0675 $X2=0 $Y2=0
cc_95 VSS N_7_c_125_n 0.00149296f $X=0.486 $Y=0.2025 $X2=0 $Y2=0
cc_96 VSS N_7_c_121_n 0.00107804f $X=0.485 $Y=0.072 $X2=0 $Y2=0
cc_97 VSS N_7_c_128_n 0.001169f $X=0.5 $Y=0.072 $X2=0 $Y2=0
cc_98 VSS N_7_c_136_p 2.88467e-19 $X=0.282 $Y=0.096 $X2=0 $Y2=0
cc_99 VSS N_7_c_99_n 3.09693e-19 $X=0.056 $Y=0.0675 $X2=0 $Y2=0
cc_100 VSS N_7_c_142_p 0.00291007f $X=0.268 $Y=0.0675 $X2=0 $Y2=0
cc_101 VSS N_7_c_138_p 0.0157549f $X=0.126 $Y=0.072 $X2=0 $Y2=0
cc_102 VSS N_7_c_109_n 8.14546e-19 $X=0.42 $Y=0.096 $X2=0 $Y2=0
cc_103 VSS N_7_c_109_n 0.00121499f $X=0.42 $Y=0.096 $X2=0 $Y2=0
cc_104 VSS N_7_c_109_n 2.88467e-19 $X=0.42 $Y=0.096 $X2=0 $Y2=0
cc_105 VSS N_7_M2_s 3.16747e-19 $X=0.449 $Y=0.0675 $X2=0 $Y2=0
cc_106 VSS N_7_c_145_p 0.00259595f $X=0.434 $Y=0.0675 $X2=0 $Y2=0
cc_107 VSS N_7_c_121_n 0.00353488f $X=0.485 $Y=0.072 $X2=0 $Y2=0
cc_108 VSS N_7_c_109_n 0.00151902f $X=0.42 $Y=0.096 $X2=0.135 $Y2=0.135
cc_109 VSS N_7_c_137_p 0.0035285f $X=0.38 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_110 VSS N_7_c_125_n 0.00328965f $X=0.486 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_111 VSS N_7_c_162_p 0.00226064f $X=0.446 $Y=0.198 $X2=0.135 $Y2=0.135
cc_112 VSS N_7_c_137_p 5.61679e-19 $X=0.38 $Y=0.2025 $X2=0 $Y2=0
cc_113 VSS N_7_c_117_n 9.95918e-19 $X=0.414 $Y=0.198 $X2=0 $Y2=0
cc_114 VSS N_7_c_106_n 2.38776e-19 $X=0.203 $Y=0.072 $X2=0.135 $Y2=0.2025
cc_115 VSS N_7_c_139_p 2.38776e-19 $X=0.2365 $Y=0.072 $X2=0.135 $Y2=0.2025
cc_116 VSS N_7_c_109_n 9.15892e-19 $X=0.42 $Y=0.096 $X2=0.081 $Y2=0.135
cc_117 VSS N_7_c_104_n 2.38776e-19 $X=0.27 $Y=0.072 $X2=0.081 $Y2=0.135
cc_118 VSS N_7_c_125_n 3.13327e-19 $X=0.486 $Y=0.2025 $X2=0 $Y2=0
cc_119 VSS N_7_c_170_p 0.0031969f $X=0.418 $Y=0.198 $X2=0 $Y2=0
cc_120 VSS N_7_c_137_p 8.27072e-19 $X=0.38 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_121 VSS N_7_M10_s 3.12293e-19 $X=0.395 $Y=0.2025 $X2=0 $Y2=0
cc_122 VSS N_7_c_137_p 0.0019103f $X=0.38 $Y=0.2025 $X2=0 $Y2=0
cc_123 VSS N_7_c_117_n 0.0031969f $X=0.414 $Y=0.198 $X2=0 $Y2=0
cc_124 N_7_c_124_n N_Y_M5_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_125 N_7_c_124_n N_Y_M14_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_126 N_7_c_124_n N_Y_c_187_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.135 $Y2=0.135
cc_127 N_7_M5_g N_Y_c_188_n 4.59284e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_128 N_7_c_124_n N_Y_c_188_n 4.80361e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_129 N_7_c_124_n N_Y_c_190_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_130 N_7_M5_g N_Y_c_191_n 4.59284e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_131 N_7_c_124_n N_Y_c_191_n 4.80361e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_132 N_7_c_124_n Y 5.0726e-19 $X=0.729 $Y=0.135 $X2=0 $Y2=0
cc_133 N_7_c_133_n N_Y_c_194_n 2.15381e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0

* END of "./OA31x2_ASAP7_75t_L.pex.sp.OA31X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA331x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:49:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA331x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA331x1_ASAP7_75t_L.pex.sp.pex"
* File: OA331x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:49:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA331X1_ASAP7_75T_L%3 2 5 7 9 12 14 15 18 19 22 26 30 32 34 39 41 42
+ 43 44 45 49 50 51 52 53 55 58 64 67 76 VSS
c43 76 VSS 0.00202532f $X=0.504 $Y=0.072
c44 75 VSS 0.00163302f $X=0.513 $Y=0.072
c45 69 VSS 6.57651e-19 $X=0.099 $Y=0.195
c46 68 VSS 6.23446e-19 $X=0.09 $Y=0.195
c47 67 VSS 0.00204357f $X=0.108 $Y=0.195
c48 64 VSS 0.00412141f $X=0.513 $Y=0.2
c49 63 VSS 0.00103118f $X=0.513 $Y=0.106
c50 62 VSS 8.11244e-19 $X=0.513 $Y=0.225
c51 60 VSS 6.94247e-19 $X=0.4785 $Y=0.234
c52 59 VSS 2.39163e-19 $X=0.471 $Y=0.234
c53 58 VSS 0.00146362f $X=0.468 $Y=0.234
c54 57 VSS 2.39163e-19 $X=0.45 $Y=0.234
c55 56 VSS 0.00617212f $X=0.447 $Y=0.234
c56 55 VSS 0.00142296f $X=0.414 $Y=0.234
c57 54 VSS 3.71649e-19 $X=0.396 $Y=0.234
c58 53 VSS 0.00311761f $X=0.393 $Y=0.234
c59 52 VSS 0.00146362f $X=0.36 $Y=0.234
c60 51 VSS 0.00340162f $X=0.342 $Y=0.234
c61 50 VSS 0.00146362f $X=0.306 $Y=0.234
c62 49 VSS 0.00256536f $X=0.288 $Y=0.234
c63 45 VSS 8.84964e-19 $X=0.261 $Y=0.234
c64 44 VSS 0.00142296f $X=0.252 $Y=0.234
c65 43 VSS 0.00360252f $X=0.234 $Y=0.234
c66 42 VSS 0.00142296f $X=0.198 $Y=0.234
c67 41 VSS 0.00312977f $X=0.18 $Y=0.234
c68 40 VSS 3.78291e-19 $X=0.148 $Y=0.234
c69 39 VSS 0.00151377f $X=0.144 $Y=0.234
c70 38 VSS 0.00171948f $X=0.126 $Y=0.234
c71 34 VSS 0.00330057f $X=0.117 $Y=0.234
c72 33 VSS 0.00590321f $X=0.504 $Y=0.234
c73 32 VSS 0.00229578f $X=0.108 $Y=0.225
c74 30 VSS 4.04879e-19 $X=0.081 $Y=0.176
c75 26 VSS 7.04746e-19 $X=0.081 $Y=0.135
c76 24 VSS 3.84635e-19 $X=0.081 $Y=0.186
c77 22 VSS 0.00701741f $X=0.484 $Y=0.2025
c78 18 VSS 0.00220219f $X=0.27 $Y=0.2025
c79 14 VSS 5.38922e-19 $X=0.287 $Y=0.2025
c80 12 VSS 0.0013176f $X=0.484 $Y=0.0675
c81 5 VSS 0.0024241f $X=0.081 $Y=0.135
c82 2 VSS 0.0649339f $X=0.081 $Y=0.0675
r83 76 77 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.072 $X2=0.5085 $Y2=0.072
r84 75 77 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.072 $X2=0.5085 $Y2=0.072
r85 72 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.072 $X2=0.504 $Y2=0.072
r86 68 69 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.195 $X2=0.099 $Y2=0.195
r87 67 69 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.195 $X2=0.099 $Y2=0.195
r88 65 68 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.195 $X2=0.09 $Y2=0.195
r89 63 64 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.106 $X2=0.513 $Y2=0.2
r90 62 64 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.2
r91 61 75 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.081 $X2=0.513 $Y2=0.072
r92 61 63 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.081 $X2=0.513 $Y2=0.106
r93 59 60 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.471
+ $Y=0.234 $X2=0.4785 $Y2=0.234
r94 58 59 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.471 $Y2=0.234
r95 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r96 56 57 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.234 $X2=0.45 $Y2=0.234
r97 55 56 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.447 $Y2=0.234
r98 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r99 53 54 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.393
+ $Y=0.234 $X2=0.396 $Y2=0.234
r100 52 53 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.393 $Y2=0.234
r101 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r102 50 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.342 $Y2=0.234
r103 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r104 47 60 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.4785 $Y2=0.234
r105 44 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.261 $Y2=0.234
r106 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r107 42 43 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.234 $Y2=0.234
r108 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r109 40 41 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.234 $X2=0.18 $Y2=0.234
r110 39 40 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.148 $Y2=0.234
r111 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r112 36 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.288 $Y2=0.234
r113 36 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.261 $Y2=0.234
r114 34 38 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.234 $X2=0.126 $Y2=0.234
r115 33 62 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.234 $X2=0.513 $Y2=0.225
r116 33 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.486 $Y2=0.234
r117 32 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.108 $Y=0.225 $X2=0.117 $Y2=0.234
r118 31 67 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.204 $X2=0.108 $Y2=0.195
r119 31 32 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.204 $X2=0.108 $Y2=0.225
r120 29 30 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.166 $X2=0.081 $Y2=0.176
r121 26 29 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.166
r122 24 65 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.186 $X2=0.081 $Y2=0.195
r123 24 30 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.186 $X2=0.081 $Y2=0.176
r124 22 47 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234
+ $X2=0.486 $Y2=0.234
r125 19 22 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.484 $Y2=0.2025
r126 18 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r127 15 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r128 14 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r129 12 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.072
+ $X2=0.486 $Y2=0.072
r130 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.484 $Y2=0.0675
r131 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r132 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r133 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA331X1_ASAP7_75T_L%A3 2 5 7 10 18 VSS
c11 10 VSS 0.0027483f $X=0.135 $Y=0.135
c12 5 VSS 0.001273f $X=0.135 $Y=0.135
c13 2 VSS 0.0593081f $X=0.135 $Y=0.0675
r14 10 18 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OA331X1_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c14 14 VSS 5.30982e-19 $X=0.189 $Y=0.155
c15 10 VSS 4.5987e-19 $X=0.189 $Y=0.135
c16 5 VSS 0.00110916f $X=0.189 $Y=0.135
c17 2 VSS 0.059482f $X=0.189 $Y=0.0675
r18 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.155
r19 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r20 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r21 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA331X1_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c12 10 VSS 4.82288e-19 $X=0.243 $Y=0.135
c13 5 VSS 0.00111383f $X=0.243 $Y=0.135
c14 2 VSS 0.060901f $X=0.243 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OA331X1_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.297 $Y=0.135
c14 5 VSS 0.00111336f $X=0.297 $Y=0.135
c15 2 VSS 0.0617786f $X=0.297 $Y=0.0675
r16 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.154
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OA331X1_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.351 $Y=0.135
c14 5 VSS 0.00112198f $X=0.351 $Y=0.135
c15 2 VSS 0.0616432f $X=0.351 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OA331X1_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c11 10 VSS 7.24259e-19 $X=0.405 $Y=0.135
c12 5 VSS 0.00113686f $X=0.405 $Y=0.135
c13 2 VSS 0.0618011f $X=0.405 $Y=0.0675
r14 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OA331X1_ASAP7_75T_L%C1 2 5 7 10 14 VSS
c8 10 VSS 0.00201948f $X=0.459 $Y=0.135
c9 5 VSS 0.00178699f $X=0.459 $Y=0.135
c10 2 VSS 0.0660367f $X=0.459 $Y=0.0675
r11 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.155
r12 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OA331X1_ASAP7_75T_L%Y 1 6 9 14 16 18 22 23 30 VSS
c7 33 VSS 9.17717e-19 $X=0.045 $Y=0.234
c8 32 VSS 0.0032947f $X=0.036 $Y=0.234
c9 30 VSS 0.0030586f $X=0.054 $Y=0.234
c10 25 VSS 9.17717e-19 $X=0.045 $Y=0.036
c11 24 VSS 0.0032947f $X=0.036 $Y=0.036
c12 23 VSS 0.0063623f $X=0.054 $Y=0.036
c13 22 VSS 0.00328209f $X=0.054 $Y=0.036
c14 18 VSS 3.56737e-19 $X=0.027 $Y=0.2145
c15 16 VSS 0.00201583f $X=0.027 $Y=0.115
c16 15 VSS 8.81034e-19 $X=0.027 $Y=0.07
c17 14 VSS 0.00385152f $X=0.03 $Y=0.143
c18 12 VSS 3.3975e-19 $X=0.027 $Y=0.225
c19 9 VSS 0.0067618f $X=0.056 $Y=0.2025
c20 6 VSS 3.7894e-19 $X=0.071 $Y=0.2025
c21 1 VSS 3.7894e-19 $X=0.071 $Y=0.0675
r22 32 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.045 $Y2=0.234
r23 30 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.045 $Y2=0.234
r24 27 32 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.036 $Y2=0.234
r25 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.045 $Y2=0.036
r26 22 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.045 $Y2=0.036
r27 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r28 19 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.036 $Y2=0.036
r29 17 18 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.204 $X2=0.027 $Y2=0.2145
r30 15 16 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.115
r31 14 17 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.143 $X2=0.027 $Y2=0.204
r32 14 16 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.143 $X2=0.027 $Y2=0.115
r33 12 27 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.234
r34 12 18 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.2145
r35 11 19 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.036
r36 11 15 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r37 9 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r38 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
r39 4 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r40 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./OA331x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA331x1_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C1 Y
* 
* Y	Y
* C1	C1
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 VSS N_3_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 noxref_12 N_A3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_A2_M2_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_12 N_A1_M3_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_13 N_B1_M4_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_12 N_B2_M5_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_13 N_B3_M6_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_3_M7_d N_C1_M7_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 VDD N_3_M8_g N_Y_M8_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M9 noxref_14 N_A3_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M10 noxref_15 N_A2_M10_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.179 $Y=0.162
M11 N_3_M11_d N_A1_M11_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M12 noxref_16 N_B1_M12_g N_3_M12_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M13 noxref_17 N_B2_M13_g noxref_16 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M14 VDD N_B3_M14_g noxref_17 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M15 N_3_M15_d N_C1_M15_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "OA331x1_ASAP7_75t_L.pex.sp.OA331X1_ASAP7_75T_L.pxi"
* BEGIN of "./OA331x1_ASAP7_75t_L.pex.sp.OA331X1_ASAP7_75T_L.pxi"
* File: OA331x1_ASAP7_75t_L.pex.sp.OA331X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:49:34 2017
* 
x_PM_OA331X1_ASAP7_75T_L%3 N_3_M0_g N_3_c_3_p N_3_M8_g N_3_M7_d N_3_c_37_p
+ N_3_M12_s N_3_M11_d N_3_c_12_p N_3_M15_d N_3_c_22_p N_3_c_4_p N_3_c_8_p
+ N_3_c_27_p N_3_c_28_p N_3_c_2_p N_3_c_31_p N_3_c_7_p N_3_c_30_p N_3_c_11_p
+ N_3_c_33_p N_3_c_34_p N_3_c_14_p N_3_c_35_p N_3_c_17_p N_3_c_36_p N_3_c_19_p
+ N_3_c_21_p N_3_c_24_p N_3_c_10_p N_3_c_32_p VSS PM_OA331X1_ASAP7_75T_L%3
x_PM_OA331X1_ASAP7_75T_L%A3 N_A3_M1_g N_A3_c_46_n N_A3_M9_g N_A3_c_47_n A3 VSS
+ PM_OA331X1_ASAP7_75T_L%A3
x_PM_OA331X1_ASAP7_75T_L%A2 N_A2_M2_g N_A2_c_61_n N_A2_M10_g N_A2_c_62_n A2 VSS
+ PM_OA331X1_ASAP7_75T_L%A2
x_PM_OA331X1_ASAP7_75T_L%A1 N_A1_M3_g N_A1_c_74_n N_A1_M11_g N_A1_c_70_n A1 VSS
+ PM_OA331X1_ASAP7_75T_L%A1
x_PM_OA331X1_ASAP7_75T_L%B1 N_B1_M4_g N_B1_c_86_n N_B1_M12_g N_B1_c_82_n B1 VSS
+ PM_OA331X1_ASAP7_75T_L%B1
x_PM_OA331X1_ASAP7_75T_L%B2 N_B2_M5_g N_B2_c_98_n N_B2_M13_g N_B2_c_95_n B2 VSS
+ PM_OA331X1_ASAP7_75T_L%B2
x_PM_OA331X1_ASAP7_75T_L%B3 N_B3_M6_g N_B3_c_111_n N_B3_M14_g N_B3_c_108_n B3
+ VSS PM_OA331X1_ASAP7_75T_L%B3
x_PM_OA331X1_ASAP7_75T_L%C1 N_C1_M7_g N_C1_c_124_n N_C1_M15_g N_C1_c_119_n C1
+ VSS PM_OA331X1_ASAP7_75T_L%C1
x_PM_OA331X1_ASAP7_75T_L%Y N_Y_M0_s N_Y_M8_s N_Y_c_126_n Y N_Y_c_130_n
+ N_Y_c_128_n N_Y_c_132_p N_Y_c_131_p N_Y_c_129_n VSS PM_OA331X1_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M1_g 0.00284417f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_3_c_2_p N_A3_M1_g 2.3886e-19 $X=0.144 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_3 N_3_c_3_p N_A3_c_46_n 9.34529e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_3_c_4_p N_A3_c_47_n 0.00221012f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_5 N_3_c_2_p N_A3_c_47_n 2.7862e-19 $X=0.144 $Y=0.234 $X2=0.135 $Y2=0.135
cc_6 N_3_M0_g N_A2_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_7 N_3_c_7_p N_A2_M2_g 3.38929e-19 $X=0.198 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_8 N_3_c_8_p A2 2.13942e-19 $X=0.081 $Y=0.176 $X2=0 $Y2=0
cc_9 N_3_c_7_p A2 0.00123064f $X=0.198 $Y=0.234 $X2=0 $Y2=0
cc_10 N_3_c_10_p A2 4.18335e-19 $X=0.108 $Y=0.195 $X2=0 $Y2=0
cc_11 N_3_c_11_p N_A1_M3_g 2.56935e-19 $X=0.252 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_12 N_3_c_12_p N_A1_c_70_n 0.0013295f $X=0.27 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_13 N_3_c_11_p N_A1_c_70_n 0.00123064f $X=0.252 $Y=0.234 $X2=0.135 $Y2=0.135
cc_14 N_3_c_14_p N_B1_M4_g 2.64276e-19 $X=0.306 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_15 N_3_c_12_p N_B1_c_82_n 0.0013295f $X=0.27 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_16 N_3_c_14_p N_B1_c_82_n 0.00124805f $X=0.306 $Y=0.234 $X2=0.135 $Y2=0.135
cc_17 N_3_c_17_p N_B2_M5_g 3.48613e-19 $X=0.36 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_18 N_3_c_17_p N_B2_c_95_n 0.00124805f $X=0.36 $Y=0.234 $X2=0.135 $Y2=0.135
cc_19 N_3_c_19_p N_B3_M6_g 2.56935e-19 $X=0.414 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_20 N_3_c_19_p N_B3_c_108_n 0.00123064f $X=0.414 $Y=0.234 $X2=0.135 $Y2=0.135
cc_21 N_3_c_21_p N_C1_M7_g 2.64276e-19 $X=0.468 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_22 N_3_c_22_p N_C1_c_119_n 0.00114532f $X=0.484 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_23 N_3_c_21_p N_C1_c_119_n 0.00124805f $X=0.468 $Y=0.234 $X2=0.135 $Y2=0.135
cc_24 N_3_c_24_p N_C1_c_119_n 0.00392202f $X=0.513 $Y=0.2 $X2=0.135 $Y2=0.135
cc_25 N_3_c_4_p N_Y_c_126_n 0.00125175f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_26 N_3_c_4_p Y 0.0036413f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_27 N_3_c_27_p N_Y_c_128_n 2.71869e-19 $X=0.108 $Y=0.225 $X2=0.135 $Y2=0.155
cc_28 N_3_c_28_p N_Y_c_129_n 9.13687e-19 $X=0.117 $Y=0.234 $X2=0 $Y2=0
cc_29 VSS N_3_c_12_p 0.00138157f $X=0.27 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_30 VSS N_3_c_30_p 2.20596e-19 $X=0.234 $Y=0.234 $X2=0 $Y2=0
cc_31 VSS N_3_c_31_p 2.20596e-19 $X=0.18 $Y=0.234 $X2=0 $Y2=0
cc_32 VSS N_3_c_32_p 2.82518e-19 $X=0.504 $Y=0.072 $X2=0 $Y2=0
cc_33 VSS N_3_c_33_p 2.23188e-19 $X=0.261 $Y=0.234 $X2=0 $Y2=0
cc_34 VSS N_3_c_34_p 2.23188e-19 $X=0.288 $Y=0.234 $X2=0 $Y2=0
cc_35 VSS N_3_c_35_p 2.23188e-19 $X=0.342 $Y=0.234 $X2=0 $Y2=0
cc_36 VSS N_3_c_36_p 2.23188e-19 $X=0.393 $Y=0.234 $X2=0 $Y2=0
cc_37 VSS N_3_c_37_p 3.11523e-19 $X=0.484 $Y=0.0675 $X2=0 $Y2=0
cc_38 VSS N_3_c_37_p 0.00333695f $X=0.484 $Y=0.0675 $X2=0.135 $Y2=0.155
cc_39 VSS N_3_c_32_p 4.47506e-19 $X=0.504 $Y=0.072 $X2=0.135 $Y2=0.155
cc_40 VSS N_3_c_31_p 3.25855e-19 $X=0.18 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_41 VSS N_3_c_30_p 3.56327e-19 $X=0.234 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_42 VSS N_3_c_35_p 3.48201e-19 $X=0.342 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_43 VSS N_3_c_36_p 3.30547e-19 $X=0.393 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_44 N_A3_M1_g N_A2_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_45 N_A3_c_46_n N_A2_c_61_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_46 N_A3_c_47_n N_A2_c_62_n 0.00286115f $X=0.135 $Y=0.135 $X2=0.484 $Y2=0.0675
cc_47 N_A3_M1_g N_A1_M3_g 2.66145e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_48 N_A3_c_47_n N_Y_c_130_n 4.26334e-19 $X=0.135 $Y=0.135 $X2=0.27 $Y2=0.2025
cc_49 VSS N_A3_c_47_n 8.88545e-19 $X=0.135 $Y=0.135 $X2=0.469 $Y2=0.2025
cc_50 N_A2_M2_g N_A1_M3_g 0.00327995f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_51 N_A2_c_61_n N_A1_c_74_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_52 N_A2_c_62_n N_A1_c_70_n 0.00482209f $X=0.189 $Y=0.135 $X2=0.484 $Y2=0.0675
cc_53 N_A2_M2_g N_B1_M4_g 2.71887e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_54 VSS N_A2_M2_g 3.57119e-19 $X=0.189 $Y=0.0675 $X2=0.484 $Y2=0.2025
cc_55 VSS N_A2_c_62_n 5.37372e-19 $X=0.189 $Y=0.135 $X2=0.484 $Y2=0.2025
cc_56 N_A1_M3_g N_B1_M4_g 0.0036939f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_57 N_A1_c_74_n N_B1_c_86_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_58 N_A1_c_70_n N_B1_c_82_n 0.00406615f $X=0.243 $Y=0.135 $X2=0.484 $Y2=0.0675
cc_59 N_A1_M3_g N_B2_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_60 VSS N_A1_c_70_n 0.00159458f $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_61 N_B1_M4_g N_B2_M5_g 0.00371573f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_62 N_B1_c_86_n N_B2_c_98_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_63 N_B1_c_82_n N_B2_c_95_n 0.00483372f $X=0.297 $Y=0.135 $X2=0.484 $Y2=0.0675
cc_64 N_B1_M4_g N_B3_M6_g 3.06651e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_65 VSS N_B1_M4_g 3.62029e-19 $X=0.297 $Y=0.0675 $X2=0.504 $Y2=0.234
cc_66 VSS N_B1_c_82_n 0.0012322f $X=0.297 $Y=0.135 $X2=0.504 $Y2=0.234
cc_67 N_B2_M5_g N_B3_M6_g 0.0036939f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_68 N_B2_c_98_n N_B3_c_111_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_69 N_B2_c_95_n N_B3_c_108_n 0.00483372f $X=0.351 $Y=0.135 $X2=0.484
+ $Y2=0.0675
cc_70 N_B2_M5_g N_C1_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_71 VSS N_B2_M5_g 2.68514e-19 $X=0.351 $Y=0.0675 $X2=0.27 $Y2=0.234
cc_72 VSS N_B2_c_95_n 0.00121543f $X=0.351 $Y=0.135 $X2=0.27 $Y2=0.234
cc_73 VSS N_B2_M5_g 2.38303e-19 $X=0.351 $Y=0.0675 $X2=0.27 $Y2=0.2025
cc_74 N_B3_M6_g N_C1_M7_g 0.00333077f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_75 N_B3_c_111_n N_C1_c_124_n 9.33263e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_76 N_B3_c_108_n N_C1_c_119_n 0.00406322f $X=0.405 $Y=0.135 $X2=0.484
+ $Y2=0.0675
cc_77 VSS N_B3_M6_g 3.47199e-19 $X=0.405 $Y=0.0675 $X2=0.484 $Y2=0.2025
cc_78 VSS N_B3_c_108_n 5.30079e-19 $X=0.405 $Y=0.135 $X2=0.484 $Y2=0.2025
cc_79 VSS N_Y_c_131_p 2.4216e-19 $X=0.054 $Y=0.036 $X2=0.469 $Y2=0.2025
cc_80 VSS N_Y_c_132_p 2.72644e-19 $X=0.054 $Y=0.036 $X2=0 $Y2=0

* END of "./OA331x1_ASAP7_75t_L.pex.sp.OA331X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA331x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:49:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA331x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA331x2_ASAP7_75t_L.pex.sp.pex"
* File: OA331x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:49:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA331X2_ASAP7_75T_L%3 2 7 10 13 15 17 20 22 23 26 27 30 34 38 42 47
+ 49 50 51 52 53 57 58 59 60 61 63 66 72 75 84 VSS
c51 84 VSS 0.00202532f $X=0.558 $Y=0.072
c52 83 VSS 0.00163302f $X=0.567 $Y=0.072
c53 77 VSS 6.57651e-19 $X=0.153 $Y=0.195
c54 76 VSS 6.23446e-19 $X=0.144 $Y=0.195
c55 75 VSS 0.00204357f $X=0.162 $Y=0.195
c56 72 VSS 0.00412141f $X=0.567 $Y=0.2
c57 71 VSS 0.00103118f $X=0.567 $Y=0.106
c58 70 VSS 8.11244e-19 $X=0.567 $Y=0.225
c59 68 VSS 6.94247e-19 $X=0.5325 $Y=0.234
c60 67 VSS 2.39163e-19 $X=0.525 $Y=0.234
c61 66 VSS 0.00146362f $X=0.522 $Y=0.234
c62 65 VSS 2.39163e-19 $X=0.504 $Y=0.234
c63 64 VSS 0.00617212f $X=0.501 $Y=0.234
c64 63 VSS 0.00142296f $X=0.468 $Y=0.234
c65 62 VSS 3.71649e-19 $X=0.45 $Y=0.234
c66 61 VSS 0.00311761f $X=0.447 $Y=0.234
c67 60 VSS 0.00146362f $X=0.414 $Y=0.234
c68 59 VSS 0.00340162f $X=0.396 $Y=0.234
c69 58 VSS 0.00146362f $X=0.36 $Y=0.234
c70 57 VSS 0.00256536f $X=0.342 $Y=0.234
c71 53 VSS 8.84964e-19 $X=0.315 $Y=0.234
c72 52 VSS 0.00142296f $X=0.306 $Y=0.234
c73 51 VSS 0.00360252f $X=0.288 $Y=0.234
c74 50 VSS 0.00142296f $X=0.252 $Y=0.234
c75 49 VSS 0.00312977f $X=0.234 $Y=0.234
c76 48 VSS 3.78291e-19 $X=0.202 $Y=0.234
c77 47 VSS 0.00151377f $X=0.198 $Y=0.234
c78 46 VSS 0.00171948f $X=0.18 $Y=0.234
c79 42 VSS 0.00318976f $X=0.171 $Y=0.234
c80 41 VSS 0.00590321f $X=0.558 $Y=0.234
c81 40 VSS 0.00196286f $X=0.162 $Y=0.225
c82 38 VSS 4.04879e-19 $X=0.135 $Y=0.176
c83 34 VSS 6.57355e-19 $X=0.135 $Y=0.135
c84 32 VSS 3.84635e-19 $X=0.135 $Y=0.186
c85 30 VSS 0.00701741f $X=0.538 $Y=0.2025
c86 26 VSS 0.00220219f $X=0.324 $Y=0.2025
c87 22 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c88 20 VSS 0.0013176f $X=0.538 $Y=0.0675
c89 13 VSS 0.00437781f $X=0.135 $Y=0.135
c90 10 VSS 0.0609638f $X=0.135 $Y=0.0675
c91 2 VSS 0.0639847f $X=0.081 $Y=0.0675
r92 84 85 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.072 $X2=0.5625 $Y2=0.072
r93 83 85 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.072 $X2=0.5625 $Y2=0.072
r94 80 84 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.072 $X2=0.558 $Y2=0.072
r95 76 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.195 $X2=0.153 $Y2=0.195
r96 75 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.195 $X2=0.153 $Y2=0.195
r97 73 76 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.195 $X2=0.144 $Y2=0.195
r98 71 72 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.106 $X2=0.567 $Y2=0.2
r99 70 72 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.225 $X2=0.567 $Y2=0.2
r100 69 83 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.567 $Y2=0.072
r101 69 71 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.567 $Y2=0.106
r102 67 68 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.525
+ $Y=0.234 $X2=0.5325 $Y2=0.234
r103 66 67 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.234 $X2=0.525 $Y2=0.234
r104 65 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.522 $Y2=0.234
r105 64 65 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.501
+ $Y=0.234 $X2=0.504 $Y2=0.234
r106 63 64 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.501 $Y2=0.234
r107 62 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r108 61 62 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.234 $X2=0.45 $Y2=0.234
r109 60 61 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.447 $Y2=0.234
r110 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r111 58 59 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.396 $Y2=0.234
r112 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r113 55 68 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.5325 $Y2=0.234
r114 52 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.315 $Y2=0.234
r115 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r116 50 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.288 $Y2=0.234
r117 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r118 48 49 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.234 $X2=0.234 $Y2=0.234
r119 47 48 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.202 $Y2=0.234
r120 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r121 44 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.342 $Y2=0.234
r122 44 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.315 $Y2=0.234
r123 42 46 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.234 $X2=0.18 $Y2=0.234
r124 41 70 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.234 $X2=0.567 $Y2=0.225
r125 41 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.54 $Y2=0.234
r126 40 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.225 $X2=0.171 $Y2=0.234
r127 39 75 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.204 $X2=0.162 $Y2=0.195
r128 39 40 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.204 $X2=0.162 $Y2=0.225
r129 37 38 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.166 $X2=0.135 $Y2=0.176
r130 34 37 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.166
r131 32 73 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.186 $X2=0.135 $Y2=0.195
r132 32 38 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.186 $X2=0.135 $Y2=0.176
r133 30 55 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r134 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.538 $Y2=0.2025
r135 26 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r136 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r137 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r138 20 80 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.072 $X2=0.54
+ $Y2=0.072
r139 17 20 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.538 $Y2=0.0675
r140 13 34 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r141 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r142 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r143 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r144 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r145 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA331X2_ASAP7_75T_L%A3 2 5 7 10 18 VSS
c11 10 VSS 0.00328756f $X=0.189 $Y=0.135
c12 5 VSS 0.00115289f $X=0.189 $Y=0.135
c13 2 VSS 0.0585388f $X=0.189 $Y=0.0675
r14 10 18 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA331X2_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c14 14 VSS 5.30982e-19 $X=0.243 $Y=0.155
c15 10 VSS 4.5987e-19 $X=0.243 $Y=0.135
c16 5 VSS 0.0011122f $X=0.243 $Y=0.135
c17 2 VSS 0.059482f $X=0.243 $Y=0.0675
r18 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.155
r19 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r20 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r21 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OA331X2_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c12 10 VSS 4.82288e-19 $X=0.297 $Y=0.135
c13 5 VSS 0.00111383f $X=0.297 $Y=0.135
c14 2 VSS 0.0608639f $X=0.297 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OA331X2_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.351 $Y=0.135
c14 5 VSS 0.00111336f $X=0.351 $Y=0.135
c15 2 VSS 0.0617786f $X=0.351 $Y=0.0675
r16 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.154
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OA331X2_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.405 $Y=0.135
c14 5 VSS 0.00112198f $X=0.405 $Y=0.135
c15 2 VSS 0.0616432f $X=0.405 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OA331X2_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c11 10 VSS 7.24259e-19 $X=0.459 $Y=0.135
c12 5 VSS 0.00113686f $X=0.459 $Y=0.135
c13 2 VSS 0.0618011f $X=0.459 $Y=0.0675
r14 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OA331X2_ASAP7_75T_L%C1 2 5 7 10 14 VSS
c8 10 VSS 0.00201948f $X=0.513 $Y=0.135
c9 5 VSS 0.00178699f $X=0.513 $Y=0.135
c10 2 VSS 0.0660367f $X=0.513 $Y=0.0675
r11 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.155
r12 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OA331X2_ASAP7_75T_L%Y 1 2 6 7 10 14 21 22 26 VSS
c12 26 VSS 0.00659662f $X=0.108 $Y=0.234
c13 24 VSS 0.00385179f $X=0.063 $Y=0.234
c14 22 VSS 0.0091267f $X=0.108 $Y=0.036
c15 21 VSS 0.00682286f $X=0.108 $Y=0.036
c16 19 VSS 0.00385179f $X=0.063 $Y=0.036
c17 18 VSS 9.92723e-19 $X=0.054 $Y=0.2145
c18 16 VSS 0.00440024f $X=0.054 $Y=0.115
c19 15 VSS 0.00219361f $X=0.054 $Y=0.07
c20 14 VSS 0.00620222f $X=0.057 $Y=0.143
c21 12 VSS 9.44835e-19 $X=0.054 $Y=0.225
c22 10 VSS 0.0101881f $X=0.108 $Y=0.2025
c23 6 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c24 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r25 24 26 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.234 $X2=0.108 $Y2=0.234
r26 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r27 19 21 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.036 $X2=0.108 $Y2=0.036
r28 17 18 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.204 $X2=0.054 $Y2=0.2145
r29 15 16 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.07 $X2=0.054 $Y2=0.115
r30 14 17 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.143 $X2=0.054 $Y2=0.204
r31 14 16 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.143 $X2=0.054 $Y2=0.115
r32 12 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.054 $Y=0.225 $X2=0.063 $Y2=0.234
r33 12 18 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.225 $X2=0.054 $Y2=0.2145
r34 11 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.054 $Y=0.045 $X2=0.063 $Y2=0.036
r35 11 15 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.045 $X2=0.054 $Y2=0.07
r36 10 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r37 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r38 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r39 5 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r40 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r41 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OA331x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA331x2_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C1 Y
* 
* Y	Y
* C1	C1
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_12 N_A3_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_A2_M3_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_12 N_A1_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_13 N_B1_M5_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_12 N_B2_M6_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_13 N_B3_M7_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_3_M8_d N_C1_M8_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 N_Y_M9_d N_3_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M10 N_Y_M10_d N_3_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M11 noxref_14 N_A3_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M12 noxref_15 N_A2_M12_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M13 N_3_M13_d N_A1_M13_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M14 noxref_16 N_B1_M14_g N_3_M14_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M15 noxref_17 N_B2_M15_g noxref_16 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M16 VDD N_B3_M16_g noxref_17 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M17 N_3_M17_d N_C1_M17_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
*
* 
* .include "OA331x2_ASAP7_75t_L.pex.sp.OA331X2_ASAP7_75T_L.pxi"
* BEGIN of "./OA331x2_ASAP7_75t_L.pex.sp.OA331X2_ASAP7_75T_L.pxi"
* File: OA331x2_ASAP7_75t_L.pex.sp.OA331X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:49:56 2017
* 
x_PM_OA331X2_ASAP7_75T_L%3 N_3_M0_g N_3_M9_g N_3_M1_g N_3_c_4_p N_3_M10_g
+ N_3_M8_d N_3_c_45_p N_3_M14_s N_3_M13_d N_3_c_13_p N_3_M17_d N_3_c_23_p
+ N_3_c_5_p N_3_c_9_p N_3_c_36_p N_3_c_3_p N_3_c_39_p N_3_c_8_p N_3_c_38_p
+ N_3_c_12_p N_3_c_41_p N_3_c_42_p N_3_c_15_p N_3_c_43_p N_3_c_18_p N_3_c_44_p
+ N_3_c_20_p N_3_c_22_p N_3_c_25_p N_3_c_11_p N_3_c_40_p VSS
+ PM_OA331X2_ASAP7_75T_L%3
x_PM_OA331X2_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_55_n N_A3_M11_g N_A3_c_56_n A3 VSS
+ PM_OA331X2_ASAP7_75T_L%A3
x_PM_OA331X2_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_69_n N_A2_M12_g N_A2_c_70_n A2 VSS
+ PM_OA331X2_ASAP7_75T_L%A2
x_PM_OA331X2_ASAP7_75T_L%A1 N_A1_M4_g N_A1_c_82_n N_A1_M13_g N_A1_c_78_n A1 VSS
+ PM_OA331X2_ASAP7_75T_L%A1
x_PM_OA331X2_ASAP7_75T_L%B1 N_B1_M5_g N_B1_c_94_n N_B1_M14_g N_B1_c_90_n B1 VSS
+ PM_OA331X2_ASAP7_75T_L%B1
x_PM_OA331X2_ASAP7_75T_L%B2 N_B2_M6_g N_B2_c_106_n N_B2_M15_g N_B2_c_103_n B2
+ VSS PM_OA331X2_ASAP7_75T_L%B2
x_PM_OA331X2_ASAP7_75T_L%B3 N_B3_M7_g N_B3_c_119_n N_B3_M16_g N_B3_c_116_n B3
+ VSS PM_OA331X2_ASAP7_75T_L%B3
x_PM_OA331X2_ASAP7_75T_L%C1 N_C1_M8_g N_C1_c_132_n N_C1_M17_g N_C1_c_127_n C1
+ VSS PM_OA331X2_ASAP7_75T_L%C1
x_PM_OA331X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_M10_d N_Y_M9_d N_Y_c_136_n Y
+ N_Y_c_139_n N_Y_c_141_n N_Y_c_142_n VSS PM_OA331X2_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_A3_M2_g 0.00284417f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_A3_M2_g 2.3886e-19 $X=0.198 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_4 N_3_c_4_p N_A3_c_55_n 9.59383e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_5 N_3_c_5_p N_A3_c_56_n 0.00221266f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_6 N_3_c_3_p N_A3_c_56_n 2.7862e-19 $X=0.198 $Y=0.234 $X2=0.189 $Y2=0.135
cc_7 N_3_M1_g N_A2_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_8 N_3_c_8_p N_A2_M3_g 3.38929e-19 $X=0.252 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_9 N_3_c_9_p A2 2.13942e-19 $X=0.135 $Y=0.176 $X2=0 $Y2=0
cc_10 N_3_c_8_p A2 0.00123064f $X=0.252 $Y=0.234 $X2=0 $Y2=0
cc_11 N_3_c_11_p A2 4.18335e-19 $X=0.162 $Y=0.195 $X2=0 $Y2=0
cc_12 N_3_c_12_p N_A1_M4_g 2.56935e-19 $X=0.306 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_13 N_3_c_13_p N_A1_c_78_n 0.0013295f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_14 N_3_c_12_p N_A1_c_78_n 0.00123064f $X=0.306 $Y=0.234 $X2=0.189 $Y2=0.135
cc_15 N_3_c_15_p N_B1_M5_g 2.64276e-19 $X=0.36 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_16 N_3_c_13_p N_B1_c_90_n 0.0013295f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_17 N_3_c_15_p N_B1_c_90_n 0.00124805f $X=0.36 $Y=0.234 $X2=0.189 $Y2=0.135
cc_18 N_3_c_18_p N_B2_M6_g 3.48613e-19 $X=0.414 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_19 N_3_c_18_p N_B2_c_103_n 0.00124805f $X=0.414 $Y=0.234 $X2=0.189 $Y2=0.135
cc_20 N_3_c_20_p N_B3_M7_g 2.56935e-19 $X=0.468 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_21 N_3_c_20_p N_B3_c_116_n 0.00123064f $X=0.468 $Y=0.234 $X2=0.189 $Y2=0.135
cc_22 N_3_c_22_p N_C1_M8_g 2.64276e-19 $X=0.522 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_23 N_3_c_23_p N_C1_c_127_n 0.00114532f $X=0.538 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_24 N_3_c_22_p N_C1_c_127_n 0.00124805f $X=0.522 $Y=0.234 $X2=0.189 $Y2=0.135
cc_25 N_3_c_25_p N_C1_c_127_n 0.00392202f $X=0.567 $Y=0.2 $X2=0.189 $Y2=0.135
cc_26 N_3_c_4_p N_Y_M1_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_27 N_3_c_4_p N_Y_M10_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_28 N_3_c_4_p N_Y_c_136_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_29 N_3_c_5_p N_Y_c_136_n 0.00141343f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_30 N_3_c_5_p Y 0.00193798f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_31 N_3_M0_g N_Y_c_139_n 4.59284e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_32 N_3_c_4_p N_Y_c_139_n 5.51214e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_33 N_3_c_4_p N_Y_c_141_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_34 N_3_M0_g N_Y_c_142_n 4.59284e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_3_c_4_p N_Y_c_142_n 5.51214e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_36 N_3_c_36_p N_Y_c_142_n 9.43741e-19 $X=0.171 $Y=0.234 $X2=0 $Y2=0
cc_37 VSS N_3_c_13_p 0.00138157f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_38 VSS N_3_c_38_p 2.20596e-19 $X=0.288 $Y=0.234 $X2=0 $Y2=0
cc_39 VSS N_3_c_39_p 2.20596e-19 $X=0.234 $Y=0.234 $X2=0 $Y2=0
cc_40 VSS N_3_c_40_p 2.82518e-19 $X=0.558 $Y=0.072 $X2=0 $Y2=0
cc_41 VSS N_3_c_41_p 2.23188e-19 $X=0.315 $Y=0.234 $X2=0 $Y2=0
cc_42 VSS N_3_c_42_p 2.23188e-19 $X=0.342 $Y=0.234 $X2=0 $Y2=0
cc_43 VSS N_3_c_43_p 2.23188e-19 $X=0.396 $Y=0.234 $X2=0 $Y2=0
cc_44 VSS N_3_c_44_p 2.23188e-19 $X=0.447 $Y=0.234 $X2=0 $Y2=0
cc_45 VSS N_3_c_45_p 3.11523e-19 $X=0.538 $Y=0.0675 $X2=0 $Y2=0
cc_46 VSS N_3_c_45_p 0.00333695f $X=0.538 $Y=0.0675 $X2=0.189 $Y2=0.155
cc_47 VSS N_3_c_40_p 4.47506e-19 $X=0.558 $Y=0.072 $X2=0.189 $Y2=0.155
cc_48 VSS N_3_c_39_p 3.25855e-19 $X=0.234 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_49 VSS N_3_c_38_p 3.56327e-19 $X=0.288 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_50 VSS N_3_c_43_p 3.48201e-19 $X=0.396 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_51 VSS N_3_c_44_p 3.30547e-19 $X=0.447 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_52 N_A3_M2_g N_A2_M3_g 0.00344695f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_53 N_A3_c_55_n N_A2_c_69_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_54 N_A3_c_56_n N_A2_c_70_n 0.00286115f $X=0.189 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_55 N_A3_M2_g N_A1_M4_g 2.66145e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_56 VSS N_A3_c_56_n 8.88545e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_57 N_A2_M3_g N_A1_M4_g 0.00327995f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_58 N_A2_c_69_n N_A1_c_82_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_59 N_A2_c_70_n N_A1_c_78_n 0.00482209f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_60 N_A2_M3_g N_B1_M5_g 2.71887e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_61 VSS N_A2_M3_g 3.57119e-19 $X=0.243 $Y=0.0675 $X2=0.341 $Y2=0.2025
cc_62 VSS N_A2_c_70_n 5.37372e-19 $X=0.243 $Y=0.135 $X2=0.341 $Y2=0.2025
cc_63 N_A1_M4_g N_B1_M5_g 0.0036939f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_64 N_A1_c_82_n N_B1_c_94_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_65 N_A1_c_78_n N_B1_c_90_n 0.00406615f $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_66 N_A1_M4_g N_B2_M6_g 3.06651e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_67 VSS N_A1_c_78_n 0.00159458f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_68 N_B1_M5_g N_B2_M6_g 0.00371573f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_69 N_B1_c_94_n N_B2_c_106_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_70 N_B1_c_90_n N_B2_c_103_n 0.00483372f $X=0.351 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_71 N_B1_M5_g N_B3_M7_g 3.06651e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_72 VSS N_B1_M5_g 3.62029e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_73 VSS N_B1_c_90_n 0.0012322f $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_74 N_B2_M6_g N_B3_M7_g 0.0036939f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_75 N_B2_c_106_n N_B3_c_119_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_76 N_B2_c_103_n N_B3_c_116_n 0.00483372f $X=0.405 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_77 N_B2_M6_g N_C1_M8_g 2.71887e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_78 VSS N_B2_M6_g 2.68514e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_79 VSS N_B2_c_103_n 0.00121543f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_80 VSS N_B2_M6_g 2.38303e-19 $X=0.405 $Y=0.0675 $X2=0.538 $Y2=0.0675
cc_81 N_B3_M7_g N_C1_M8_g 0.00333077f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_82 N_B3_c_119_n N_C1_c_132_n 9.33263e-19 $X=0.459 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_83 N_B3_c_116_n N_C1_c_127_n 0.00406322f $X=0.459 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_84 VSS N_B3_M7_g 3.47199e-19 $X=0.459 $Y=0.0675 $X2=0.538 $Y2=0.0675
cc_85 VSS N_B3_c_116_n 5.30079e-19 $X=0.459 $Y=0.135 $X2=0.538 $Y2=0.0675
cc_86 VSS N_Y_c_139_n 2.80341e-19 $X=0.108 $Y=0.036 $X2=0 $Y2=0

* END of "./OA331x2_ASAP7_75t_L.pex.sp.OA331X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA332x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:50:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA332x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA332x1_ASAP7_75t_L.pex.sp.pex"
* File: OA332x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:50:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA332X1_ASAP7_75T_L%3 2 5 7 9 10 13 14 15 18 19 22 26 30 31 32 38 43
+ 44 45 46 47 51 52 53 54 55 57 59 61 62 68 69 70 74 75 VSS
c55 75 VSS 0.00412141f $X=0.567 $Y=0.2
c56 74 VSS 0.00112176f $X=0.567 $Y=0.106
c57 73 VSS 9.6701e-19 $X=0.567 $Y=0.225
c58 71 VSS 4.93718e-20 $X=0.557 $Y=0.072
c59 70 VSS 4.1269e-19 $X=0.556 $Y=0.072
c60 69 VSS 8.46035e-21 $X=0.522 $Y=0.072
c61 68 VSS 4.70878e-19 $X=0.504 $Y=0.072
c62 63 VSS 0.0019286f $X=0.558 $Y=0.072
c63 62 VSS 0.00146362f $X=0.522 $Y=0.234
c64 61 VSS 0.00296425f $X=0.504 $Y=0.234
c65 60 VSS 3.35992e-19 $X=0.471 $Y=0.234
c66 59 VSS 0.00142296f $X=0.468 $Y=0.234
c67 58 VSS 0.00672869f $X=0.45 $Y=0.234
c68 57 VSS 0.00142296f $X=0.414 $Y=0.234
c69 56 VSS 3.35992e-19 $X=0.396 $Y=0.234
c70 55 VSS 0.00311761f $X=0.393 $Y=0.234
c71 54 VSS 0.00146362f $X=0.36 $Y=0.234
c72 53 VSS 0.00340162f $X=0.342 $Y=0.234
c73 52 VSS 0.00146362f $X=0.306 $Y=0.234
c74 51 VSS 0.00256536f $X=0.288 $Y=0.234
c75 47 VSS 8.84964e-19 $X=0.261 $Y=0.234
c76 46 VSS 0.00142296f $X=0.252 $Y=0.234
c77 45 VSS 0.00360252f $X=0.234 $Y=0.234
c78 44 VSS 0.00142296f $X=0.198 $Y=0.234
c79 43 VSS 0.00331443f $X=0.18 $Y=0.234
c80 42 VSS 1.51923e-19 $X=0.146 $Y=0.234
c81 38 VSS 0.00233672f $X=0.144 $Y=0.234
c82 37 VSS 0.00702647f $X=0.558 $Y=0.234
c83 36 VSS 9.0336e-19 $X=0.135 $Y=0.225
c84 34 VSS 0.00182969f $X=0.11 $Y=0.198
c85 33 VSS 8.41473e-20 $X=0.094 $Y=0.198
c86 32 VSS 4.67384e-20 $X=0.09 $Y=0.198
c87 31 VSS 0.00174552f $X=0.126 $Y=0.198
c88 30 VSS 5.06098e-19 $X=0.081 $Y=0.1765
c89 26 VSS 5.20501e-19 $X=0.081 $Y=0.135
c90 24 VSS 4.85855e-19 $X=0.081 $Y=0.189
c91 22 VSS 0.0038436f $X=0.538 $Y=0.2025
c92 18 VSS 0.00220219f $X=0.27 $Y=0.2025
c93 14 VSS 5.38922e-19 $X=0.287 $Y=0.2025
c94 13 VSS 0.0023085f $X=0.486 $Y=0.0675
c95 9 VSS 5.70099e-19 $X=0.503 $Y=0.0675
c96 5 VSS 0.0017666f $X=0.081 $Y=0.135
c97 2 VSS 0.0645889f $X=0.081 $Y=0.0675
r98 74 75 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.106 $X2=0.567 $Y2=0.2
r99 73 75 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.225 $X2=0.567 $Y2=0.2
r100 72 74 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.567 $Y2=0.106
r101 70 71 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.556
+ $Y=0.072 $X2=0.557 $Y2=0.072
r102 69 70 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.072 $X2=0.556 $Y2=0.072
r103 68 69 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.072 $X2=0.522 $Y2=0.072
r104 65 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.072 $X2=0.504 $Y2=0.072
r105 63 72 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.072 $X2=0.567 $Y2=0.081
r106 63 71 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.072 $X2=0.557 $Y2=0.072
r107 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.522 $Y2=0.234
r108 60 61 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.471
+ $Y=0.234 $X2=0.504 $Y2=0.234
r109 59 60 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.471 $Y2=0.234
r110 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r111 57 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.45 $Y2=0.234
r112 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r113 55 56 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.393
+ $Y=0.234 $X2=0.396 $Y2=0.234
r114 54 55 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.393 $Y2=0.234
r115 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r116 52 53 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.342 $Y2=0.234
r117 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r118 49 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.522 $Y2=0.234
r119 46 47 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.261 $Y2=0.234
r120 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r121 44 45 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.234 $Y2=0.234
r122 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r123 42 43 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.146
+ $Y=0.234 $X2=0.18 $Y2=0.234
r124 40 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.288 $Y2=0.234
r125 40 47 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.261 $Y2=0.234
r126 38 42 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.146 $Y2=0.234
r127 37 73 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.234 $X2=0.567 $Y2=0.225
r128 37 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.54 $Y2=0.234
r129 36 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.225 $X2=0.144 $Y2=0.234
r130 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.207 $X2=0.135 $Y2=0.225
r131 33 34 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.198 $X2=0.11 $Y2=0.198
r132 32 33 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.198 $X2=0.094 $Y2=0.198
r133 31 35 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.126 $Y=0.198 $X2=0.135 $Y2=0.207
r134 31 34 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.198 $X2=0.11 $Y2=0.198
r135 29 30 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.164 $X2=0.081 $Y2=0.1765
r136 26 29 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.164
r137 24 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.189 $X2=0.09 $Y2=0.198
r138 24 30 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.189 $X2=0.081 $Y2=0.1765
r139 22 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r140 19 22 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.538 $Y2=0.2025
r141 18 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r142 15 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r143 14 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r144 13 65 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.072
+ $X2=0.486 $Y2=0.072
r145 10 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.486 $Y2=0.0675
r146 9 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.0675 $X2=0.486 $Y2=0.0675
r147 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r148 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r149 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA332X1_ASAP7_75T_L%A3 2 5 7 10 16 VSS
c10 10 VSS 0.00251553f $X=0.135 $Y=0.135
c11 5 VSS 0.00122791f $X=0.135 $Y=0.135
c12 2 VSS 0.0596346f $X=0.135 $Y=0.0675
r13 10 16 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.155
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OA332X1_ASAP7_75T_L%A2 2 5 7 10 16 VSS
c16 16 VSS 4.40527e-19 $X=0.189 $Y=0.155
c17 10 VSS 0.00192154f $X=0.189 $Y=0.135
c18 5 VSS 0.00110907f $X=0.189 $Y=0.135
c19 2 VSS 0.059482f $X=0.189 $Y=0.0675
r20 10 16 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.155
r21 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA332X1_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c12 10 VSS 4.82288e-19 $X=0.243 $Y=0.135
c13 5 VSS 0.00111383f $X=0.243 $Y=0.135
c14 2 VSS 0.0608471f $X=0.243 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OA332X1_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.297 $Y=0.135
c14 5 VSS 0.00111336f $X=0.297 $Y=0.135
c15 2 VSS 0.0617786f $X=0.297 $Y=0.0675
r16 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.154
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OA332X1_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.351 $Y=0.135
c14 5 VSS 0.00112198f $X=0.351 $Y=0.135
c15 2 VSS 0.0616432f $X=0.351 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OA332X1_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c12 10 VSS 7.27237e-19 $X=0.405 $Y=0.135
c13 5 VSS 0.00111185f $X=0.405 $Y=0.135
c14 2 VSS 0.0615515f $X=0.405 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OA332X1_ASAP7_75T_L%C2 2 5 7 10 14 VSS
c11 10 VSS 0.00167719f $X=0.459 $Y=0.135
c12 5 VSS 0.00113407f $X=0.459 $Y=0.135
c13 2 VSS 0.0618699f $X=0.459 $Y=0.0675
r14 10 14 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.156
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OA332X1_ASAP7_75T_L%C1 2 5 7 10 14 VSS
c11 10 VSS 4.90626e-19 $X=0.513 $Y=0.135
c12 5 VSS 0.00170409f $X=0.513 $Y=0.135
c13 2 VSS 0.0662985f $X=0.513 $Y=0.0675
r14 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OA332X1_ASAP7_75T_L%Y 1 6 9 14 16 21 22 26 VSS
c8 26 VSS 0.0078719f $X=0.054 $Y=0.234
c9 24 VSS 0.00318685f $X=0.027 $Y=0.234
c10 22 VSS 0.00525295f $X=0.054 $Y=0.036
c11 21 VSS 0.00548172f $X=0.054 $Y=0.036
c12 19 VSS 0.00317012f $X=0.027 $Y=0.036
c13 18 VSS 4.26553e-19 $X=0.018 $Y=0.216
c14 16 VSS 0.00230477f $X=0.018 $Y=0.119
c15 15 VSS 0.00107066f $X=0.018 $Y=0.07
c16 14 VSS 0.00393433f $X=0.0195 $Y=0.1395
c17 12 VSS 4.02856e-19 $X=0.018 $Y=0.225
c18 9 VSS 0.00568786f $X=0.056 $Y=0.2025
c19 6 VSS 2.55988e-19 $X=0.071 $Y=0.2025
c20 1 VSS 3.02808e-19 $X=0.071 $Y=0.0675
r21 24 26 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.054 $Y2=0.234
r22 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r23 19 21 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.054 $Y2=0.036
r24 17 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.207 $X2=0.018 $Y2=0.216
r25 15 16 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.119
r26 14 17 4.58333 $w=1.8e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.207
r27 14 16 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.119
r28 12 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r29 12 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.216
r30 11 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r31 11 15 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r32 9 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r33 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
r34 4 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r35 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./OA332x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA332x1_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 VSS N_3_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 noxref_13 N_A3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_A2_M2_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_13 N_A1_M3_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_14 N_B1_M4_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_13 N_B2_M5_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_14 N_B3_M6_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_3_M7_d N_C2_M7_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 noxref_14 N_C1_M8_g N_3_M8_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 VDD N_3_M9_g N_Y_M9_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M10 noxref_15 N_A3_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M11 noxref_16 N_A2_M11_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.179 $Y=0.162
M12 N_3_M12_d N_A1_M12_g noxref_16 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M13 noxref_17 N_B1_M13_g N_3_M13_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M14 noxref_18 N_B2_M14_g noxref_17 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M15 VDD N_B3_M15_g noxref_18 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M16 noxref_19 N_C2_M16_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M17 N_3_M17_d N_C1_M17_g noxref_19 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
*
* 
* .include "OA332x1_ASAP7_75t_L.pex.sp.OA332X1_ASAP7_75T_L.pxi"
* BEGIN of "./OA332x1_ASAP7_75t_L.pex.sp.OA332X1_ASAP7_75T_L.pxi"
* File: OA332x1_ASAP7_75t_L.pex.sp.OA332X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:50:18 2017
* 
x_PM_OA332X1_ASAP7_75T_L%3 N_3_M0_g N_3_c_2_p N_3_M9_g N_3_M8_s N_3_M7_d
+ N_3_c_42_p N_3_M13_s N_3_M12_d N_3_c_11_p N_3_M17_d N_3_c_24_p N_3_c_3_p
+ N_3_c_7_p N_3_c_4_p N_3_c_31_p N_3_c_32_p N_3_c_35_p N_3_c_6_p N_3_c_34_p
+ N_3_c_10_p N_3_c_37_p N_3_c_38_p N_3_c_13_p N_3_c_39_p N_3_c_16_p N_3_c_40_p
+ N_3_c_18_p N_3_c_20_p N_3_c_55_p N_3_c_22_p N_3_c_36_p N_3_c_23_p N_3_c_41_p
+ N_3_c_48_p N_3_c_27_p VSS PM_OA332X1_ASAP7_75T_L%3
x_PM_OA332X1_ASAP7_75T_L%A3 N_A3_M1_g N_A3_c_57_n N_A3_M10_g N_A3_c_58_n A3 VSS
+ PM_OA332X1_ASAP7_75T_L%A3
x_PM_OA332X1_ASAP7_75T_L%A2 N_A2_M2_g N_A2_c_72_n N_A2_M11_g N_A2_c_73_n A2 VSS
+ PM_OA332X1_ASAP7_75T_L%A2
x_PM_OA332X1_ASAP7_75T_L%A1 N_A1_M3_g N_A1_c_87_n N_A1_M12_g N_A1_c_83_n A1 VSS
+ PM_OA332X1_ASAP7_75T_L%A1
x_PM_OA332X1_ASAP7_75T_L%B1 N_B1_M4_g N_B1_c_99_n N_B1_M13_g N_B1_c_95_n B1 VSS
+ PM_OA332X1_ASAP7_75T_L%B1
x_PM_OA332X1_ASAP7_75T_L%B2 N_B2_M5_g N_B2_c_111_n N_B2_M14_g N_B2_c_108_n B2
+ VSS PM_OA332X1_ASAP7_75T_L%B2
x_PM_OA332X1_ASAP7_75T_L%B3 N_B3_M6_g N_B3_c_124_n N_B3_M15_g N_B3_c_121_n B3
+ VSS PM_OA332X1_ASAP7_75T_L%B3
x_PM_OA332X1_ASAP7_75T_L%C2 N_C2_M7_g N_C2_c_136_n N_C2_M16_g N_C2_c_133_n C2
+ VSS PM_OA332X1_ASAP7_75T_L%C2
x_PM_OA332X1_ASAP7_75T_L%C1 N_C1_M8_g N_C1_c_151_n N_C1_M17_g N_C1_c_145_n C1
+ VSS PM_OA332X1_ASAP7_75T_L%C1
x_PM_OA332X1_ASAP7_75T_L%Y N_Y_M0_s N_Y_M9_s N_Y_c_154_n Y N_Y_c_159_n
+ N_Y_c_161_p N_Y_c_160_p N_Y_c_156_n VSS PM_OA332X1_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M1_g 0.00286002f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_3_c_2_p N_A3_c_57_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_3_c_3_p N_A3_c_58_n 0.00196469f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_3_c_4_p N_A3_c_58_n 0.00133324f $X=0.126 $Y=0.198 $X2=0.135 $Y2=0.135
cc_5 N_3_M0_g N_A2_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 N_3_c_6_p N_A2_M2_g 3.38929e-19 $X=0.198 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_7 N_3_c_7_p A2 2.69033e-19 $X=0.081 $Y=0.1765 $X2=0.135 $Y2=0.155
cc_8 N_3_c_4_p A2 7.10035e-19 $X=0.126 $Y=0.198 $X2=0.135 $Y2=0.155
cc_9 N_3_c_6_p A2 0.00123604f $X=0.198 $Y=0.234 $X2=0.135 $Y2=0.155
cc_10 N_3_c_10_p N_A1_M3_g 2.56935e-19 $X=0.252 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_11 N_3_c_11_p N_A1_c_83_n 0.0013295f $X=0.27 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_12 N_3_c_10_p N_A1_c_83_n 0.00123064f $X=0.252 $Y=0.234 $X2=0.135 $Y2=0.135
cc_13 N_3_c_13_p N_B1_M4_g 2.64276e-19 $X=0.306 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_14 N_3_c_11_p N_B1_c_95_n 0.0013295f $X=0.27 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_15 N_3_c_13_p N_B1_c_95_n 0.00124805f $X=0.306 $Y=0.234 $X2=0.135 $Y2=0.135
cc_16 N_3_c_16_p N_B2_M5_g 3.48613e-19 $X=0.36 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_17 N_3_c_16_p N_B2_c_108_n 0.00124805f $X=0.36 $Y=0.234 $X2=0.135 $Y2=0.135
cc_18 N_3_c_18_p N_B3_M6_g 2.56935e-19 $X=0.414 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_19 N_3_c_18_p N_B3_c_121_n 0.00123064f $X=0.414 $Y=0.234 $X2=0.135 $Y2=0.135
cc_20 N_3_c_20_p N_C2_M7_g 2.56935e-19 $X=0.468 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_21 N_3_c_20_p N_C2_c_133_n 0.00123064f $X=0.468 $Y=0.234 $X2=0.135 $Y2=0.135
cc_22 N_3_c_22_p N_C1_M8_g 2.64276e-19 $X=0.522 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_23 N_3_c_23_p N_C1_M8_g 2.76185e-19 $X=0.522 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_24 N_3_c_24_p N_C1_c_145_n 0.0013399f $X=0.538 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_25 N_3_c_22_p N_C1_c_145_n 0.00124805f $X=0.522 $Y=0.234 $X2=0.135 $Y2=0.135
cc_26 N_3_c_23_p N_C1_c_145_n 0.0012322f $X=0.522 $Y=0.072 $X2=0.135 $Y2=0.135
cc_27 N_3_c_27_p N_C1_c_145_n 0.00392202f $X=0.567 $Y=0.2 $X2=0.135 $Y2=0.135
cc_28 N_3_c_3_p N_Y_c_154_n 0.00143087f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_29 N_3_c_3_p Y 0.00278222f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_30 N_3_M0_g N_Y_c_156_n 2.34993e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_3_c_31_p N_Y_c_156_n 0.00197676f $X=0.09 $Y=0.198 $X2=0 $Y2=0
cc_32 N_3_c_32_p N_Y_c_156_n 7.93849e-19 $X=0.144 $Y=0.234 $X2=0 $Y2=0
cc_33 VSS N_3_c_11_p 0.00138157f $X=0.27 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_34 VSS N_3_c_34_p 2.30767e-19 $X=0.234 $Y=0.234 $X2=0.135 $Y2=0.155
cc_35 VSS N_3_c_35_p 2.30767e-19 $X=0.18 $Y=0.234 $X2=0 $Y2=0
cc_36 VSS N_3_c_36_p 2.9669e-19 $X=0.504 $Y=0.072 $X2=0 $Y2=0
cc_37 VSS N_3_c_37_p 2.23188e-19 $X=0.261 $Y=0.234 $X2=0 $Y2=0
cc_38 VSS N_3_c_38_p 2.23188e-19 $X=0.288 $Y=0.234 $X2=0 $Y2=0
cc_39 VSS N_3_c_39_p 2.23188e-19 $X=0.342 $Y=0.234 $X2=0 $Y2=0
cc_40 VSS N_3_c_40_p 2.23188e-19 $X=0.393 $Y=0.234 $X2=0 $Y2=0
cc_41 VSS N_3_c_41_p 2.47657e-19 $X=0.556 $Y=0.072 $X2=0 $Y2=0
cc_42 VSS N_3_c_42_p 0.00333582f $X=0.486 $Y=0.0675 $X2=0 $Y2=0
cc_43 VSS N_3_c_36_p 4.54465e-19 $X=0.504 $Y=0.072 $X2=0 $Y2=0
cc_44 VSS N_3_c_23_p 0.00365373f $X=0.522 $Y=0.072 $X2=0 $Y2=0
cc_45 VSS N_3_c_42_p 0.00371671f $X=0.486 $Y=0.0675 $X2=0 $Y2=0
cc_46 VSS N_3_c_24_p 0.00138157f $X=0.538 $Y=0.2025 $X2=0 $Y2=0
cc_47 VSS N_3_c_41_p 0.00260156f $X=0.556 $Y=0.072 $X2=0 $Y2=0
cc_48 VSS N_3_c_48_p 3.97918e-19 $X=0.567 $Y=0.106 $X2=0 $Y2=0
cc_49 VSS N_3_c_42_p 0.00250965f $X=0.486 $Y=0.0675 $X2=0 $Y2=0
cc_50 VSS N_3_c_36_p 0.00365373f $X=0.504 $Y=0.072 $X2=0 $Y2=0
cc_51 VSS N_3_c_35_p 3.56327e-19 $X=0.18 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_52 VSS N_3_c_34_p 3.56327e-19 $X=0.234 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_53 VSS N_3_c_39_p 3.48201e-19 $X=0.342 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_54 VSS N_3_c_40_p 3.30547e-19 $X=0.393 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_55 VSS N_3_c_55_p 3.30547e-19 $X=0.504 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_56 N_A3_M1_g N_A2_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_57 N_A3_c_57_n N_A2_c_72_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_58 N_A3_c_58_n N_A2_c_73_n 0.00392079f $X=0.135 $Y=0.135 $X2=0.469 $Y2=0.0675
cc_59 N_A3_M1_g N_A1_M3_g 2.66145e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_60 N_A3_c_58_n N_Y_c_159_n 4.54513e-19 $X=0.135 $Y=0.135 $X2=0.27 $Y2=0.2025
cc_61 VSS N_A3_c_58_n 0.00114532f $X=0.135 $Y=0.135 $X2=0.523 $Y2=0.2025
cc_62 N_A2_M2_g N_A1_M3_g 0.00327995f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_63 N_A2_c_72_n N_A1_c_87_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_64 N_A2_c_73_n N_A1_c_83_n 0.00464977f $X=0.189 $Y=0.135 $X2=0.469 $Y2=0.0675
cc_65 N_A2_M2_g N_B1_M4_g 2.71887e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_66 VSS N_A2_c_73_n 0.0011319f $X=0.189 $Y=0.135 $X2=0.523 $Y2=0.2025
cc_67 VSS N_A2_M2_g 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0.538 $Y2=0.2025
cc_68 VSS N_A2_c_73_n 0.00125352f $X=0.189 $Y=0.135 $X2=0.538 $Y2=0.2025
cc_69 VSS N_A2_c_73_n 4.64812e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_70 N_A1_M3_g N_B1_M4_g 0.0036939f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_71 N_A1_c_87_n N_B1_c_99_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_72 N_A1_c_83_n N_B1_c_95_n 0.00406615f $X=0.243 $Y=0.135 $X2=0.469 $Y2=0.0675
cc_73 N_A1_M3_g N_B2_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_74 VSS N_A1_c_83_n 0.00159458f $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_75 N_B1_M4_g N_B2_M5_g 0.00371573f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_76 N_B1_c_99_n N_B2_c_111_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_77 N_B1_c_95_n N_B2_c_108_n 0.00483372f $X=0.297 $Y=0.135 $X2=0.469
+ $Y2=0.0675
cc_78 N_B1_M4_g N_B3_M6_g 3.06651e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_79 VSS N_B1_M4_g 3.62029e-19 $X=0.297 $Y=0.0675 $X2=0.094 $Y2=0.198
cc_80 VSS N_B1_c_95_n 0.0012322f $X=0.297 $Y=0.135 $X2=0.094 $Y2=0.198
cc_81 N_B2_M5_g N_B3_M6_g 0.0036939f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_82 N_B2_c_111_n N_B3_c_124_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_83 N_B2_c_108_n N_B3_c_121_n 0.00483372f $X=0.351 $Y=0.135 $X2=0.469
+ $Y2=0.0675
cc_84 N_B2_M5_g N_C2_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_85 VSS N_B2_M5_g 2.68514e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.225
cc_86 VSS N_B2_c_108_n 0.00121543f $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.225
cc_87 VSS N_B2_M5_g 2.38303e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_88 N_B3_M6_g N_C2_M7_g 0.00333077f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_89 N_B3_c_124_n N_C2_c_136_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_90 N_B3_c_121_n N_C2_c_133_n 0.00406615f $X=0.405 $Y=0.135 $X2=0.469
+ $Y2=0.0675
cc_91 N_B3_M6_g N_C1_M8_g 2.71887e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_92 VSS N_B3_M6_g 3.47199e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_93 VSS N_B3_c_121_n 5.30079e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_94 N_C2_M7_g N_C1_M8_g 0.0036939f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_95 N_C2_c_136_n N_C1_c_151_n 9.33263e-19 $X=0.459 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_96 N_C2_c_133_n N_C1_c_145_n 0.00477924f $X=0.459 $Y=0.135 $X2=0.469
+ $Y2=0.0675
cc_97 VSS N_C2_M7_g 3.57119e-19 $X=0.459 $Y=0.0675 $X2=0.126 $Y2=0.198
cc_98 VSS N_C2_c_133_n 5.37372e-19 $X=0.459 $Y=0.135 $X2=0.126 $Y2=0.198
cc_99 VSS N_C1_M8_g 2.15135e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_100 VSS N_Y_c_160_p 2.2337e-19 $X=0.054 $Y=0.036 $X2=0.523 $Y2=0.2025
cc_101 VSS N_Y_c_161_p 2.82839e-19 $X=0.054 $Y=0.036 $X2=0 $Y2=0

* END of "./OA332x1_ASAP7_75t_L.pex.sp.OA332X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA332x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:50:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA332x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA332x2_ASAP7_75t_L.pex.sp.pex"
* File: OA332x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:50:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA332X2_ASAP7_75T_L%3 2 7 10 13 15 17 18 21 22 23 26 27 30 34 38 39
+ 40 46 51 52 53 54 55 59 60 61 62 63 65 67 69 70 76 77 78 82 83 VSS
c65 83 VSS 0.00412141f $X=0.621 $Y=0.2
c66 82 VSS 0.00112176f $X=0.621 $Y=0.106
c67 81 VSS 9.6701e-19 $X=0.621 $Y=0.225
c68 79 VSS 4.93718e-20 $X=0.611 $Y=0.072
c69 78 VSS 4.1269e-19 $X=0.61 $Y=0.072
c70 77 VSS 8.46035e-21 $X=0.576 $Y=0.072
c71 76 VSS 4.70878e-19 $X=0.558 $Y=0.072
c72 71 VSS 0.0019286f $X=0.612 $Y=0.072
c73 70 VSS 0.00146362f $X=0.576 $Y=0.234
c74 69 VSS 0.00296425f $X=0.558 $Y=0.234
c75 68 VSS 3.35992e-19 $X=0.525 $Y=0.234
c76 67 VSS 0.00142296f $X=0.522 $Y=0.234
c77 66 VSS 0.00672869f $X=0.504 $Y=0.234
c78 65 VSS 0.00142296f $X=0.468 $Y=0.234
c79 64 VSS 3.35992e-19 $X=0.45 $Y=0.234
c80 63 VSS 0.00311761f $X=0.447 $Y=0.234
c81 62 VSS 0.00146362f $X=0.414 $Y=0.234
c82 61 VSS 0.00340162f $X=0.396 $Y=0.234
c83 60 VSS 0.00146362f $X=0.36 $Y=0.234
c84 59 VSS 0.00256536f $X=0.342 $Y=0.234
c85 55 VSS 8.84964e-19 $X=0.315 $Y=0.234
c86 54 VSS 0.00142296f $X=0.306 $Y=0.234
c87 53 VSS 0.00360252f $X=0.288 $Y=0.234
c88 52 VSS 0.00142296f $X=0.252 $Y=0.234
c89 51 VSS 0.00331443f $X=0.234 $Y=0.234
c90 50 VSS 1.51923e-19 $X=0.2 $Y=0.234
c91 46 VSS 0.00233672f $X=0.198 $Y=0.234
c92 45 VSS 0.00702647f $X=0.612 $Y=0.234
c93 44 VSS 9.0336e-19 $X=0.189 $Y=0.225
c94 42 VSS 0.00182969f $X=0.164 $Y=0.198
c95 41 VSS 8.41473e-20 $X=0.148 $Y=0.198
c96 40 VSS 4.67384e-20 $X=0.144 $Y=0.198
c97 39 VSS 0.00174552f $X=0.18 $Y=0.198
c98 38 VSS 5.06098e-19 $X=0.135 $Y=0.1765
c99 34 VSS 5.77929e-19 $X=0.135 $Y=0.135
c100 32 VSS 4.85855e-19 $X=0.135 $Y=0.189
c101 30 VSS 0.0038436f $X=0.592 $Y=0.2025
c102 26 VSS 0.00220219f $X=0.324 $Y=0.2025
c103 22 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c104 21 VSS 0.0023085f $X=0.54 $Y=0.0675
c105 17 VSS 5.70099e-19 $X=0.557 $Y=0.0675
c106 13 VSS 0.00396933f $X=0.135 $Y=0.135
c107 10 VSS 0.0608916f $X=0.135 $Y=0.0675
c108 2 VSS 0.0615048f $X=0.081 $Y=0.0675
r109 82 83 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.106 $X2=0.621 $Y2=0.2
r110 81 83 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.2
r111 80 82 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.081 $X2=0.621 $Y2=0.106
r112 78 79 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.61
+ $Y=0.072 $X2=0.611 $Y2=0.072
r113 77 78 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.072 $X2=0.61 $Y2=0.072
r114 76 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.072 $X2=0.576 $Y2=0.072
r115 73 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.072 $X2=0.558 $Y2=0.072
r116 71 80 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.072 $X2=0.621 $Y2=0.081
r117 71 79 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.072 $X2=0.611 $Y2=0.072
r118 69 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.576 $Y2=0.234
r119 68 69 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.525
+ $Y=0.234 $X2=0.558 $Y2=0.234
r120 67 68 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.234 $X2=0.525 $Y2=0.234
r121 66 67 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.522 $Y2=0.234
r122 65 66 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.504 $Y2=0.234
r123 64 65 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r124 63 64 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.234 $X2=0.45 $Y2=0.234
r125 62 63 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.447 $Y2=0.234
r126 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r127 60 61 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.396 $Y2=0.234
r128 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r129 57 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.576 $Y2=0.234
r130 54 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.315 $Y2=0.234
r131 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r132 52 53 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.288 $Y2=0.234
r133 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r134 50 51 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.2
+ $Y=0.234 $X2=0.234 $Y2=0.234
r135 48 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.342 $Y2=0.234
r136 48 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.315 $Y2=0.234
r137 46 50 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.2 $Y2=0.234
r138 45 81 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r139 45 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r140 44 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.225 $X2=0.198 $Y2=0.234
r141 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.207 $X2=0.189 $Y2=0.225
r142 41 42 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.198 $X2=0.164 $Y2=0.198
r143 40 41 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.198 $X2=0.148 $Y2=0.198
r144 39 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.198 $X2=0.189 $Y2=0.207
r145 39 42 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.198 $X2=0.164 $Y2=0.198
r146 37 38 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.164 $X2=0.135 $Y2=0.1765
r147 34 37 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.164
r148 32 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.189 $X2=0.144 $Y2=0.198
r149 32 38 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.135 $Y2=0.1765
r150 30 57 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r151 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2025 $X2=0.592 $Y2=0.2025
r152 26 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r153 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r154 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r155 21 73 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.072 $X2=0.54
+ $Y2=0.072
r156 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r157 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r158 13 34 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r159 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r160 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r161 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r162 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r163 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA332X2_ASAP7_75T_L%A3 2 5 7 10 16 VSS
c11 10 VSS 0.00277936f $X=0.189 $Y=0.135
c12 5 VSS 0.0011078f $X=0.189 $Y=0.135
c13 2 VSS 0.0588833f $X=0.189 $Y=0.0675
r14 10 16 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA332X2_ASAP7_75T_L%A2 2 5 7 10 16 VSS
c16 16 VSS 4.40527e-19 $X=0.243 $Y=0.155
c17 10 VSS 0.00192154f $X=0.243 $Y=0.135
c18 5 VSS 0.00111216f $X=0.243 $Y=0.135
c19 2 VSS 0.059482f $X=0.243 $Y=0.0675
r20 10 16 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.155
r21 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OA332X2_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c12 10 VSS 4.82288e-19 $X=0.297 $Y=0.135
c13 5 VSS 0.00111383f $X=0.297 $Y=0.135
c14 2 VSS 0.0608471f $X=0.297 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OA332X2_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.351 $Y=0.135
c14 5 VSS 0.00111336f $X=0.351 $Y=0.135
c15 2 VSS 0.0617786f $X=0.351 $Y=0.0675
r16 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.154
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OA332X2_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.405 $Y=0.135
c14 5 VSS 0.00112198f $X=0.405 $Y=0.135
c15 2 VSS 0.0616432f $X=0.405 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OA332X2_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c12 10 VSS 7.27237e-19 $X=0.459 $Y=0.135
c13 5 VSS 0.00111185f $X=0.459 $Y=0.135
c14 2 VSS 0.0615515f $X=0.459 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OA332X2_ASAP7_75T_L%C2 2 5 7 10 14 VSS
c11 10 VSS 0.00167719f $X=0.513 $Y=0.135
c12 5 VSS 0.00113407f $X=0.513 $Y=0.135
c13 2 VSS 0.0618699f $X=0.513 $Y=0.0675
r14 10 14 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.156
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OA332X2_ASAP7_75T_L%C1 2 5 7 10 14 VSS
c11 10 VSS 4.90626e-19 $X=0.567 $Y=0.135
c12 5 VSS 0.00170409f $X=0.567 $Y=0.135
c13 2 VSS 0.0662985f $X=0.567 $Y=0.0675
r14 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
.ends

.subckt PM_OA332X2_ASAP7_75T_L%Y 1 2 6 7 10 14 16 21 22 26 VSS
c17 26 VSS 0.0154624f $X=0.108 $Y=0.234
c18 24 VSS 0.0032101f $X=0.027 $Y=0.234
c19 22 VSS 0.00902033f $X=0.108 $Y=0.036
c20 21 VSS 0.0131561f $X=0.108 $Y=0.036
c21 19 VSS 0.00320021f $X=0.027 $Y=0.036
c22 18 VSS 4.26553e-19 $X=0.018 $Y=0.216
c23 16 VSS 0.00278197f $X=0.018 $Y=0.119
c24 15 VSS 0.00126561f $X=0.018 $Y=0.07
c25 14 VSS 0.00449127f $X=0.0195 $Y=0.1395
c26 12 VSS 4.02856e-19 $X=0.018 $Y=0.225
c27 10 VSS 0.0102944f $X=0.108 $Y=0.2025
c28 6 VSS 5.25448e-19 $X=0.125 $Y=0.2025
c29 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r30 24 26 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.108 $Y2=0.234
r31 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r32 19 21 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.108 $Y2=0.036
r33 17 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.207 $X2=0.018 $Y2=0.216
r34 15 16 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.119
r35 14 17 4.58333 $w=1.8e-08 $l=6.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.207
r36 14 16 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.1395 $X2=0.018 $Y2=0.119
r37 12 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r38 12 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.216
r39 11 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r40 11 15 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r41 10 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r42 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r43 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r44 5 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r45 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r46 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OA332x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA332x2_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_13 N_A3_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_A2_M3_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_13 N_A1_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_14 N_B1_M5_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_13 N_B2_M6_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_14 N_B3_M7_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_3_M8_d N_C2_M8_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 noxref_14 N_C1_M9_g N_3_M9_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M10 N_Y_M10_d N_3_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M11 N_Y_M11_d N_3_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M12 noxref_15 N_A3_M12_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M13 noxref_16 N_A2_M13_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M14 N_3_M14_d N_A1_M14_g noxref_16 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M15 noxref_17 N_B1_M15_g N_3_M15_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M16 noxref_18 N_B2_M16_g noxref_17 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M17 VDD N_B3_M17_g noxref_18 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M18 noxref_19 N_C2_M18_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M19 N_3_M19_d N_C1_M19_g noxref_19 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
*
* 
* .include "OA332x2_ASAP7_75t_L.pex.sp.OA332X2_ASAP7_75T_L.pxi"
* BEGIN of "./OA332x2_ASAP7_75t_L.pex.sp.OA332X2_ASAP7_75T_L.pxi"
* File: OA332x2_ASAP7_75t_L.pex.sp.OA332X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:50:41 2017
* 
x_PM_OA332X2_ASAP7_75T_L%3 N_3_M0_g N_3_M10_g N_3_M1_g N_3_c_3_p N_3_M11_g
+ N_3_M9_s N_3_M8_d N_3_c_52_p N_3_M15_s N_3_M14_d N_3_c_12_p N_3_M19_d
+ N_3_c_25_p N_3_c_4_p N_3_c_8_p N_3_c_5_p N_3_c_41_p N_3_c_42_p N_3_c_45_p
+ N_3_c_7_p N_3_c_44_p N_3_c_11_p N_3_c_47_p N_3_c_48_p N_3_c_14_p N_3_c_49_p
+ N_3_c_17_p N_3_c_50_p N_3_c_19_p N_3_c_21_p N_3_c_65_p N_3_c_23_p N_3_c_46_p
+ N_3_c_24_p N_3_c_51_p N_3_c_58_p N_3_c_28_p VSS PM_OA332X2_ASAP7_75T_L%3
x_PM_OA332X2_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_68_n N_A3_M12_g N_A3_c_69_n A3 VSS
+ PM_OA332X2_ASAP7_75T_L%A3
x_PM_OA332X2_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_83_n N_A2_M13_g N_A2_c_84_n A2 VSS
+ PM_OA332X2_ASAP7_75T_L%A2
x_PM_OA332X2_ASAP7_75T_L%A1 N_A1_M4_g N_A1_c_98_n N_A1_M14_g N_A1_c_94_n A1 VSS
+ PM_OA332X2_ASAP7_75T_L%A1
x_PM_OA332X2_ASAP7_75T_L%B1 N_B1_M5_g N_B1_c_110_n N_B1_M15_g N_B1_c_106_n B1
+ VSS PM_OA332X2_ASAP7_75T_L%B1
x_PM_OA332X2_ASAP7_75T_L%B2 N_B2_M6_g N_B2_c_122_n N_B2_M16_g N_B2_c_119_n B2
+ VSS PM_OA332X2_ASAP7_75T_L%B2
x_PM_OA332X2_ASAP7_75T_L%B3 N_B3_M7_g N_B3_c_135_n N_B3_M17_g N_B3_c_132_n B3
+ VSS PM_OA332X2_ASAP7_75T_L%B3
x_PM_OA332X2_ASAP7_75T_L%C2 N_C2_M8_g N_C2_c_147_n N_C2_M18_g N_C2_c_144_n C2
+ VSS PM_OA332X2_ASAP7_75T_L%C2
x_PM_OA332X2_ASAP7_75T_L%C1 N_C1_M9_g N_C1_c_162_n N_C1_M19_g N_C1_c_156_n C1
+ VSS PM_OA332X2_ASAP7_75T_L%C1
x_PM_OA332X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_M11_d N_Y_M10_d N_Y_c_167_n Y
+ N_Y_c_179_n N_Y_c_171_n N_Y_c_173_n N_Y_c_174_n VSS PM_OA332X2_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A3_M2_g 2.13359e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_A3_M2_g 0.00286002f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_A3_c_68_n 9.59209e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_4 N_3_c_4_p N_A3_c_69_n 0.00196691f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_5 N_3_c_5_p N_A3_c_69_n 0.00133324f $X=0.18 $Y=0.198 $X2=0.189 $Y2=0.135
cc_6 N_3_M1_g N_A2_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_7 N_3_c_7_p N_A2_M3_g 3.38929e-19 $X=0.252 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_8 N_3_c_8_p A2 2.69033e-19 $X=0.135 $Y=0.1765 $X2=0.189 $Y2=0.155
cc_9 N_3_c_5_p A2 7.10035e-19 $X=0.18 $Y=0.198 $X2=0.189 $Y2=0.155
cc_10 N_3_c_7_p A2 0.00123604f $X=0.252 $Y=0.234 $X2=0.189 $Y2=0.155
cc_11 N_3_c_11_p N_A1_M4_g 2.56935e-19 $X=0.306 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_12 N_3_c_12_p N_A1_c_94_n 0.0013295f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_13 N_3_c_11_p N_A1_c_94_n 0.00123064f $X=0.306 $Y=0.234 $X2=0.189 $Y2=0.135
cc_14 N_3_c_14_p N_B1_M5_g 2.64276e-19 $X=0.36 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_15 N_3_c_12_p N_B1_c_106_n 0.0013295f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_16 N_3_c_14_p N_B1_c_106_n 0.00124805f $X=0.36 $Y=0.234 $X2=0.189 $Y2=0.135
cc_17 N_3_c_17_p N_B2_M6_g 3.48613e-19 $X=0.414 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_18 N_3_c_17_p N_B2_c_119_n 0.00124805f $X=0.414 $Y=0.234 $X2=0.189 $Y2=0.135
cc_19 N_3_c_19_p N_B3_M7_g 2.56935e-19 $X=0.468 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_20 N_3_c_19_p N_B3_c_132_n 0.00123064f $X=0.468 $Y=0.234 $X2=0.189 $Y2=0.135
cc_21 N_3_c_21_p N_C2_M8_g 2.56935e-19 $X=0.522 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_22 N_3_c_21_p N_C2_c_144_n 0.00123064f $X=0.522 $Y=0.234 $X2=0.189 $Y2=0.135
cc_23 N_3_c_23_p N_C1_M9_g 2.64276e-19 $X=0.576 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_24 N_3_c_24_p N_C1_M9_g 2.76185e-19 $X=0.576 $Y=0.072 $X2=0.189 $Y2=0.0675
cc_25 N_3_c_25_p N_C1_c_156_n 0.0013399f $X=0.592 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_26 N_3_c_23_p N_C1_c_156_n 0.00124805f $X=0.576 $Y=0.234 $X2=0.189 $Y2=0.135
cc_27 N_3_c_24_p N_C1_c_156_n 0.0012322f $X=0.576 $Y=0.072 $X2=0.189 $Y2=0.135
cc_28 N_3_c_28_p N_C1_c_156_n 0.00392202f $X=0.621 $Y=0.2 $X2=0.189 $Y2=0.135
cc_29 N_3_c_3_p N_Y_M1_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_30 N_3_c_3_p N_Y_M11_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_31 N_3_c_3_p N_Y_c_167_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_32 N_3_c_4_p N_Y_c_167_n 0.00156987f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_33 N_3_c_3_p Y 3.36333e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_34 N_3_c_4_p Y 9.49917e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_35 N_3_M0_g N_Y_c_171_n 4.59284e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_3_c_3_p N_Y_c_171_n 5.35059e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_37 N_3_c_3_p N_Y_c_173_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_38 N_3_M0_g N_Y_c_174_n 4.59284e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_3_M1_g N_Y_c_174_n 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_40 N_3_c_3_p N_Y_c_174_n 5.94649e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_41 N_3_c_41_p N_Y_c_174_n 0.00197676f $X=0.144 $Y=0.198 $X2=0 $Y2=0
cc_42 N_3_c_42_p N_Y_c_174_n 8.21768e-19 $X=0.198 $Y=0.234 $X2=0 $Y2=0
cc_43 VSS N_3_c_12_p 0.00138157f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_44 VSS N_3_c_44_p 2.30767e-19 $X=0.288 $Y=0.234 $X2=0.189 $Y2=0.155
cc_45 VSS N_3_c_45_p 2.30767e-19 $X=0.234 $Y=0.234 $X2=0 $Y2=0
cc_46 VSS N_3_c_46_p 2.9669e-19 $X=0.558 $Y=0.072 $X2=0 $Y2=0
cc_47 VSS N_3_c_47_p 2.23188e-19 $X=0.315 $Y=0.234 $X2=0 $Y2=0
cc_48 VSS N_3_c_48_p 2.23188e-19 $X=0.342 $Y=0.234 $X2=0 $Y2=0
cc_49 VSS N_3_c_49_p 2.23188e-19 $X=0.396 $Y=0.234 $X2=0 $Y2=0
cc_50 VSS N_3_c_50_p 2.23188e-19 $X=0.447 $Y=0.234 $X2=0 $Y2=0
cc_51 VSS N_3_c_51_p 2.47657e-19 $X=0.61 $Y=0.072 $X2=0 $Y2=0
cc_52 VSS N_3_c_52_p 0.00333582f $X=0.54 $Y=0.0675 $X2=0 $Y2=0
cc_53 VSS N_3_c_46_p 4.54465e-19 $X=0.558 $Y=0.072 $X2=0 $Y2=0
cc_54 VSS N_3_c_24_p 0.00365373f $X=0.576 $Y=0.072 $X2=0 $Y2=0
cc_55 VSS N_3_c_52_p 0.00371671f $X=0.54 $Y=0.0675 $X2=0 $Y2=0
cc_56 VSS N_3_c_25_p 0.00138157f $X=0.592 $Y=0.2025 $X2=0 $Y2=0
cc_57 VSS N_3_c_51_p 0.00260156f $X=0.61 $Y=0.072 $X2=0 $Y2=0
cc_58 VSS N_3_c_58_p 3.97918e-19 $X=0.621 $Y=0.106 $X2=0 $Y2=0
cc_59 VSS N_3_c_52_p 0.00250965f $X=0.54 $Y=0.0675 $X2=0 $Y2=0
cc_60 VSS N_3_c_46_p 0.00365373f $X=0.558 $Y=0.072 $X2=0 $Y2=0
cc_61 VSS N_3_c_45_p 3.56327e-19 $X=0.234 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_62 VSS N_3_c_44_p 3.56327e-19 $X=0.288 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_63 VSS N_3_c_49_p 3.48201e-19 $X=0.396 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_64 VSS N_3_c_50_p 3.30547e-19 $X=0.447 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_65 VSS N_3_c_65_p 3.30547e-19 $X=0.558 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_66 N_A3_M2_g N_A2_M3_g 0.00344695f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_67 N_A3_c_68_n N_A2_c_83_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_68 N_A3_c_69_n N_A2_c_84_n 0.00392079f $X=0.189 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_69 N_A3_M2_g N_A1_M4_g 2.66145e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_70 N_A3_c_69_n N_Y_c_179_n 2.24689e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_71 VSS N_A3_c_69_n 0.00114532f $X=0.189 $Y=0.135 $X2=0.54 $Y2=0.0675
cc_72 N_A2_M3_g N_A1_M4_g 0.00327995f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_73 N_A2_c_83_n N_A1_c_98_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_74 N_A2_c_84_n N_A1_c_94_n 0.00464977f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_75 N_A2_M3_g N_B1_M5_g 2.71887e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_76 VSS N_A2_c_84_n 0.0011319f $X=0.243 $Y=0.135 $X2=0.54 $Y2=0.0675
cc_77 VSS N_A2_M3_g 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0.341 $Y2=0.2025
cc_78 VSS N_A2_c_84_n 0.00125352f $X=0.243 $Y=0.135 $X2=0.341 $Y2=0.2025
cc_79 VSS N_A2_c_84_n 4.64812e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_80 N_A1_M4_g N_B1_M5_g 0.0036939f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_81 N_A1_c_98_n N_B1_c_110_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_82 N_A1_c_94_n N_B1_c_106_n 0.00406615f $X=0.297 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_83 N_A1_M4_g N_B2_M6_g 3.06651e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_84 VSS N_A1_c_94_n 0.00159458f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_85 N_B1_M5_g N_B2_M6_g 0.00371573f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_86 N_B1_c_110_n N_B2_c_122_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_87 N_B1_c_106_n N_B2_c_119_n 0.00483372f $X=0.351 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_88 N_B1_M5_g N_B3_M7_g 3.06651e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_89 VSS N_B1_M5_g 3.62029e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_90 VSS N_B1_c_106_n 0.0012322f $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_91 N_B2_M6_g N_B3_M7_g 0.0036939f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_92 N_B2_c_122_n N_B3_c_135_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_93 N_B2_c_119_n N_B3_c_132_n 0.00483372f $X=0.405 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_94 N_B2_M6_g N_C2_M8_g 2.71887e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_95 VSS N_B2_M6_g 2.68514e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_96 VSS N_B2_c_119_n 0.00121543f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_97 VSS N_B2_M6_g 2.38303e-19 $X=0.405 $Y=0.0675 $X2=0.307 $Y2=0.2025
cc_98 N_B3_M7_g N_C2_M8_g 0.00333077f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_99 N_B3_c_135_n N_C2_c_147_n 8.86777e-19 $X=0.459 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_100 N_B3_c_132_n N_C2_c_144_n 0.00406615f $X=0.459 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_101 N_B3_M7_g N_C1_M9_g 2.71887e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_102 VSS N_B3_M7_g 3.47199e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_103 VSS N_B3_c_132_n 5.30079e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_104 N_C2_M8_g N_C1_M9_g 0.0036939f $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_105 N_C2_c_147_n N_C1_c_162_n 9.33263e-19 $X=0.513 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_106 N_C2_c_144_n N_C1_c_156_n 0.00477924f $X=0.513 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_107 VSS N_C2_M8_g 3.57119e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_108 VSS N_C2_c_144_n 5.37372e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_109 VSS N_C1_M9_g 2.15135e-19 $X=0.567 $Y=0.0675 $X2=0.592 $Y2=0.2025
cc_110 VSS N_Y_c_173_n 2.23372e-19 $X=0.108 $Y=0.036 $X2=0.54 $Y2=0.0675
cc_111 VSS N_Y_c_171_n 2.93728e-19 $X=0.108 $Y=0.036 $X2=0.54 $Y2=0.0675

* END of "./OA332x2_ASAP7_75t_L.pex.sp.OA332X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA333x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:51:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA333x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA333x1_ASAP7_75t_L.pex.sp.pex"
* File: OA333x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:51:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA333X1_ASAP7_75T_L%3 2 5 7 9 10 13 14 17 19 20 23 24 27 31 35 37 39
+ 44 46 47 48 49 50 54 55 56 57 58 60 62 63 64 65 66 70 79 80 81 87 90 VSS
c57 92 VSS 6.57651e-19 $X=0.099 $Y=0.195
c58 91 VSS 6.23446e-19 $X=0.09 $Y=0.195
c59 90 VSS 0.00204357f $X=0.108 $Y=0.195
c60 87 VSS 0.00412141f $X=0.621 $Y=0.2
c61 86 VSS 0.00112176f $X=0.621 $Y=0.106
c62 85 VSS 9.76731e-19 $X=0.621 $Y=0.225
c63 83 VSS 4.0892e-19 $X=0.585 $Y=0.072
c64 82 VSS 3.28227e-19 $X=0.576 $Y=0.072
c65 81 VSS 1.7724e-19 $X=0.569 $Y=0.072
c66 80 VSS 4.2636e-19 $X=0.558 $Y=0.072
c67 79 VSS 8.46035e-21 $X=0.522 $Y=0.072
c68 78 VSS 3.93699e-19 $X=0.504 $Y=0.072
c69 70 VSS 3.25927e-19 $X=0.486 $Y=0.072
c70 68 VSS 0.00347481f $X=0.612 $Y=0.072
c71 67 VSS 8.36318e-19 $X=0.585 $Y=0.234
c72 66 VSS 0.00142296f $X=0.576 $Y=0.234
c73 65 VSS 0.00344621f $X=0.558 $Y=0.234
c74 64 VSS 0.00142296f $X=0.522 $Y=0.234
c75 63 VSS 0.00329285f $X=0.504 $Y=0.234
c76 62 VSS 0.00142296f $X=0.468 $Y=0.234
c77 61 VSS 0.00688205f $X=0.45 $Y=0.234
c78 60 VSS 0.00142296f $X=0.414 $Y=0.234
c79 59 VSS 2.83817e-19 $X=0.396 $Y=0.234
c80 58 VSS 0.00320869f $X=0.394 $Y=0.234
c81 57 VSS 0.00146362f $X=0.36 $Y=0.234
c82 56 VSS 0.00339482f $X=0.342 $Y=0.234
c83 55 VSS 0.00146362f $X=0.306 $Y=0.234
c84 54 VSS 0.00346424f $X=0.288 $Y=0.234
c85 50 VSS 0.00146362f $X=0.252 $Y=0.234
c86 49 VSS 1.46299e-19 $X=0.234 $Y=0.234
c87 48 VSS 0.00340809f $X=0.232 $Y=0.234
c88 47 VSS 0.00142296f $X=0.198 $Y=0.234
c89 46 VSS 0.0032221f $X=0.18 $Y=0.234
c90 45 VSS 2.39163e-19 $X=0.147 $Y=0.234
c91 44 VSS 0.00151377f $X=0.144 $Y=0.234
c92 43 VSS 0.00171948f $X=0.126 $Y=0.234
c93 39 VSS 0.00329953f $X=0.117 $Y=0.234
c94 38 VSS 0.00606378f $X=0.612 $Y=0.234
c95 37 VSS 0.00229578f $X=0.108 $Y=0.225
c96 35 VSS 4.45367e-19 $X=0.081 $Y=0.175
c97 31 VSS 6.4323e-19 $X=0.081 $Y=0.135
c98 29 VSS 4.25123e-19 $X=0.081 $Y=0.186
c99 27 VSS 0.00251001f $X=0.592 $Y=0.2025
c100 23 VSS 0.0022026f $X=0.27 $Y=0.2025
c101 19 VSS 5.38922e-19 $X=0.287 $Y=0.2025
c102 17 VSS 0.00113516f $X=0.592 $Y=0.0675
c103 13 VSS 0.0023085f $X=0.486 $Y=0.0675
c104 9 VSS 5.91014e-19 $X=0.503 $Y=0.0675
c105 5 VSS 0.0024241f $X=0.081 $Y=0.135
c106 2 VSS 0.0649339f $X=0.081 $Y=0.0675
r107 91 92 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.195 $X2=0.099 $Y2=0.195
r108 90 92 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.195 $X2=0.099 $Y2=0.195
r109 88 91 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.195 $X2=0.09 $Y2=0.195
r110 86 87 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.106 $X2=0.621 $Y2=0.2
r111 85 87 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.2
r112 84 86 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.081 $X2=0.621 $Y2=0.106
r113 82 83 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.072 $X2=0.585 $Y2=0.072
r114 81 82 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.569
+ $Y=0.072 $X2=0.576 $Y2=0.072
r115 80 81 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.072 $X2=0.569 $Y2=0.072
r116 79 80 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.072 $X2=0.558 $Y2=0.072
r117 78 79 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.072 $X2=0.522 $Y2=0.072
r118 76 83 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.072 $X2=0.585 $Y2=0.072
r119 70 78 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.072 $X2=0.504 $Y2=0.072
r120 68 84 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.072 $X2=0.621 $Y2=0.081
r121 68 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.072 $X2=0.594 $Y2=0.072
r122 66 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.234 $X2=0.585 $Y2=0.234
r123 65 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.576 $Y2=0.234
r124 64 65 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.234 $X2=0.558 $Y2=0.234
r125 63 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.522 $Y2=0.234
r126 62 63 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.504 $Y2=0.234
r127 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r128 60 61 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.45 $Y2=0.234
r129 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r130 58 59 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.394
+ $Y=0.234 $X2=0.396 $Y2=0.234
r131 57 58 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.394 $Y2=0.234
r132 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r133 55 56 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.342 $Y2=0.234
r134 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r135 52 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.585 $Y2=0.234
r136 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r137 48 49 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.232
+ $Y=0.234 $X2=0.234 $Y2=0.234
r138 47 48 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.232 $Y2=0.234
r139 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r140 45 46 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.147
+ $Y=0.234 $X2=0.18 $Y2=0.234
r141 44 45 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.147 $Y2=0.234
r142 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r143 41 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.288 $Y2=0.234
r144 41 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.252 $Y2=0.234
r145 39 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.234 $X2=0.126 $Y2=0.234
r146 38 85 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r147 38 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r148 37 39 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.108 $Y=0.225 $X2=0.117 $Y2=0.234
r149 36 90 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.204 $X2=0.108 $Y2=0.195
r150 36 37 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.204 $X2=0.108 $Y2=0.225
r151 34 35 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.164 $X2=0.081 $Y2=0.175
r152 31 34 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.164
r153 29 88 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.186 $X2=0.081 $Y2=0.195
r154 29 35 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.186 $X2=0.081 $Y2=0.175
r155 27 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r156 24 27 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2025 $X2=0.592 $Y2=0.2025
r157 23 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r158 20 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r159 19 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r160 17 76 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.072
+ $X2=0.594 $Y2=0.072
r161 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0675 $X2=0.592 $Y2=0.0675
r162 13 70 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.072
+ $X2=0.486 $Y2=0.072
r163 10 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.486 $Y2=0.0675
r164 9 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.0675 $X2=0.486 $Y2=0.0675
r165 5 31 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r166 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r167 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA333X1_ASAP7_75T_L%C3 2 5 7 10 16 VSS
c11 10 VSS 0.00264963f $X=0.135 $Y=0.135
c12 5 VSS 0.001273f $X=0.135 $Y=0.135
c13 2 VSS 0.0593081f $X=0.135 $Y=0.0675
r14 10 16 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.156
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OA333X1_ASAP7_75T_L%C2 2 5 7 10 16 VSS
c16 16 VSS 5.62086e-19 $X=0.183 $Y=0.154
c17 10 VSS 0.0019135f $X=0.189 $Y=0.135
c18 5 VSS 0.00110916f $X=0.189 $Y=0.135
c19 2 VSS 0.059482f $X=0.189 $Y=0.0675
r20 10 16 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.154
r21 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA333X1_ASAP7_75T_L%C1 2 5 7 10 14 VSS
c12 10 VSS 4.82288e-19 $X=0.243 $Y=0.135
c13 5 VSS 0.00113015f $X=0.243 $Y=0.135
c14 2 VSS 0.0608209f $X=0.243 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OA333X1_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.297 $Y=0.135
c14 5 VSS 0.00111823f $X=0.297 $Y=0.135
c15 2 VSS 0.0617786f $X=0.297 $Y=0.0675
r16 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.154
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OA333X1_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.351 $Y=0.135
c14 5 VSS 0.00112198f $X=0.351 $Y=0.135
c15 2 VSS 0.0616432f $X=0.351 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OA333X1_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c12 10 VSS 7.27237e-19 $X=0.405 $Y=0.135
c13 5 VSS 0.00111185f $X=0.405 $Y=0.135
c14 2 VSS 0.0615515f $X=0.405 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OA333X1_ASAP7_75T_L%A3 2 5 7 10 VSS
c12 10 VSS 7.27237e-19 $X=0.462 $Y=0.119
c13 5 VSS 0.00111774f $X=0.459 $Y=0.135
c14 2 VSS 0.0615416f $X=0.459 $Y=0.0675
r15 10 13 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.119 $X2=0.459 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OA333X1_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c12 10 VSS 4.78074e-19 $X=0.513 $Y=0.135
c13 5 VSS 0.00114557f $X=0.513 $Y=0.135
c14 2 VSS 0.0623815f $X=0.513 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OA333X1_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c9 10 VSS 4.90626e-19 $X=0.567 $Y=0.135
c10 5 VSS 0.00171677f $X=0.567 $Y=0.135
c11 2 VSS 0.0671256f $X=0.567 $Y=0.0675
r12 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.155
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
.ends

.subckt PM_OA333X1_ASAP7_75T_L%Y 1 6 9 14 16 18 22 23 30 VSS
c7 33 VSS 9.17717e-19 $X=0.045 $Y=0.234
c8 32 VSS 0.0032947f $X=0.036 $Y=0.234
c9 30 VSS 0.0030586f $X=0.054 $Y=0.234
c10 25 VSS 9.17717e-19 $X=0.045 $Y=0.036
c11 24 VSS 0.0032947f $X=0.036 $Y=0.036
c12 23 VSS 0.00636224f $X=0.054 $Y=0.036
c13 22 VSS 0.00327906f $X=0.054 $Y=0.036
c14 18 VSS 3.56737e-19 $X=0.027 $Y=0.2145
c15 16 VSS 0.00201583f $X=0.027 $Y=0.115
c16 15 VSS 8.84258e-19 $X=0.027 $Y=0.07
c17 14 VSS 0.00385152f $X=0.03 $Y=0.143
c18 12 VSS 3.3975e-19 $X=0.027 $Y=0.225
c19 9 VSS 0.00676077f $X=0.056 $Y=0.2025
c20 6 VSS 3.7894e-19 $X=0.071 $Y=0.2025
c21 1 VSS 3.7894e-19 $X=0.071 $Y=0.0675
r22 32 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.045 $Y2=0.234
r23 30 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.045 $Y2=0.234
r24 27 32 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.036 $Y2=0.234
r25 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.045 $Y2=0.036
r26 22 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.045 $Y2=0.036
r27 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r28 19 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.036 $Y2=0.036
r29 17 18 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.204 $X2=0.027 $Y2=0.2145
r30 15 16 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.115
r31 14 17 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.143 $X2=0.027 $Y2=0.204
r32 14 16 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.143 $X2=0.027 $Y2=0.115
r33 12 27 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.234
r34 12 18 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.2145
r35 11 19 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.036
r36 11 15 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r37 9 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r38 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
r39 4 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r40 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./OA333x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA333x1_ASAP7_75t_L  VSS VDD C3 C2 C1 B1 B2 B3 A3 A2 A1 Y
* 
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* B3	B3
* B2	B2
* B1	B1
* C1	C1
* C2	C2
* C3	C3
M0 VSS N_3_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 noxref_14 N_C3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_C2_M2_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_14 N_C1_M3_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_15 N_B1_M4_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_14 N_B2_M5_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_15 N_B3_M6_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_3_M7_d N_A3_M7_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 noxref_15 N_A2_M8_g N_3_M8_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 N_3_M9_d N_A1_M9_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M10 VDD N_3_M10_g N_Y_M10_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M11 noxref_16 N_C3_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M12 noxref_17 N_C2_M12_g noxref_16 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.179 $Y=0.162
M13 N_3_M13_d N_C1_M13_g noxref_17 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M14 noxref_18 N_B1_M14_g N_3_M14_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M15 noxref_19 N_B2_M15_g noxref_18 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M16 VDD N_B3_M16_g noxref_19 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M17 noxref_20 N_A3_M17_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M18 noxref_21 N_A2_M18_g noxref_20 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
M19 N_3_M19_d N_A1_M19_g noxref_21 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
*
* 
* .include "OA333x1_ASAP7_75t_L.pex.sp.OA333X1_ASAP7_75T_L.pxi"
* BEGIN of "./OA333x1_ASAP7_75t_L.pex.sp.OA333X1_ASAP7_75T_L.pxi"
* File: OA333x1_ASAP7_75t_L.pex.sp.OA333X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:51:03 2017
* 
x_PM_OA333X1_ASAP7_75T_L%3 N_3_M0_g N_3_c_3_p N_3_M10_g N_3_M8_s N_3_M7_d
+ N_3_c_44_p N_3_M9_d N_3_c_47_p N_3_M14_s N_3_M13_d N_3_c_12_p N_3_M19_d
+ N_3_c_28_p N_3_c_4_p N_3_c_8_p N_3_c_34_p N_3_c_35_p N_3_c_2_p N_3_c_38_p
+ N_3_c_7_p N_3_c_37_p N_3_c_39_p N_3_c_11_p N_3_c_40_p N_3_c_14_p N_3_c_42_p
+ N_3_c_17_p N_3_c_43_p N_3_c_19_p N_3_c_21_p N_3_c_56_p N_3_c_23_p N_3_c_57_p
+ N_3_c_27_p N_3_c_41_p N_3_c_24_p N_3_c_51_p N_3_c_30_p N_3_c_31_p N_3_c_10_p
+ VSS PM_OA333X1_ASAP7_75T_L%3
x_PM_OA333X1_ASAP7_75T_L%C3 N_C3_M1_g N_C3_c_60_n N_C3_M11_g N_C3_c_61_n C3 VSS
+ PM_OA333X1_ASAP7_75T_L%C3
x_PM_OA333X1_ASAP7_75T_L%C2 N_C2_M2_g N_C2_c_75_n N_C2_M12_g N_C2_c_76_n C2 VSS
+ PM_OA333X1_ASAP7_75T_L%C2
x_PM_OA333X1_ASAP7_75T_L%C1 N_C1_M3_g N_C1_c_90_n N_C1_M13_g N_C1_c_86_n C1 VSS
+ PM_OA333X1_ASAP7_75T_L%C1
x_PM_OA333X1_ASAP7_75T_L%B1 N_B1_M4_g N_B1_c_102_n N_B1_M14_g N_B1_c_98_n B1 VSS
+ PM_OA333X1_ASAP7_75T_L%B1
x_PM_OA333X1_ASAP7_75T_L%B2 N_B2_M5_g N_B2_c_114_n N_B2_M15_g N_B2_c_111_n B2
+ VSS PM_OA333X1_ASAP7_75T_L%B2
x_PM_OA333X1_ASAP7_75T_L%B3 N_B3_M6_g N_B3_c_127_n N_B3_M16_g N_B3_c_124_n B3
+ VSS PM_OA333X1_ASAP7_75T_L%B3
x_PM_OA333X1_ASAP7_75T_L%A3 N_A3_M7_g N_A3_c_139_n N_A3_M17_g A3 VSS
+ PM_OA333X1_ASAP7_75T_L%A3
x_PM_OA333X1_ASAP7_75T_L%A2 N_A2_M8_g N_A2_c_153_n N_A2_M18_g N_A2_c_149_n A2
+ VSS PM_OA333X1_ASAP7_75T_L%A2
x_PM_OA333X1_ASAP7_75T_L%A1 N_A1_M9_g N_A1_c_166_n N_A1_M19_g N_A1_c_160_n A1
+ VSS PM_OA333X1_ASAP7_75T_L%A1
x_PM_OA333X1_ASAP7_75T_L%Y N_Y_M0_s N_Y_M10_s N_Y_c_168_n Y N_Y_c_172_n
+ N_Y_c_170_n N_Y_c_174_p N_Y_c_173_p N_Y_c_171_n VSS PM_OA333X1_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_C3_M1_g 0.00284417f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_3_c_2_p N_C3_M1_g 2.40674e-19 $X=0.144 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_3 N_3_c_3_p N_C3_c_60_n 9.34529e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_3_c_4_p N_C3_c_61_n 0.00216032f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_5 N_3_c_2_p N_C3_c_61_n 2.68686e-19 $X=0.144 $Y=0.234 $X2=0.135 $Y2=0.135
cc_6 N_3_M0_g N_C2_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_7 N_3_c_7_p N_C2_M2_g 3.38929e-19 $X=0.198 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_8 N_3_c_8_p C2 2.35508e-19 $X=0.081 $Y=0.175 $X2=0.127 $Y2=0.156
cc_9 N_3_c_7_p C2 0.00123604f $X=0.198 $Y=0.234 $X2=0.127 $Y2=0.156
cc_10 N_3_c_10_p C2 4.18335e-19 $X=0.108 $Y=0.195 $X2=0.127 $Y2=0.156
cc_11 N_3_c_11_p N_C1_M3_g 2.64276e-19 $X=0.252 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_12 N_3_c_12_p N_C1_c_86_n 0.0013295f $X=0.27 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_13 N_3_c_11_p N_C1_c_86_n 0.00124805f $X=0.252 $Y=0.234 $X2=0.135 $Y2=0.135
cc_14 N_3_c_14_p N_B1_M4_g 2.64276e-19 $X=0.306 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_15 N_3_c_12_p N_B1_c_98_n 0.0013295f $X=0.27 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_16 N_3_c_14_p N_B1_c_98_n 0.00124805f $X=0.306 $Y=0.234 $X2=0.135 $Y2=0.135
cc_17 N_3_c_17_p N_B2_M5_g 3.48613e-19 $X=0.36 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_18 N_3_c_17_p N_B2_c_111_n 0.00124805f $X=0.36 $Y=0.234 $X2=0.135 $Y2=0.135
cc_19 N_3_c_19_p N_B3_M6_g 2.56935e-19 $X=0.414 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_20 N_3_c_19_p N_B3_c_124_n 0.00123064f $X=0.414 $Y=0.234 $X2=0.135 $Y2=0.135
cc_21 N_3_c_21_p N_A3_M7_g 2.45924e-19 $X=0.468 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_22 N_3_c_21_p A3 0.00123064f $X=0.468 $Y=0.234 $X2=0.135 $Y2=0.135
cc_23 N_3_c_23_p N_A2_M8_g 3.38929e-19 $X=0.522 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_24 N_3_c_24_p N_A2_M8_g 2.76185e-19 $X=0.522 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_25 N_3_c_23_p N_A2_c_149_n 0.00123064f $X=0.522 $Y=0.234 $X2=0.135 $Y2=0.135
cc_26 N_3_c_24_p N_A2_c_149_n 0.0012322f $X=0.522 $Y=0.072 $X2=0.135 $Y2=0.135
cc_27 N_3_c_27_p N_A1_M9_g 2.56935e-19 $X=0.576 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_28 N_3_c_28_p N_A1_c_160_n 0.0013295f $X=0.592 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_29 N_3_c_27_p N_A1_c_160_n 0.00123064f $X=0.576 $Y=0.234 $X2=0.135 $Y2=0.135
cc_30 N_3_c_30_p N_A1_c_160_n 0.00121543f $X=0.569 $Y=0.072 $X2=0.135 $Y2=0.135
cc_31 N_3_c_31_p N_A1_c_160_n 0.00392202f $X=0.621 $Y=0.2 $X2=0.135 $Y2=0.135
cc_32 N_3_c_4_p N_Y_c_168_n 0.00125175f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_33 N_3_c_4_p Y 0.0036413f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_34 N_3_c_34_p N_Y_c_170_n 2.71869e-19 $X=0.108 $Y=0.225 $X2=0 $Y2=0
cc_35 N_3_c_35_p N_Y_c_171_n 9.1444e-19 $X=0.117 $Y=0.234 $X2=0 $Y2=0
cc_36 VSS N_3_c_12_p 0.00138157f $X=0.27 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_37 VSS N_3_c_37_p 2.20236e-19 $X=0.232 $Y=0.234 $X2=0.127 $Y2=0.156
cc_38 VSS N_3_c_38_p 2.20236e-19 $X=0.18 $Y=0.234 $X2=0 $Y2=0
cc_39 VSS N_3_c_39_p 2.30729e-19 $X=0.234 $Y=0.234 $X2=0 $Y2=0
cc_40 VSS N_3_c_40_p 2.30729e-19 $X=0.288 $Y=0.234 $X2=0 $Y2=0
cc_41 VSS N_3_c_41_p 3.14723e-19 $X=0.486 $Y=0.072 $X2=0 $Y2=0
cc_42 VSS N_3_c_42_p 2.30729e-19 $X=0.342 $Y=0.234 $X2=0 $Y2=0
cc_43 VSS N_3_c_43_p 2.30729e-19 $X=0.394 $Y=0.234 $X2=0 $Y2=0
cc_44 VSS N_3_c_44_p 0.003332f $X=0.486 $Y=0.0675 $X2=0 $Y2=0
cc_45 VSS N_3_c_41_p 4.6373e-19 $X=0.486 $Y=0.072 $X2=0 $Y2=0
cc_46 VSS N_3_c_44_p 0.00250965f $X=0.486 $Y=0.0675 $X2=0 $Y2=0
cc_47 VSS N_3_c_47_p 3.14809e-19 $X=0.592 $Y=0.0675 $X2=0 $Y2=0
cc_48 VSS N_3_c_41_p 0.00881219f $X=0.486 $Y=0.072 $X2=0 $Y2=0
cc_49 VSS N_3_c_44_p 0.00355403f $X=0.486 $Y=0.0675 $X2=0 $Y2=0
cc_50 VSS N_3_c_47_p 0.00337424f $X=0.592 $Y=0.0675 $X2=0 $Y2=0
cc_51 VSS N_3_c_51_p 0.00233206f $X=0.558 $Y=0.072 $X2=0 $Y2=0
cc_52 VSS N_3_c_38_p 3.41091e-19 $X=0.18 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_53 VSS N_3_c_37_p 3.56327e-19 $X=0.232 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_54 VSS N_3_c_42_p 3.34078e-19 $X=0.342 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_55 VSS N_3_c_43_p 3.4467e-19 $X=0.394 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_56 VSS N_3_c_56_p 3.48201e-19 $X=0.504 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_57 VSS N_3_c_57_p 3.48201e-19 $X=0.558 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_58 N_C3_M1_g N_C2_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_59 N_C3_c_60_n N_C2_c_75_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_60 N_C3_c_61_n N_C2_c_76_n 0.00392079f $X=0.135 $Y=0.135 $X2=0.469 $Y2=0.0675
cc_61 N_C3_M1_g N_C1_M3_g 2.66145e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_62 N_C3_c_61_n N_Y_c_172_n 4.286e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_63 VSS N_C3_c_61_n 0.00114532f $X=0.135 $Y=0.135 $X2=0.287 $Y2=0.2025
cc_64 N_C2_M2_g N_C1_M3_g 0.00327995f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_65 N_C2_c_75_n N_C1_c_90_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_66 N_C2_c_76_n N_C1_c_86_n 0.0046535f $X=0.189 $Y=0.135 $X2=0.469 $Y2=0.0675
cc_67 N_C2_M2_g N_B1_M4_g 2.71887e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_68 VSS N_C2_c_76_n 0.0011319f $X=0.189 $Y=0.135 $X2=0.287 $Y2=0.2025
cc_69 VSS N_C2_M2_g 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_70 VSS N_C2_c_76_n 0.00125352f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_71 VSS N_C2_c_76_n 5.07686e-19 $X=0.189 $Y=0.135 $X2=0.592 $Y2=0.2025
cc_72 N_C1_M3_g N_B1_M4_g 0.0036939f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_73 N_C1_c_90_n N_B1_c_102_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_74 N_C1_c_86_n N_B1_c_98_n 0.00406615f $X=0.243 $Y=0.135 $X2=0.469 $Y2=0.0675
cc_75 N_C1_M3_g N_B2_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_76 VSS N_C1_c_86_n 0.00151583f $X=0.243 $Y=0.135 $X2=0.592 $Y2=0.2025
cc_77 N_B1_M4_g N_B2_M5_g 0.00371573f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_78 N_B1_c_102_n N_B2_c_114_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_79 N_B1_c_98_n N_B2_c_111_n 0.00483372f $X=0.297 $Y=0.135 $X2=0.469
+ $Y2=0.0675
cc_80 N_B1_M4_g N_B3_M6_g 3.06651e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_81 VSS N_B1_M4_g 3.62029e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.175
cc_82 VSS N_B1_c_98_n 0.0012322f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.175
cc_83 N_B2_M5_g N_B3_M6_g 0.0036939f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_84 N_B2_c_114_n N_B3_c_127_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_85 N_B2_c_111_n N_B3_c_124_n 0.00483372f $X=0.351 $Y=0.135 $X2=0.469
+ $Y2=0.0675
cc_86 N_B2_M5_g N_A3_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_87 VSS N_B2_M5_g 2.68514e-19 $X=0.351 $Y=0.0675 $X2=0.612 $Y2=0.234
cc_88 VSS N_B2_c_111_n 0.00121543f $X=0.351 $Y=0.135 $X2=0.612 $Y2=0.234
cc_89 VSS N_B2_M5_g 2.38303e-19 $X=0.351 $Y=0.0675 $X2=0.27 $Y2=0.2025
cc_90 N_B3_M6_g N_A3_M7_g 0.00333077f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_91 N_B3_c_127_n N_A3_c_139_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_92 N_B3_c_124_n A3 0.00406615f $X=0.405 $Y=0.135 $X2=0.469 $Y2=0.0675
cc_93 N_B3_M6_g N_A2_M8_g 2.71887e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_94 VSS N_B3_M6_g 3.47199e-19 $X=0.405 $Y=0.0675 $X2=0.592 $Y2=0.2025
cc_95 VSS N_B3_c_124_n 5.30079e-19 $X=0.405 $Y=0.135 $X2=0.592 $Y2=0.2025
cc_96 N_A3_M7_g N_A2_M8_g 0.0036939f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_97 N_A3_c_139_n N_A2_c_153_n 8.86777e-19 $X=0.459 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_98 A3 N_A2_c_149_n 0.00483372f $X=0.462 $Y=0.119 $X2=0.469 $Y2=0.0675
cc_99 N_A3_M7_g N_A1_M9_g 3.06651e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_100 VSS N_A3_M7_g 3.37279e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_101 VSS A3 5.22785e-19 $X=0.462 $Y=0.119 $X2=0.081 $Y2=0.135
cc_102 N_A2_M8_g N_A1_M9_g 0.00376655f $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_103 N_A2_c_153_n N_A1_c_166_n 9.33263e-19 $X=0.513 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_104 N_A2_c_149_n N_A1_c_160_n 0.0048308f $X=0.513 $Y=0.135 $X2=0.469
+ $Y2=0.0675
cc_105 VSS N_A2_M8_g 2.38303e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_106 VSS N_Y_c_173_p 2.87474e-19 $X=0.054 $Y=0.036 $X2=0.287 $Y2=0.2025
cc_107 VSS N_Y_c_174_p 2.75937e-19 $X=0.054 $Y=0.036 $X2=0.27 $Y2=0.2025

* END of "./OA333x1_ASAP7_75t_L.pex.sp.OA333X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA333x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:51:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA333x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA333x2_ASAP7_75t_L.pex.sp.pex"
* File: OA333x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:51:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA333X2_ASAP7_75T_L%3 2 7 10 13 15 17 18 21 22 25 27 28 31 32 35 39
+ 43 47 52 54 55 56 57 58 62 63 64 65 66 68 70 71 72 73 74 78 87 88 89 95 98 VSS
c65 100 VSS 6.57651e-19 $X=0.153 $Y=0.195
c66 99 VSS 6.23446e-19 $X=0.144 $Y=0.195
c67 98 VSS 0.00204357f $X=0.162 $Y=0.195
c68 95 VSS 0.00412141f $X=0.675 $Y=0.2
c69 94 VSS 0.00112176f $X=0.675 $Y=0.106
c70 93 VSS 9.76731e-19 $X=0.675 $Y=0.225
c71 91 VSS 4.0892e-19 $X=0.639 $Y=0.072
c72 90 VSS 3.28227e-19 $X=0.63 $Y=0.072
c73 89 VSS 1.7724e-19 $X=0.623 $Y=0.072
c74 88 VSS 4.2636e-19 $X=0.612 $Y=0.072
c75 87 VSS 8.46035e-21 $X=0.576 $Y=0.072
c76 86 VSS 3.93699e-19 $X=0.558 $Y=0.072
c77 78 VSS 3.25927e-19 $X=0.54 $Y=0.072
c78 76 VSS 0.00347481f $X=0.666 $Y=0.072
c79 75 VSS 8.36318e-19 $X=0.639 $Y=0.234
c80 74 VSS 0.00142296f $X=0.63 $Y=0.234
c81 73 VSS 0.00344621f $X=0.612 $Y=0.234
c82 72 VSS 0.00142296f $X=0.576 $Y=0.234
c83 71 VSS 0.00329285f $X=0.558 $Y=0.234
c84 70 VSS 0.00142296f $X=0.522 $Y=0.234
c85 69 VSS 0.00688205f $X=0.504 $Y=0.234
c86 68 VSS 0.00142296f $X=0.468 $Y=0.234
c87 67 VSS 2.83817e-19 $X=0.45 $Y=0.234
c88 66 VSS 0.00320869f $X=0.448 $Y=0.234
c89 65 VSS 0.00146362f $X=0.414 $Y=0.234
c90 64 VSS 0.00339482f $X=0.396 $Y=0.234
c91 63 VSS 0.00146362f $X=0.36 $Y=0.234
c92 62 VSS 0.00346424f $X=0.342 $Y=0.234
c93 58 VSS 0.00146362f $X=0.306 $Y=0.234
c94 57 VSS 1.46299e-19 $X=0.288 $Y=0.234
c95 56 VSS 0.00340809f $X=0.286 $Y=0.234
c96 55 VSS 0.00142296f $X=0.252 $Y=0.234
c97 54 VSS 0.0032221f $X=0.234 $Y=0.234
c98 53 VSS 2.39163e-19 $X=0.201 $Y=0.234
c99 52 VSS 0.00151377f $X=0.198 $Y=0.234
c100 51 VSS 0.00171948f $X=0.18 $Y=0.234
c101 47 VSS 0.00318978f $X=0.171 $Y=0.234
c102 46 VSS 0.00606378f $X=0.666 $Y=0.234
c103 45 VSS 0.00196286f $X=0.162 $Y=0.225
c104 43 VSS 4.45367e-19 $X=0.135 $Y=0.175
c105 39 VSS 5.9584e-19 $X=0.135 $Y=0.135
c106 37 VSS 4.25123e-19 $X=0.135 $Y=0.186
c107 35 VSS 0.00251001f $X=0.646 $Y=0.2025
c108 31 VSS 0.0022026f $X=0.324 $Y=0.2025
c109 27 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c110 25 VSS 0.00113516f $X=0.646 $Y=0.0675
c111 21 VSS 0.0023085f $X=0.54 $Y=0.0675
c112 17 VSS 5.91014e-19 $X=0.557 $Y=0.0675
c113 13 VSS 0.00437781f $X=0.135 $Y=0.135
c114 10 VSS 0.0609638f $X=0.135 $Y=0.0675
c115 2 VSS 0.0639847f $X=0.081 $Y=0.0675
r116 99 100 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.195 $X2=0.153 $Y2=0.195
r117 98 100 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.195 $X2=0.153 $Y2=0.195
r118 96 99 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.195 $X2=0.144 $Y2=0.195
r119 94 95 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.106 $X2=0.675 $Y2=0.2
r120 93 95 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.225 $X2=0.675 $Y2=0.2
r121 92 94 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.081 $X2=0.675 $Y2=0.106
r122 90 91 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.072 $X2=0.639 $Y2=0.072
r123 89 90 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.623
+ $Y=0.072 $X2=0.63 $Y2=0.072
r124 88 89 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.072 $X2=0.623 $Y2=0.072
r125 87 88 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.072 $X2=0.612 $Y2=0.072
r126 86 87 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.072 $X2=0.576 $Y2=0.072
r127 84 91 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.072 $X2=0.639 $Y2=0.072
r128 78 86 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.072 $X2=0.558 $Y2=0.072
r129 76 92 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.072 $X2=0.675 $Y2=0.081
r130 76 84 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.072 $X2=0.648 $Y2=0.072
r131 74 75 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.234 $X2=0.639 $Y2=0.234
r132 73 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.63 $Y2=0.234
r133 72 73 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.234 $X2=0.612 $Y2=0.234
r134 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.576 $Y2=0.234
r135 70 71 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.234 $X2=0.558 $Y2=0.234
r136 69 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.522 $Y2=0.234
r137 68 69 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.504 $Y2=0.234
r138 67 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r139 66 67 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.448
+ $Y=0.234 $X2=0.45 $Y2=0.234
r140 65 66 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.448 $Y2=0.234
r141 64 65 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r142 63 64 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.396 $Y2=0.234
r143 62 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r144 60 75 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.639 $Y2=0.234
r145 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r146 56 57 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.286
+ $Y=0.234 $X2=0.288 $Y2=0.234
r147 55 56 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.286 $Y2=0.234
r148 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r149 53 54 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.201
+ $Y=0.234 $X2=0.234 $Y2=0.234
r150 52 53 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.201 $Y2=0.234
r151 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r152 49 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.342 $Y2=0.234
r153 49 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.306 $Y2=0.234
r154 47 51 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.234 $X2=0.18 $Y2=0.234
r155 46 93 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.234 $X2=0.675 $Y2=0.225
r156 46 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.234 $X2=0.648 $Y2=0.234
r157 45 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.225 $X2=0.171 $Y2=0.234
r158 44 98 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.204 $X2=0.162 $Y2=0.195
r159 44 45 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.204 $X2=0.162 $Y2=0.225
r160 42 43 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.164 $X2=0.135 $Y2=0.175
r161 39 42 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.164
r162 37 96 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.186 $X2=0.135 $Y2=0.195
r163 37 43 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.186 $X2=0.135 $Y2=0.175
r164 35 60 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234
+ $X2=0.648 $Y2=0.234
r165 32 35 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.646 $Y2=0.2025
r166 31 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r167 28 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r168 27 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r169 25 84 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.072
+ $X2=0.648 $Y2=0.072
r170 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.646 $Y2=0.0675
r171 21 78 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.072 $X2=0.54
+ $Y2=0.072
r172 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r173 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r174 13 39 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r175 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r176 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r177 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r178 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r179 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA333X2_ASAP7_75T_L%C3 2 5 7 10 16 VSS
c12 10 VSS 0.00283088f $X=0.189 $Y=0.135
c13 5 VSS 0.00115289f $X=0.189 $Y=0.135
c14 2 VSS 0.0585388f $X=0.189 $Y=0.0675
r15 10 16 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.156
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA333X2_ASAP7_75T_L%C2 2 5 7 10 16 VSS
c16 16 VSS 5.62086e-19 $X=0.237 $Y=0.154
c17 10 VSS 0.0019135f $X=0.243 $Y=0.135
c18 5 VSS 0.0011122f $X=0.243 $Y=0.135
c19 2 VSS 0.059482f $X=0.243 $Y=0.0675
r20 10 16 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.154
r21 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OA333X2_ASAP7_75T_L%C1 2 5 7 10 14 VSS
c12 10 VSS 4.82288e-19 $X=0.297 $Y=0.135
c13 5 VSS 0.00113015f $X=0.297 $Y=0.135
c14 2 VSS 0.0608209f $X=0.297 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OA333X2_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.351 $Y=0.135
c14 5 VSS 0.00111823f $X=0.351 $Y=0.135
c15 2 VSS 0.0617786f $X=0.351 $Y=0.0675
r16 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.154
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OA333X2_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.405 $Y=0.135
c14 5 VSS 0.00112198f $X=0.405 $Y=0.135
c15 2 VSS 0.0616432f $X=0.405 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OA333X2_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c12 10 VSS 7.27237e-19 $X=0.459 $Y=0.135
c13 5 VSS 0.00111185f $X=0.459 $Y=0.135
c14 2 VSS 0.0615515f $X=0.459 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OA333X2_ASAP7_75T_L%A3 2 5 7 10 VSS
c12 10 VSS 7.27237e-19 $X=0.516 $Y=0.119
c13 5 VSS 0.00111774f $X=0.513 $Y=0.135
c14 2 VSS 0.0615416f $X=0.513 $Y=0.0675
r15 10 13 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.119 $X2=0.513 $Y2=0.135
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OA333X2_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c12 10 VSS 4.78074e-19 $X=0.567 $Y=0.135
c13 5 VSS 0.00114557f $X=0.567 $Y=0.135
c14 2 VSS 0.0623815f $X=0.567 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
.ends

.subckt PM_OA333X2_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c9 10 VSS 4.90626e-19 $X=0.621 $Y=0.135
c10 5 VSS 0.00171677f $X=0.621 $Y=0.135
c11 2 VSS 0.0671256f $X=0.621 $Y=0.0675
r12 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.155
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
.ends

.subckt PM_OA333X2_ASAP7_75T_L%Y 1 2 6 7 10 14 16 21 22 26 VSS
c14 26 VSS 0.00659662f $X=0.108 $Y=0.234
c15 24 VSS 0.00385179f $X=0.063 $Y=0.234
c16 22 VSS 0.00894858f $X=0.108 $Y=0.036
c17 21 VSS 0.00681978f $X=0.108 $Y=0.036
c18 19 VSS 0.00385179f $X=0.063 $Y=0.036
c19 18 VSS 9.92723e-19 $X=0.054 $Y=0.2145
c20 16 VSS 0.00422063f $X=0.054 $Y=0.115
c21 15 VSS 0.00219361f $X=0.054 $Y=0.07
c22 14 VSS 0.00602261f $X=0.057 $Y=0.143
c23 12 VSS 9.44835e-19 $X=0.054 $Y=0.225
c24 10 VSS 0.0101881f $X=0.108 $Y=0.2025
c25 6 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c26 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r27 24 26 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.234 $X2=0.108 $Y2=0.234
r28 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r29 19 21 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.036 $X2=0.108 $Y2=0.036
r30 17 18 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.204 $X2=0.054 $Y2=0.2145
r31 15 16 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.07 $X2=0.054 $Y2=0.115
r32 14 17 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.143 $X2=0.054 $Y2=0.204
r33 14 16 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.143 $X2=0.054 $Y2=0.115
r34 12 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.054 $Y=0.225 $X2=0.063 $Y2=0.234
r35 12 18 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.225 $X2=0.054 $Y2=0.2145
r36 11 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.054 $Y=0.045 $X2=0.063 $Y2=0.036
r37 11 15 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.045 $X2=0.054 $Y2=0.07
r38 10 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r39 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r40 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r41 5 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r42 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r43 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OA333x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA333x2_ASAP7_75t_L  VSS VDD C3 C2 C1 B1 B2 B3 A3 A2 A1 Y
* 
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* B3	B3
* B2	B2
* B1	B1
* C1	C1
* C2	C2
* C3	C3
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_14 N_C3_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_C2_M3_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_14 N_C1_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_15 N_B1_M5_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_14 N_B2_M6_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_15 N_B3_M7_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_3_M8_d N_A3_M8_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 noxref_15 N_A2_M9_g N_3_M9_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M10 N_3_M10_d N_A1_M10_g noxref_15 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.611 $Y=0.027
M11 N_Y_M11_d N_3_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M12 N_Y_M12_d N_3_M12_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M13 noxref_16 N_C3_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M14 noxref_17 N_C2_M14_g noxref_16 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M15 N_3_M15_d N_C1_M15_g noxref_17 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M16 noxref_18 N_B1_M16_g N_3_M16_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M17 noxref_19 N_B2_M17_g noxref_18 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M18 VDD N_B3_M18_g noxref_19 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M19 noxref_20 N_A3_M19_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M20 noxref_21 N_A2_M20_g noxref_20 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M21 N_3_M21_d N_A1_M21_g noxref_21 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.611 $Y=0.162
*
* 
* .include "OA333x2_ASAP7_75t_L.pex.sp.OA333X2_ASAP7_75T_L.pxi"
* BEGIN of "./OA333x2_ASAP7_75t_L.pex.sp.OA333X2_ASAP7_75T_L.pxi"
* File: OA333x2_ASAP7_75t_L.pex.sp.OA333X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:51:26 2017
* 
x_PM_OA333X2_ASAP7_75T_L%3 N_3_M0_g N_3_M11_g N_3_M1_g N_3_c_4_p N_3_M12_g
+ N_3_M9_s N_3_M8_d N_3_c_52_p N_3_M10_d N_3_c_55_p N_3_M16_s N_3_M15_d
+ N_3_c_13_p N_3_M21_d N_3_c_29_p N_3_c_5_p N_3_c_9_p N_3_c_43_p N_3_c_3_p
+ N_3_c_46_p N_3_c_8_p N_3_c_45_p N_3_c_47_p N_3_c_12_p N_3_c_48_p N_3_c_15_p
+ N_3_c_50_p N_3_c_18_p N_3_c_51_p N_3_c_20_p N_3_c_22_p N_3_c_64_p N_3_c_24_p
+ N_3_c_65_p N_3_c_28_p N_3_c_49_p N_3_c_25_p N_3_c_59_p N_3_c_31_p N_3_c_32_p
+ N_3_c_11_p VSS PM_OA333X2_ASAP7_75T_L%3
x_PM_OA333X2_ASAP7_75T_L%C3 N_C3_M2_g N_C3_c_69_n N_C3_M13_g N_C3_c_70_n C3 VSS
+ PM_OA333X2_ASAP7_75T_L%C3
x_PM_OA333X2_ASAP7_75T_L%C2 N_C2_M3_g N_C2_c_84_n N_C2_M14_g N_C2_c_85_n C2 VSS
+ PM_OA333X2_ASAP7_75T_L%C2
x_PM_OA333X2_ASAP7_75T_L%C1 N_C1_M4_g N_C1_c_99_n N_C1_M15_g N_C1_c_95_n C1 VSS
+ PM_OA333X2_ASAP7_75T_L%C1
x_PM_OA333X2_ASAP7_75T_L%B1 N_B1_M5_g N_B1_c_111_n N_B1_M16_g N_B1_c_107_n B1
+ VSS PM_OA333X2_ASAP7_75T_L%B1
x_PM_OA333X2_ASAP7_75T_L%B2 N_B2_M6_g N_B2_c_123_n N_B2_M17_g N_B2_c_120_n B2
+ VSS PM_OA333X2_ASAP7_75T_L%B2
x_PM_OA333X2_ASAP7_75T_L%B3 N_B3_M7_g N_B3_c_136_n N_B3_M18_g N_B3_c_133_n B3
+ VSS PM_OA333X2_ASAP7_75T_L%B3
x_PM_OA333X2_ASAP7_75T_L%A3 N_A3_M8_g N_A3_c_148_n N_A3_M19_g A3 VSS
+ PM_OA333X2_ASAP7_75T_L%A3
x_PM_OA333X2_ASAP7_75T_L%A2 N_A2_M9_g N_A2_c_162_n N_A2_M20_g N_A2_c_158_n A2
+ VSS PM_OA333X2_ASAP7_75T_L%A2
x_PM_OA333X2_ASAP7_75T_L%A1 N_A1_M10_g N_A1_c_175_n N_A1_M21_g N_A1_c_169_n A1
+ VSS PM_OA333X2_ASAP7_75T_L%A1
x_PM_OA333X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_M12_d N_Y_M11_d N_Y_c_179_n Y
+ N_Y_c_188_n N_Y_c_182_n N_Y_c_184_n N_Y_c_185_n VSS PM_OA333X2_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_C3_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_C3_M2_g 0.00284417f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_C3_M2_g 2.40674e-19 $X=0.198 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_4 N_3_c_4_p N_C3_c_69_n 9.59383e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_5 N_3_c_5_p N_C3_c_70_n 0.00216301f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_6 N_3_c_3_p N_C3_c_70_n 2.68686e-19 $X=0.198 $Y=0.234 $X2=0.189 $Y2=0.135
cc_7 N_3_M1_g N_C2_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_8 N_3_c_8_p N_C2_M3_g 3.38929e-19 $X=0.252 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_9 N_3_c_9_p C2 2.35508e-19 $X=0.135 $Y=0.175 $X2=0.181 $Y2=0.156
cc_10 N_3_c_8_p C2 0.00123604f $X=0.252 $Y=0.234 $X2=0.181 $Y2=0.156
cc_11 N_3_c_11_p C2 4.18335e-19 $X=0.162 $Y=0.195 $X2=0.181 $Y2=0.156
cc_12 N_3_c_12_p N_C1_M4_g 2.64276e-19 $X=0.306 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_13 N_3_c_13_p N_C1_c_95_n 0.0013295f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_14 N_3_c_12_p N_C1_c_95_n 0.00124805f $X=0.306 $Y=0.234 $X2=0.189 $Y2=0.135
cc_15 N_3_c_15_p N_B1_M5_g 2.64276e-19 $X=0.36 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_16 N_3_c_13_p N_B1_c_107_n 0.0013295f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_17 N_3_c_15_p N_B1_c_107_n 0.00124805f $X=0.36 $Y=0.234 $X2=0.189 $Y2=0.135
cc_18 N_3_c_18_p N_B2_M6_g 3.48613e-19 $X=0.414 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_19 N_3_c_18_p N_B2_c_120_n 0.00124805f $X=0.414 $Y=0.234 $X2=0.189 $Y2=0.135
cc_20 N_3_c_20_p N_B3_M7_g 2.56935e-19 $X=0.468 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_21 N_3_c_20_p N_B3_c_133_n 0.00123064f $X=0.468 $Y=0.234 $X2=0.189 $Y2=0.135
cc_22 N_3_c_22_p N_A3_M8_g 2.45924e-19 $X=0.522 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_23 N_3_c_22_p A3 0.00123064f $X=0.522 $Y=0.234 $X2=0.189 $Y2=0.135
cc_24 N_3_c_24_p N_A2_M9_g 3.38929e-19 $X=0.576 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_25 N_3_c_25_p N_A2_M9_g 2.76185e-19 $X=0.576 $Y=0.072 $X2=0.189 $Y2=0.0675
cc_26 N_3_c_24_p N_A2_c_158_n 0.00123064f $X=0.576 $Y=0.234 $X2=0.189 $Y2=0.135
cc_27 N_3_c_25_p N_A2_c_158_n 0.0012322f $X=0.576 $Y=0.072 $X2=0.189 $Y2=0.135
cc_28 N_3_c_28_p N_A1_M10_g 2.56935e-19 $X=0.63 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_29 N_3_c_29_p N_A1_c_169_n 0.0013295f $X=0.646 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_30 N_3_c_28_p N_A1_c_169_n 0.00123064f $X=0.63 $Y=0.234 $X2=0.189 $Y2=0.135
cc_31 N_3_c_31_p N_A1_c_169_n 0.00121543f $X=0.623 $Y=0.072 $X2=0.189 $Y2=0.135
cc_32 N_3_c_32_p N_A1_c_169_n 0.00392202f $X=0.675 $Y=0.2 $X2=0.189 $Y2=0.135
cc_33 N_3_c_4_p N_Y_M1_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_34 N_3_c_4_p N_Y_M12_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_35 N_3_c_4_p N_Y_c_179_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_36 N_3_c_5_p N_Y_c_179_n 0.00141343f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_37 N_3_c_5_p Y 0.00193798f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_38 N_3_M0_g N_Y_c_182_n 4.59284e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_3_c_4_p N_Y_c_182_n 5.51214e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_40 N_3_c_4_p N_Y_c_184_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_41 N_3_M0_g N_Y_c_185_n 4.59284e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_42 N_3_c_4_p N_Y_c_185_n 5.51214e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_43 N_3_c_43_p N_Y_c_185_n 9.4488e-19 $X=0.171 $Y=0.234 $X2=0 $Y2=0
cc_44 VSS N_3_c_13_p 0.00138157f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.135
cc_45 VSS N_3_c_45_p 2.20236e-19 $X=0.286 $Y=0.234 $X2=0.181 $Y2=0.156
cc_46 VSS N_3_c_46_p 2.20236e-19 $X=0.234 $Y=0.234 $X2=0 $Y2=0
cc_47 VSS N_3_c_47_p 2.30729e-19 $X=0.288 $Y=0.234 $X2=0 $Y2=0
cc_48 VSS N_3_c_48_p 2.30729e-19 $X=0.342 $Y=0.234 $X2=0 $Y2=0
cc_49 VSS N_3_c_49_p 3.14723e-19 $X=0.54 $Y=0.072 $X2=0 $Y2=0
cc_50 VSS N_3_c_50_p 2.30729e-19 $X=0.396 $Y=0.234 $X2=0 $Y2=0
cc_51 VSS N_3_c_51_p 2.30729e-19 $X=0.448 $Y=0.234 $X2=0 $Y2=0
cc_52 VSS N_3_c_52_p 0.003332f $X=0.54 $Y=0.0675 $X2=0 $Y2=0
cc_53 VSS N_3_c_49_p 4.6373e-19 $X=0.54 $Y=0.072 $X2=0 $Y2=0
cc_54 VSS N_3_c_52_p 0.00250965f $X=0.54 $Y=0.0675 $X2=0 $Y2=0
cc_55 VSS N_3_c_55_p 3.14809e-19 $X=0.646 $Y=0.0675 $X2=0 $Y2=0
cc_56 VSS N_3_c_49_p 0.00881219f $X=0.54 $Y=0.072 $X2=0 $Y2=0
cc_57 VSS N_3_c_52_p 0.00355403f $X=0.54 $Y=0.0675 $X2=0 $Y2=0
cc_58 VSS N_3_c_55_p 0.00337424f $X=0.646 $Y=0.0675 $X2=0 $Y2=0
cc_59 VSS N_3_c_59_p 0.00233206f $X=0.612 $Y=0.072 $X2=0 $Y2=0
cc_60 VSS N_3_c_46_p 3.41091e-19 $X=0.234 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_61 VSS N_3_c_45_p 3.56327e-19 $X=0.286 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_62 VSS N_3_c_50_p 3.34078e-19 $X=0.396 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_63 VSS N_3_c_51_p 3.4467e-19 $X=0.448 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_64 VSS N_3_c_64_p 3.48201e-19 $X=0.558 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_65 VSS N_3_c_65_p 3.48201e-19 $X=0.612 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_66 N_C3_M2_g N_C2_M3_g 0.00344695f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_67 N_C3_c_69_n N_C2_c_84_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_68 N_C3_c_70_n N_C2_c_85_n 0.00392079f $X=0.189 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_69 N_C3_M2_g N_C1_M4_g 2.66145e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_70 N_C3_c_70_n N_Y_c_188_n 3.60572e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_71 VSS N_C3_c_70_n 0.00114532f $X=0.189 $Y=0.135 $X2=0.54 $Y2=0.0675
cc_72 N_C2_M3_g N_C1_M4_g 0.00327995f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_73 N_C2_c_84_n N_C1_c_99_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_74 N_C2_c_85_n N_C1_c_95_n 0.0046535f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_75 N_C2_M3_g N_B1_M5_g 2.71887e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_76 VSS N_C2_c_85_n 0.0011319f $X=0.243 $Y=0.135 $X2=0.54 $Y2=0.0675
cc_77 VSS N_C2_M3_g 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0.631 $Y2=0.0675
cc_78 VSS N_C2_c_85_n 0.00125352f $X=0.243 $Y=0.135 $X2=0.631 $Y2=0.0675
cc_79 VSS N_C2_c_85_n 5.07686e-19 $X=0.243 $Y=0.135 $X2=0.646 $Y2=0.0675
cc_80 N_C1_M4_g N_B1_M5_g 0.0036939f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_81 N_C1_c_99_n N_B1_c_111_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_82 N_C1_c_95_n N_B1_c_107_n 0.00406615f $X=0.297 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_83 N_C1_M4_g N_B2_M6_g 3.06651e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_84 VSS N_C1_c_95_n 0.00151583f $X=0.297 $Y=0.135 $X2=0.646 $Y2=0.0675
cc_85 N_B1_M5_g N_B2_M6_g 0.00371573f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_86 N_B1_c_111_n N_B2_c_123_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_87 N_B1_c_107_n N_B2_c_120_n 0.00483372f $X=0.351 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_88 N_B1_M5_g N_B3_M7_g 3.06651e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_89 VSS N_B1_M5_g 3.62029e-19 $X=0.351 $Y=0.0675 $X2=0.646 $Y2=0.2025
cc_90 VSS N_B1_c_107_n 0.0012322f $X=0.351 $Y=0.135 $X2=0.646 $Y2=0.2025
cc_91 N_B2_M6_g N_B3_M7_g 0.0036939f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_92 N_B2_c_123_n N_B3_c_136_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_93 N_B2_c_120_n N_B3_c_133_n 0.00483372f $X=0.405 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_94 N_B2_M6_g N_A3_M8_g 2.71887e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_95 VSS N_B2_M6_g 2.68514e-19 $X=0.405 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_96 VSS N_B2_c_120_n 0.00121543f $X=0.405 $Y=0.135 $X2=0.135 $Y2=0.135
cc_97 VSS N_B2_M6_g 2.38303e-19 $X=0.405 $Y=0.0675 $X2=0.646 $Y2=0.0675
cc_98 N_B3_M7_g N_A3_M8_g 0.00333077f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_99 N_B3_c_136_n N_A3_c_148_n 8.86777e-19 $X=0.459 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_100 N_B3_c_133_n A3 0.00406615f $X=0.459 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_101 N_B3_M7_g N_A2_M9_g 2.71887e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_102 VSS N_B3_M7_g 3.47199e-19 $X=0.459 $Y=0.0675 $X2=0.646 $Y2=0.0675
cc_103 VSS N_B3_c_133_n 5.30079e-19 $X=0.459 $Y=0.135 $X2=0.646 $Y2=0.0675
cc_104 N_A3_M8_g N_A2_M9_g 0.0036939f $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_105 N_A3_c_148_n N_A2_c_162_n 8.86777e-19 $X=0.513 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_106 A3 N_A2_c_158_n 0.00483372f $X=0.516 $Y=0.119 $X2=0.135 $Y2=0.0675
cc_107 N_A3_M8_g N_A1_M10_g 3.06651e-19 $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_108 VSS N_A3_M8_g 3.37279e-19 $X=0.513 $Y=0.0675 $X2=0.324 $Y2=0.2025
cc_109 VSS A3 5.22785e-19 $X=0.516 $Y=0.119 $X2=0.324 $Y2=0.2025
cc_110 N_A2_M9_g N_A1_M10_g 0.00376655f $X=0.567 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_111 N_A2_c_162_n N_A1_c_175_n 9.33263e-19 $X=0.567 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_112 N_A2_c_158_n N_A1_c_169_n 0.0048308f $X=0.567 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_113 VSS N_A2_M9_g 2.38303e-19 $X=0.567 $Y=0.0675 $X2=0.307 $Y2=0.2025
cc_114 VSS N_Y_c_184_n 2.23372e-19 $X=0.108 $Y=0.036 $X2=0.54 $Y2=0.0675
cc_115 VSS N_Y_c_182_n 2.83698e-19 $X=0.108 $Y=0.036 $X2=0.54 $Y2=0.0675

* END of "./OA333x2_ASAP7_75t_L.pex.sp.OA333X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OA33x2_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:51:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OA33x2_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OA33x2_ASAP7_75t_L.pex.sp.pex"
* File: OA33x2_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:51:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OA33X2_ASAP7_75T_L%3 2 7 10 13 15 17 18 21 22 25 27 28 31 33 34 35 37
+ 42 44 45 46 47 50 52 53 54 55 65 66 67 69 74 76 81 VSS
c55 82 VSS 4.63222e-19 $X=0.144 $Y=0.135
c56 81 VSS 8.47687e-19 $X=0.153 $Y=0.135
c57 76 VSS 3.28353e-19 $X=0.135 $Y=0.135
c58 74 VSS 0.00433728f $X=0.513 $Y=0.2
c59 73 VSS 0.00114071f $X=0.513 $Y=0.106
c60 72 VSS 0.0011536f $X=0.513 $Y=0.225
c61 70 VSS 4.305e-19 $X=0.477 $Y=0.072
c62 69 VSS 5.17397e-19 $X=0.468 $Y=0.072
c63 68 VSS 2.28963e-19 $X=0.45 $Y=0.072
c64 67 VSS 3.30152e-19 $X=0.446 $Y=0.072
c65 66 VSS 8.46035e-21 $X=0.414 $Y=0.072
c66 65 VSS 4.59335e-19 $X=0.396 $Y=0.072
c67 57 VSS 0.00364426f $X=0.504 $Y=0.072
c68 56 VSS 0.00338644f $X=0.486 $Y=0.234
c69 55 VSS 0.00142296f $X=0.468 $Y=0.234
c70 54 VSS 0.00344621f $X=0.45 $Y=0.234
c71 53 VSS 0.00142296f $X=0.414 $Y=0.234
c72 52 VSS 0.00291823f $X=0.396 $Y=0.234
c73 51 VSS 3.54965e-19 $X=0.364 $Y=0.234
c74 50 VSS 0.00146362f $X=0.36 $Y=0.234
c75 49 VSS 0.00274772f $X=0.342 $Y=0.234
c76 48 VSS 0.00106066f $X=0.315 $Y=0.234
c77 47 VSS 0.00142296f $X=0.306 $Y=0.234
c78 46 VSS 0.00376615f $X=0.288 $Y=0.234
c79 45 VSS 0.00142296f $X=0.252 $Y=0.234
c80 44 VSS 0.00329341f $X=0.234 $Y=0.234
c81 43 VSS 3.78291e-19 $X=0.202 $Y=0.234
c82 42 VSS 0.00146362f $X=0.198 $Y=0.234
c83 41 VSS 0.00294815f $X=0.18 $Y=0.234
c84 37 VSS 0.00270205f $X=0.162 $Y=0.234
c85 36 VSS 0.00579233f $X=0.504 $Y=0.234
c86 35 VSS 2.58269e-19 $X=0.153 $Y=0.2
c87 34 VSS 0.00132502f $X=0.153 $Y=0.189
c88 33 VSS 0.00127834f $X=0.153 $Y=0.225
c89 31 VSS 0.00218387f $X=0.324 $Y=0.2025
c90 27 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c91 25 VSS 0.0028295f $X=0.484 $Y=0.0675
c92 21 VSS 0.00244125f $X=0.378 $Y=0.0675
c93 17 VSS 5.75997e-19 $X=0.395 $Y=0.0675
c94 13 VSS 0.00419265f $X=0.135 $Y=0.135
c95 10 VSS 0.0590374f $X=0.135 $Y=0.0675
c96 2 VSS 0.06187f $X=0.081 $Y=0.0675
r97 82 83 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.1485 $Y2=0.135
r98 81 83 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.135 $X2=0.1485 $Y2=0.135
r99 76 82 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.144 $Y2=0.135
r100 73 74 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.106 $X2=0.513 $Y2=0.2
r101 72 74 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.2
r102 71 73 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.081 $X2=0.513 $Y2=0.106
r103 69 70 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.072 $X2=0.477 $Y2=0.072
r104 68 69 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.072 $X2=0.468 $Y2=0.072
r105 67 68 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.446
+ $Y=0.072 $X2=0.45 $Y2=0.072
r106 66 67 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.072 $X2=0.446 $Y2=0.072
r107 65 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.072 $X2=0.414 $Y2=0.072
r108 63 70 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.072 $X2=0.477 $Y2=0.072
r109 59 65 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.396 $Y2=0.072
r110 57 71 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.072 $X2=0.513 $Y2=0.081
r111 57 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.072 $X2=0.486 $Y2=0.072
r112 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.486 $Y2=0.234
r113 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r114 53 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.45 $Y2=0.234
r115 52 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r116 51 52 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.364
+ $Y=0.234 $X2=0.396 $Y2=0.234
r117 50 51 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.364 $Y2=0.234
r118 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r119 47 48 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.315 $Y2=0.234
r120 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r121 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.288 $Y2=0.234
r122 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r123 43 44 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.234 $X2=0.234 $Y2=0.234
r124 42 43 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.202 $Y2=0.234
r125 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r126 39 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.342 $Y2=0.234
r127 39 48 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.315 $Y2=0.234
r128 37 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r129 36 72 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.234 $X2=0.513 $Y2=0.225
r130 36 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.486 $Y2=0.234
r131 34 35 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.189 $X2=0.153 $Y2=0.2
r132 33 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.153 $Y=0.225 $X2=0.162 $Y2=0.234
r133 33 35 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.225 $X2=0.153 $Y2=0.2
r134 32 81 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.144 $X2=0.153 $Y2=0.135
r135 32 34 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.144 $X2=0.153 $Y2=0.189
r136 31 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r137 28 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r138 27 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r139 25 63 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.072
+ $X2=0.486 $Y2=0.072
r140 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.484 $Y2=0.0675
r141 21 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.072
+ $X2=0.378 $Y2=0.072
r142 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.378 $Y2=0.0675
r143 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.0675 $X2=0.378 $Y2=0.0675
r144 13 76 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r145 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r146 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r147 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r148 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r149 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OA33X2_ASAP7_75T_L%A1 2 5 7 10 13 16 VSS
c13 16 VSS 2.89025e-20 $X=0.189 $Y=0.1305
c14 13 VSS 3.18228e-19 $X=0.189 $Y=0.135
c15 10 VSS 0.00255456f $X=0.189 $Y=0.102
c16 5 VSS 0.00122965f $X=0.189 $Y=0.135
c17 2 VSS 0.0561685f $X=0.189 $Y=0.0675
r18 15 16 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.1305
r19 13 16 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.1305
r20 10 15 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.102 $X2=0.189 $Y2=0.126
r21 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OA33X2_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c13 10 VSS 0.00156318f $X=0.243 $Y=0.135
c14 5 VSS 0.00108057f $X=0.243 $Y=0.135
c15 2 VSS 0.057046f $X=0.243 $Y=0.0675
r16 10 14 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.174
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OA33X2_ASAP7_75T_L%A3 2 5 7 10 15 18 VSS
c15 18 VSS 1.57367e-19 $X=0.297 $Y=0.1205
c16 15 VSS 2.29342e-19 $X=0.297 $Y=0.135
c17 10 VSS 0.00114798f $X=0.298 $Y=0.102
c18 5 VSS 0.00110907f $X=0.297 $Y=0.135
c19 2 VSS 0.058107f $X=0.297 $Y=0.0675
r20 17 18 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.1205
r21 15 18 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.1205
r22 10 17 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.102 $X2=0.297 $Y2=0.106
r23 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r24 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r25 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OA33X2_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c13 10 VSS 5.11375e-19 $X=0.351 $Y=0.135
c14 5 VSS 0.00110628f $X=0.351 $Y=0.135
c15 2 VSS 0.0591416f $X=0.351 $Y=0.0675
r16 10 14 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.148
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OA33X2_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c12 10 VSS 4.78074e-19 $X=0.405 $Y=0.135
c13 5 VSS 0.00114557f $X=0.405 $Y=0.135
c14 2 VSS 0.0593862f $X=0.405 $Y=0.0675
r15 10 14 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.17
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OA33X2_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c9 10 VSS 7.06488e-19 $X=0.459 $Y=0.135
c10 5 VSS 0.00171018f $X=0.459 $Y=0.135
c11 2 VSS 0.0629181f $X=0.459 $Y=0.0675
r12 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.154
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OA33X2_ASAP7_75T_L%Y 1 2 6 7 10 14 16 18 19 23 24 26 30 39 VSS
c18 39 VSS 0.00143505f $X=0.108 $Y=0.216
c19 33 VSS 0.00229462f $X=0.0805 $Y=0.234
c20 32 VSS 0.00605721f $X=0.062 $Y=0.234
c21 31 VSS 0.00319807f $X=0.027 $Y=0.234
c22 30 VSS 0.00368818f $X=0.099 $Y=0.234
c23 26 VSS 0.00277019f $X=0.085 $Y=0.036
c24 25 VSS 0.00605721f $X=0.062 $Y=0.036
c25 24 VSS 0.00902111f $X=0.108 $Y=0.036
c26 23 VSS 0.00424555f $X=0.108 $Y=0.036
c27 21 VSS 0.00320021f $X=0.027 $Y=0.036
c28 20 VSS 7.68735e-19 $X=0.018 $Y=0.207
c29 19 VSS 0.00246086f $X=0.018 $Y=0.189
c30 18 VSS 8.11473e-19 $X=0.018 $Y=0.144
c31 16 VSS 8.76885e-19 $X=0.018 $Y=0.086
c32 15 VSS 0.00126561f $X=0.018 $Y=0.07
c33 14 VSS 0.00227807f $X=0.02 $Y=0.102
c34 12 VSS 6.2588e-19 $X=0.018 $Y=0.225
c35 10 VSS 0.0105087f $X=0.108 $Y=0.2025
c36 6 VSS 5.945e-19 $X=0.125 $Y=0.2025
c37 1 VSS 5.58795e-19 $X=0.125 $Y=0.0675
r38 37 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.225 $X2=0.108 $Y2=0.216
r39 32 33 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.062
+ $Y=0.234 $X2=0.0805 $Y2=0.234
r40 31 32 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.062 $Y2=0.234
r41 30 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.099 $Y=0.234 $X2=0.108 $Y2=0.225
r42 30 33 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.234 $X2=0.0805 $Y2=0.234
r43 25 26 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.062
+ $Y=0.036 $X2=0.085 $Y2=0.036
r44 23 26 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.085 $Y2=0.036
r45 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r46 21 25 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.062 $Y2=0.036
r47 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.207
r48 18 19 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.189
r49 17 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.144
r50 15 16 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.086
r51 14 17 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.102 $X2=0.018 $Y2=0.126
r52 14 16 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.102 $X2=0.018 $Y2=0.086
r53 12 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r54 12 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.207
r55 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r56 11 15 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r57 10 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.216 $X2=0.108
+ $Y2=0.216
r58 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r59 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r60 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r61 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r62 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OA33x2_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OA33x2_ASAP7_75t_L  VSS VDD A1 A2 A3 B3 B2 B1 Y
* 
* Y	Y
* B1	B1
* B2	B2
* B3	B3
* A3	A3
* A2	A2
* A1	A1
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_11 N_A1_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_A2_M3_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_11 N_A3_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 N_3_M5_d N_B3_M5_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_11 N_B2_M6_g N_3_M6_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_3_M7_d N_B1_M7_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_Y_M8_d N_3_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M9 N_Y_M9_d N_3_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M10 noxref_12 N_A1_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M11 noxref_13 N_A2_M11_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M12 N_3_M12_d N_A3_M12_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M13 noxref_14 N_B3_M13_g N_3_M13_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M14 noxref_15 N_B2_M14_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M15 VDD N_B1_M15_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "OA33x2_ASAP7_75t_L.pex.sp.OA33X2_ASAP7_75T_L.pxi"
* BEGIN of "./OA33x2_ASAP7_75t_L.pex.sp.OA33X2_ASAP7_75T_L.pxi"
* File: OA33x2_ASAP7_75t_L.pex.sp.OA33X2_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:51:48 2017
* 
x_PM_OA33X2_ASAP7_75T_L%3 N_3_M0_g N_3_M8_g N_3_M1_g N_3_c_4_p N_3_M9_g N_3_M6_s
+ N_3_M5_d N_3_c_42_p N_3_M7_d N_3_c_45_p N_3_M13_s N_3_M12_d N_3_c_13_p
+ N_3_c_40_p N_3_c_5_p N_3_c_41_p N_3_c_37_p N_3_c_3_p N_3_c_52_p N_3_c_9_p
+ N_3_c_53_p N_3_c_11_p N_3_c_15_p N_3_c_54_p N_3_c_18_p N_3_c_55_p N_3_c_22_p
+ N_3_c_12_p N_3_c_19_p N_3_c_49_p N_3_c_23_p N_3_c_26_p N_3_c_32_p N_3_c_7_p
+ VSS PM_OA33X2_ASAP7_75T_L%3
x_PM_OA33X2_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_59_n N_A1_M10_g A1 N_A1_c_60_n
+ N_A1_c_62_n VSS PM_OA33X2_ASAP7_75T_L%A1
x_PM_OA33X2_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_73_n N_A2_M11_g N_A2_c_71_n A2 VSS
+ PM_OA33X2_ASAP7_75T_L%A2
x_PM_OA33X2_ASAP7_75T_L%A3 N_A3_M4_g N_A3_c_88_n N_A3_M12_g A3 N_A3_c_84_n
+ N_A3_c_92_p VSS PM_OA33X2_ASAP7_75T_L%A3
x_PM_OA33X2_ASAP7_75T_L%B3 N_B3_M5_g N_B3_c_102_n N_B3_M13_g N_B3_c_98_n B3 VSS
+ PM_OA33X2_ASAP7_75T_L%B3
x_PM_OA33X2_ASAP7_75T_L%B2 N_B2_M6_g N_B2_c_116_n N_B2_M14_g N_B2_c_112_n B2 VSS
+ PM_OA33X2_ASAP7_75T_L%B2
x_PM_OA33X2_ASAP7_75T_L%B1 N_B1_M7_g N_B1_c_129_n N_B1_M15_g N_B1_c_124_n B1 VSS
+ PM_OA33X2_ASAP7_75T_L%B1
x_PM_OA33X2_ASAP7_75T_L%Y N_Y_M1_d N_Y_M0_d N_Y_M9_d N_Y_M8_d N_Y_c_133_n Y
+ N_Y_c_146_n N_Y_c_136_n N_Y_c_137_n N_Y_c_148_p N_Y_c_138_n N_Y_c_139_n
+ N_Y_c_141_n N_Y_c_142_n VSS PM_OA33X2_ASAP7_75T_L%Y
cc_1 N_3_M0_g N_A1_M2_g 2.13359e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_A1_M2_g 0.00268443f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_A1_M2_g 2.64276e-19 $X=0.198 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_4 N_3_c_4_p N_A1_c_59_n 0.00111954f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_5 N_3_c_5_p N_A1_c_60_n 0.0030573f $X=0.153 $Y=0.189 $X2=0.189 $Y2=0.135
cc_6 N_3_c_3_p N_A1_c_60_n 0.00125352f $X=0.198 $Y=0.234 $X2=0.189 $Y2=0.135
cc_7 N_3_c_7_p N_A1_c_62_n 0.0030573f $X=0.153 $Y=0.135 $X2=0.189 $Y2=0.1305
cc_8 N_3_M1_g N_A2_M3_g 2.13359e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_9 N_3_c_9_p N_A2_M3_g 3.38929e-19 $X=0.252 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_10 N_3_c_9_p N_A2_c_71_n 0.00123604f $X=0.252 $Y=0.234 $X2=0.189 $Y2=0.102
cc_11 N_3_c_11_p N_A3_M4_g 2.56935e-19 $X=0.306 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_12 N_3_c_12_p A3 2.64308e-19 $X=0.396 $Y=0.072 $X2=0.189 $Y2=0.102
cc_13 N_3_c_13_p N_A3_c_84_n 0.0013295f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.126
cc_14 N_3_c_11_p N_A3_c_84_n 0.00123604f $X=0.306 $Y=0.234 $X2=0.189 $Y2=0.126
cc_15 N_3_c_15_p N_B3_M5_g 2.64276e-19 $X=0.36 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_16 N_3_c_13_p N_B3_c_98_n 0.0013295f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.102
cc_17 N_3_c_15_p N_B3_c_98_n 0.00124805f $X=0.36 $Y=0.234 $X2=0.189 $Y2=0.102
cc_18 N_3_c_18_p N_B2_M6_g 3.38929e-19 $X=0.414 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_19 N_3_c_19_p N_B2_M6_g 2.76185e-19 $X=0.414 $Y=0.072 $X2=0.189 $Y2=0.0675
cc_20 N_3_c_18_p N_B2_c_112_n 0.00123064f $X=0.414 $Y=0.234 $X2=0.189 $Y2=0.102
cc_21 N_3_c_19_p N_B2_c_112_n 0.0012322f $X=0.414 $Y=0.072 $X2=0.189 $Y2=0.102
cc_22 N_3_c_22_p N_B1_M7_g 2.56935e-19 $X=0.468 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_23 N_3_c_23_p N_B1_M7_g 3.51973e-19 $X=0.468 $Y=0.072 $X2=0.189 $Y2=0.0675
cc_24 N_3_c_22_p N_B1_c_124_n 0.00123064f $X=0.468 $Y=0.234 $X2=0.189 $Y2=0.102
cc_25 N_3_c_23_p N_B1_c_124_n 0.00121543f $X=0.468 $Y=0.072 $X2=0.189 $Y2=0.102
cc_26 N_3_c_26_p N_B1_c_124_n 0.00392202f $X=0.513 $Y=0.2 $X2=0.189 $Y2=0.102
cc_27 N_3_c_4_p N_Y_M1_d 3.80485e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_28 N_3_c_4_p N_Y_M9_d 3.80277e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_29 N_3_c_4_p N_Y_c_133_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.102
cc_30 N_3_c_5_p N_Y_c_133_n 0.00142255f $X=0.153 $Y=0.189 $X2=0.189 $Y2=0.102
cc_31 N_3_c_4_p Y 4.11298e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_32 N_3_c_32_p N_Y_c_136_n 2.07283e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_33 N_3_c_5_p N_Y_c_137_n 3.92722e-19 $X=0.153 $Y=0.189 $X2=0 $Y2=0
cc_34 N_3_c_4_p N_Y_c_138_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_35 N_3_M0_g N_Y_c_139_n 3.21831e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_3_c_4_p N_Y_c_139_n 5.00341e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_37 N_3_c_37_p N_Y_c_141_n 0.00111507f $X=0.162 $Y=0.234 $X2=0 $Y2=0
cc_38 N_3_M0_g N_Y_c_142_n 3.68592e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_3_c_4_p N_Y_c_142_n 7.28855e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_40 N_3_c_40_p N_Y_c_142_n 0.00111507f $X=0.153 $Y=0.225 $X2=0 $Y2=0
cc_41 N_3_c_41_p N_Y_c_142_n 0.00111507f $X=0.153 $Y=0.2 $X2=0 $Y2=0
cc_42 VSS N_3_c_42_p 0.00364243f $X=0.378 $Y=0.0675 $X2=0 $Y2=0
cc_43 VSS N_3_c_13_p 0.00107252f $X=0.324 $Y=0.2025 $X2=0 $Y2=0
cc_44 VSS N_3_c_12_p 3.61571e-19 $X=0.396 $Y=0.072 $X2=0 $Y2=0
cc_45 VSS N_3_c_45_p 3.09693e-19 $X=0.484 $Y=0.0675 $X2=0 $Y2=0
cc_46 VSS N_3_c_19_p 0.00351217f $X=0.414 $Y=0.072 $X2=0 $Y2=0
cc_47 VSS N_3_c_42_p 0.0035539f $X=0.378 $Y=0.0675 $X2=0 $Y2=0
cc_48 VSS N_3_c_45_p 0.00339796f $X=0.484 $Y=0.0675 $X2=0 $Y2=0
cc_49 VSS N_3_c_49_p 0.00233206f $X=0.446 $Y=0.072 $X2=0 $Y2=0
cc_50 VSS N_3_c_42_p 0.00250965f $X=0.378 $Y=0.0675 $X2=0 $Y2=0
cc_51 VSS N_3_c_12_p 0.00351217f $X=0.396 $Y=0.072 $X2=0 $Y2=0
cc_52 VSS N_3_c_52_p 3.25855e-19 $X=0.234 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_53 VSS N_3_c_53_p 3.56327e-19 $X=0.288 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_54 VSS N_3_c_54_p 3.19955e-19 $X=0.396 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_55 VSS N_3_c_55_p 3.48201e-19 $X=0.45 $Y=0.234 $X2=0.189 $Y2=0.0675
cc_56 N_A1_M2_g N_A2_M3_g 0.00328721f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_57 N_A1_c_59_n N_A2_c_73_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_58 A1 N_A2_c_71_n 0.00582194f $X=0.189 $Y=0.102 $X2=0.135 $Y2=0.0675
cc_59 N_A1_M2_g N_A3_M4_g 2.48122e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_60 A1 N_Y_c_146_n 2.87432e-19 $X=0.189 $Y=0.102 $X2=0 $Y2=0
cc_61 VSS A1 0.00114532f $X=0.189 $Y=0.102 $X2=0.361 $Y2=0.0675
cc_62 N_A2_M3_g N_A3_M4_g 0.00312021f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_63 N_A2_c_73_n N_A3_c_88_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_64 N_A2_c_71_n A3 0.00581002f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_65 N_A2_M3_g N_B3_M5_g 2.53865e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_66 VSS N_A2_c_71_n 0.00114532f $X=0.243 $Y=0.135 $X2=0.361 $Y2=0.0675
cc_67 VSS N_A2_M3_g 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_68 VSS N_A2_c_71_n 0.00125352f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_69 N_A3_M4_g N_B3_M5_g 0.00353416f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_70 N_A3_c_88_n N_B3_c_102_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_71 N_A3_c_92_p N_B3_c_98_n 0.00389526f $X=0.297 $Y=0.1205 $X2=0.135
+ $Y2=0.0675
cc_72 N_A3_M4_g N_B2_M6_g 2.88628e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_73 VSS A3 9.86946e-19 $X=0.298 $Y=0.102 $X2=0.469 $Y2=0.0675
cc_74 VSS N_A3_M4_g 2.64276e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_75 VSS A3 0.00125352f $X=0.298 $Y=0.102 $X2=0 $Y2=0
cc_76 N_B3_M5_g N_B2_M6_g 0.00355599f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_77 N_B3_c_102_n N_B2_c_116_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_78 N_B3_c_98_n N_B2_c_112_n 0.00483372f $X=0.351 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_79 N_B3_M5_g N_B1_M7_g 2.88628e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_80 VSS N_B3_M5_g 3.57119e-19 $X=0.351 $Y=0.0675 $X2=0.324 $Y2=0.2025
cc_81 VSS N_B3_c_98_n 5.37372e-19 $X=0.351 $Y=0.135 $X2=0.324 $Y2=0.2025
cc_82 N_B2_M6_g N_B1_M7_g 0.00353416f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_83 N_B2_c_116_n N_B1_c_129_n 9.33263e-19 $X=0.405 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_84 N_B2_c_112_n N_B1_c_124_n 0.0048308f $X=0.405 $Y=0.135 $X2=0.135
+ $Y2=0.0675
cc_85 VSS N_B2_M6_g 2.08515e-19 $X=0.405 $Y=0.0675 $X2=0.307 $Y2=0.2025
cc_86 VSS N_Y_c_138_n 2.23372e-19 $X=0.108 $Y=0.036 $X2=0.361 $Y2=0.0675
cc_87 VSS N_Y_c_148_p 2.92912e-19 $X=0.108 $Y=0.036 $X2=0.484 $Y2=0.0675

* END of "./OA33x2_ASAP7_75t_L.pex.sp.OA33X2_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI211xp5_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:52:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI211xp5_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI211xp5_ASAP7_75t_L.pex.sp.pex"
* File: OAI211xp5_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:52:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI211XP5_ASAP7_75T_L%A2 2 5 7 11 16 21 24 26 VSS
c12 26 VSS 0.00462465f $X=0.027 $Y=0.135
c13 24 VSS 4.81186e-19 $X=0.0605 $Y=0.135
c14 23 VSS 5.77998e-19 $X=0.04 $Y=0.135
c15 21 VSS 2.24273e-19 $X=0.081 $Y=0.135
c16 16 VSS 5.19709e-19 $X=0.027 $Y=0.116
c17 11 VSS 0.00256757f $X=0.023 $Y=0.083
c18 9 VSS 4.97319e-19 $X=0.027 $Y=0.126
c19 5 VSS 0.00258107f $X=0.081 $Y=0.135
c20 2 VSS 0.0662757f $X=0.081 $Y=0.0675
r21 23 24 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.135 $X2=0.0605 $Y2=0.135
r22 21 24 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0605 $Y2=0.135
r23 19 26 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.135 $X2=0.027 $Y2=0.135
r24 19 23 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.135 $X2=0.04 $Y2=0.135
r25 15 16 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.106 $X2=0.027 $Y2=0.116
r26 11 15 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.083 $X2=0.027 $Y2=0.106
r27 9 26 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.126 $X2=0.027 $Y2=0.135
r28 9 16 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.126 $X2=0.027 $Y2=0.116
r29 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r30 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r31 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI211XP5_ASAP7_75T_L%A1 2 5 7 10 16 18 VSS
c14 18 VSS 1.73756e-19 $X=0.135 $Y=0.1655
c15 16 VSS 7.88062e-19 $X=0.134 $Y=0.187
c16 10 VSS 4.56151e-19 $X=0.135 $Y=0.135
c17 5 VSS 0.00117984f $X=0.135 $Y=0.135
c18 2 VSS 0.0602081f $X=0.135 $Y=0.0675
r19 17 18 1.45988 $w=1.8e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.1655
r20 16 18 1.45988 $w=1.8e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.187 $X2=0.135 $Y2=0.1655
r21 10 17 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r22 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r23 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r24 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI211XP5_ASAP7_75T_L%B 2 5 7 10 14 VSS
c12 10 VSS 9.85944e-19 $X=0.189 $Y=0.135
c13 5 VSS 0.00116143f $X=0.189 $Y=0.135
c14 2 VSS 0.059171f $X=0.189 $Y=0.0675
r15 10 14 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.148
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI211XP5_ASAP7_75T_L%C 2 5 7 10 VSS
c10 10 VSS 9.75038e-19 $X=0.241 $Y=0.123
c11 5 VSS 0.00172166f $X=0.243 $Y=0.135
c12 2 VSS 0.0618315f $X=0.243 $Y=0.0675
r13 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.123 $X2=0.243 $Y2=0.135
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI211XP5_ASAP7_75T_L%Y 1 2 5 6 9 11 12 15 24 27 29 31 37 38 39 41 42
+ 43 48 50 VSS
c26 52 VSS 7.14098e-19 $X=0.297 $Y=0.2125
c27 50 VSS 0.00150919f $X=0.297 $Y=0.139
c28 49 VSS 0.00131846f $X=0.297 $Y=0.106
c29 48 VSS 0.0027951f $X=0.299 $Y=0.172
c30 46 VSS 6.07272e-19 $X=0.297 $Y=0.225
c31 44 VSS 0.00236172f $X=0.27 $Y=0.072
c32 43 VSS 5.17397e-19 $X=0.252 $Y=0.072
c33 42 VSS 0.00175846f $X=0.234 $Y=0.072
c34 41 VSS 5.17397e-19 $X=0.198 $Y=0.072
c35 40 VSS 2.28963e-19 $X=0.18 $Y=0.072
c36 39 VSS 4.67884e-19 $X=0.176 $Y=0.072
c37 38 VSS 8.46035e-21 $X=0.144 $Y=0.072
c38 37 VSS 7.15352e-19 $X=0.126 $Y=0.072
c39 32 VSS 0.00390806f $X=0.288 $Y=0.072
c40 31 VSS 0.00146362f $X=0.252 $Y=0.234
c41 30 VSS 0.00346254f $X=0.234 $Y=0.234
c42 29 VSS 0.00146362f $X=0.198 $Y=0.234
c43 28 VSS 0.00577782f $X=0.18 $Y=0.234
c44 27 VSS 0.00146362f $X=0.144 $Y=0.234
c45 26 VSS 0.00257933f $X=0.126 $Y=0.234
c46 25 VSS 9.06382e-19 $X=0.099 $Y=0.234
c47 24 VSS 0.00532554f $X=0.09 $Y=0.234
c48 16 VSS 0.00884695f $X=0.288 $Y=0.234
c49 15 VSS 0.00790803f $X=0.216 $Y=0.216
c50 11 VSS 5.3314e-19 $X=0.233 $Y=0.216
c51 9 VSS 0.00348545f $X=0.056 $Y=0.216
c52 6 VSS 2.6657e-19 $X=0.071 $Y=0.216
c53 5 VSS 0.00210856f $X=0.108 $Y=0.0675
c54 1 VSS 6.64001e-19 $X=0.125 $Y=0.0675
r55 51 52 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.2 $X2=0.297 $Y2=0.2125
r56 49 50 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.139
r57 48 51 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.172 $X2=0.297 $Y2=0.2
r58 48 50 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.172 $X2=0.297 $Y2=0.139
r59 46 52 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.2125
r60 45 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.081 $X2=0.297 $Y2=0.106
r61 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.072 $X2=0.27 $Y2=0.072
r62 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.252 $Y2=0.072
r63 41 42 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.072 $X2=0.234 $Y2=0.072
r64 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.072 $X2=0.198 $Y2=0.072
r65 39 40 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.072 $X2=0.18 $Y2=0.072
r66 38 39 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.176 $Y2=0.072
r67 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.144 $Y2=0.072
r68 34 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.126 $Y2=0.072
r69 32 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.072 $X2=0.297 $Y2=0.081
r70 32 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.27 $Y2=0.072
r71 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r72 28 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r73 27 28 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.18 $Y2=0.234
r74 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r75 25 26 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.234 $X2=0.126 $Y2=0.234
r76 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.099 $Y2=0.234
r77 22 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.234 $Y2=0.234
r78 22 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.198 $Y2=0.234
r79 18 24 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.09 $Y2=0.234
r80 16 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.234 $X2=0.297 $Y2=0.225
r81 16 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.252 $Y2=0.234
r82 15 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r83 12 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.216 $X2=0.216 $Y2=0.216
r84 11 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.216 $X2=0.216 $Y2=0.216
r85 9 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r86 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.216 $X2=0.056 $Y2=0.216
r87 5 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072 $X2=0.108
+ $Y2=0.072
r88 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r89 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OAI211xp5_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI211xp5_ASAP7_75t_L  VSS VDD A2 A1 B C Y
* 
* Y	Y
* C	C
* B	B
* A1	A1
* A2	A2
M0 N_Y_M0_d N_A2_M0_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_7 N_A1_M1_g N_Y_M1_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_9 N_B_M2_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_C_M3_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 noxref_10 N_A2_M4_g N_Y_M4_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M5 VDD N_A1_M5_g noxref_10 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M6 N_Y_M6_d N_B_M6_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.189
M7 VDD N_C_M7_g N_Y_M7_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.189
*
* 
* .include "OAI211xp5_ASAP7_75t_L.pex.sp.OAI211XP5_ASAP7_75T_L.pxi"
* BEGIN of "./OAI211xp5_ASAP7_75t_L.pex.sp.OAI211XP5_ASAP7_75T_L.pxi"
* File: OAI211xp5_ASAP7_75t_L.pex.sp.OAI211XP5_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:52:11 2017
* 
x_PM_OAI211XP5_ASAP7_75T_L%A2 N_A2_M0_g N_A2_c_2_p N_A2_M4_g A2 N_A2_c_3_p
+ N_A2_c_4_p N_A2_c_9_p N_A2_c_5_p VSS PM_OAI211XP5_ASAP7_75T_L%A2
x_PM_OAI211XP5_ASAP7_75T_L%A1 N_A1_M1_g N_A1_c_14_n N_A1_M5_g N_A1_c_15_n A1
+ N_A1_c_17_n VSS PM_OAI211XP5_ASAP7_75T_L%A1
x_PM_OAI211XP5_ASAP7_75T_L%B N_B_M2_g N_B_c_29_n N_B_M6_g N_B_c_30_n B VSS
+ PM_OAI211XP5_ASAP7_75T_L%B
x_PM_OAI211XP5_ASAP7_75T_L%C N_C_M3_g N_C_c_41_n N_C_M7_g C VSS
+ PM_OAI211XP5_ASAP7_75T_L%C
x_PM_OAI211XP5_ASAP7_75T_L%Y N_Y_M1_s N_Y_M0_d N_Y_c_67_n N_Y_M4_s N_Y_c_49_n
+ N_Y_M7_s N_Y_M6_d N_Y_c_56_n N_Y_c_50_n N_Y_c_52_n N_Y_c_57_n N_Y_c_62_n
+ N_Y_c_72_n N_Y_c_54_n N_Y_c_73_n N_Y_c_59_n N_Y_c_74_p N_Y_c_64_n Y N_Y_c_66_n
+ VSS PM_OAI211XP5_ASAP7_75T_L%Y
cc_1 N_A2_M0_g N_A1_M1_g 0.00364065f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A2_c_2_p N_A1_c_14_n 9.83624e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A2_c_3_p N_A1_c_15_n 4.14444e-19 $X=0.027 $Y=0.116 $X2=0.135 $Y2=0.135
cc_4 N_A2_c_4_p N_A1_c_15_n 6.03818e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_5 N_A2_c_5_p N_A1_c_17_n 0.00108013f $X=0.027 $Y=0.135 $X2=0.135 $Y2=0.1655
cc_6 N_A2_M0_g N_B_M2_g 2.6588e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_7 VSS A2 0.00163906f $X=0.023 $Y=0.083 $X2=0 $Y2=0
cc_8 VSS N_A2_M0_g 4.01862e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.1655
cc_9 VSS N_A2_c_9_p 9.66105e-19 $X=0.0605 $Y=0.135 $X2=0.135 $Y2=0.1655
cc_10 N_A2_c_5_p N_Y_c_49_n 3.85925e-19 $X=0.027 $Y=0.135 $X2=0.135 $Y2=0.135
cc_11 N_A2_M0_g N_Y_c_50_n 4.01862e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_12 N_A2_c_9_p N_Y_c_50_n 9.13307e-19 $X=0.0605 $Y=0.135 $X2=0 $Y2=0
cc_13 N_A1_M1_g N_B_M2_g 0.0032267f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_A1_c_14_n N_B_c_29_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 N_A1_c_15_n N_B_c_30_n 0.00454568f $X=0.135 $Y=0.135 $X2=0.027 $Y2=0.083
cc_16 N_A1_M1_g N_C_M3_g 2.60137e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 VSS N_A1_M1_g 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0.027 $Y2=0.116
cc_18 N_A1_M1_g N_Y_c_52_n 2.64276e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 A1 N_Y_c_52_n 0.00124805f $X=0.134 $Y=0.187 $X2=0 $Y2=0
cc_20 N_A1_M1_g N_Y_c_54_n 2.76185e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_21 N_A1_c_15_n N_Y_c_54_n 0.0012322f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_22 N_B_M2_g N_C_M3_g 0.0033937f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_23 N_B_c_29_n N_C_c_41_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_B_c_30_n C 0.0046131f $X=0.189 $Y=0.135 $X2=0.027 $Y2=0.083
cc_25 N_B_c_30_n N_Y_c_56_n 3.31541e-19 $X=0.189 $Y=0.135 $X2=0.027 $Y2=0.106
cc_26 N_B_M2_g N_Y_c_57_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_B_c_30_n N_Y_c_57_n 0.00124805f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_28 N_B_M2_g N_Y_c_59_n 3.51973e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_29 N_B_c_30_n N_Y_c_59_n 0.00121543f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_30 C N_Y_c_56_n 3.31541e-19 $X=0.241 $Y=0.123 $X2=0.135 $Y2=0.187
cc_31 N_C_M3_g N_Y_c_62_n 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_32 C N_Y_c_62_n 0.00124805f $X=0.241 $Y=0.123 $X2=0 $Y2=0
cc_33 N_C_M3_g N_Y_c_64_n 3.51973e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_34 C N_Y_c_64_n 0.00121543f $X=0.241 $Y=0.123 $X2=0 $Y2=0
cc_35 C N_Y_c_66_n 0.00440946f $X=0.241 $Y=0.123 $X2=0 $Y2=0
cc_36 VSS N_Y_c_67_n 0.0036868f $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.135
cc_37 VSS N_Y_c_67_n 0.00189275f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_38 VSS N_Y_c_67_n 0.00359726f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_39 VSS N_Y_c_67_n 6.35113e-19 $X=0.099 $Y=0.036 $X2=0.081 $Y2=0.135
cc_40 VSS N_Y_c_49_n 8.7738e-19 $X=0.054 $Y=0.036 $X2=0.027 $Y2=0.126
cc_41 VSS N_Y_c_72_n 0.00666759f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_42 VSS N_Y_c_73_n 0.00262229f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_43 VSS N_Y_c_74_p 4.30621e-19 $X=0.234 $Y=0.072 $X2=0.081 $Y2=0.0675

* END of "./OAI211xp5_ASAP7_75t_L.pex.sp.OAI211XP5_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI21x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:52:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI21x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI21x1_ASAP7_75t_L.pex.sp.pex"
* File: OAI21x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:52:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI21X1_ASAP7_75T_L%B 2 5 7 10 13 15 19 20 21 25 26 28 29 30 31 32 33
+ 34 35 36 39 41 42 VSS
c38 42 VSS 1.30627e-19 $X=0.351 $Y=0.119
c39 39 VSS 2.04795e-19 $X=0.351 $Y=0.136
c40 36 VSS 1.62028e-19 $X=0.3375 $Y=0.072
c41 35 VSS 2.77255e-19 $X=0.333 $Y=0.072
c42 34 VSS 7.99121e-21 $X=0.306 $Y=0.072
c43 33 VSS 0.00327176f $X=0.288 $Y=0.072
c44 32 VSS 2.08366e-19 $X=0.256 $Y=0.072
c45 31 VSS 1.73836e-19 $X=0.227 $Y=0.072
c46 30 VSS 0.0016554f $X=0.19 $Y=0.072
c47 29 VSS 0.00126552f $X=0.163 $Y=0.072
c48 28 VSS 4.27363e-19 $X=0.126 $Y=0.072
c49 27 VSS 5.57344e-19 $X=0.099 $Y=0.072
c50 26 VSS 8.76255e-19 $X=0.09 $Y=0.072
c51 25 VSS 0.00103635f $X=0.342 $Y=0.072
c52 21 VSS 7.55716e-20 $X=0.081 $Y=0.11725
c53 19 VSS 0.00142772f $X=0.0835 $Y=0.1355
c54 13 VSS 0.00242651f $X=0.351 $Y=0.135
c55 10 VSS 0.0654437f $X=0.351 $Y=0.0675
c56 5 VSS 0.00246842f $X=0.081 $Y=0.135
c57 2 VSS 0.0651019f $X=0.081 $Y=0.0675
r58 41 42 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.099 $X2=0.351 $Y2=0.119
r59 39 42 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.136 $X2=0.351 $Y2=0.119
r60 37 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.099
r61 35 36 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.072 $X2=0.3375 $Y2=0.072
r62 34 35 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.072 $X2=0.333 $Y2=0.072
r63 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.306 $Y2=0.072
r64 32 33 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.072 $X2=0.288 $Y2=0.072
r65 31 32 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.227
+ $Y=0.072 $X2=0.256 $Y2=0.072
r66 30 31 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.19
+ $Y=0.072 $X2=0.227 $Y2=0.072
r67 29 30 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.163
+ $Y=0.072 $X2=0.19 $Y2=0.072
r68 28 29 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.163 $Y2=0.072
r69 27 28 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.072 $X2=0.126 $Y2=0.072
r70 26 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.099 $Y2=0.072
r71 25 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.072 $X2=0.351 $Y2=0.081
r72 25 36 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.072 $X2=0.3375 $Y2=0.072
r73 20 21 1.2392 $w=1.8e-08 $l=1.825e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.099 $X2=0.081 $Y2=0.11725
r74 19 21 1.2392 $w=1.8e-08 $l=1.825e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.1355 $X2=0.081 $Y2=0.11725
r75 17 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.081 $X2=0.09 $Y2=0.072
r76 17 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.081 $X2=0.081 $Y2=0.099
r77 13 39 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.136 $X2=0.351
+ $Y2=0.136
r78 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r79 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r80 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.136 $X2=0.081
+ $Y2=0.136
r81 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r82 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI21X1_ASAP7_75T_L%A1 2 5 7 10 13 15 20 24 25 26 27 28 29 30 33 39
+ 40 VSS
c36 41 VSS 1.80714e-19 $X=0.297 $Y=0.18
c37 40 VSS 1.83154e-19 $X=0.297 $Y=0.171
c38 39 VSS 3.74688e-20 $X=0.297 $Y=0.154
c39 33 VSS 1.56099e-19 $X=0.297 $Y=0.136
c40 31 VSS 1.70674e-19 $X=0.297 $Y=0.189
c41 30 VSS 9.36428e-19 $X=0.256 $Y=0.198
c42 29 VSS 0.00235496f $X=0.227 $Y=0.198
c43 28 VSS 6.28049e-19 $X=0.19 $Y=0.198
c44 27 VSS 1.08538e-19 $X=0.163 $Y=0.198
c45 26 VSS 1.13858e-19 $X=0.144 $Y=0.198
c46 25 VSS 3.61504e-19 $X=0.288 $Y=0.198
c47 24 VSS 1.80714e-19 $X=0.135 $Y=0.18
c48 20 VSS 0.00167247f $X=0.1345 $Y=0.1355
c49 18 VSS 1.70674e-19 $X=0.135 $Y=0.189
c50 13 VSS 0.00167162f $X=0.297 $Y=0.135
c51 10 VSS 0.0606704f $X=0.297 $Y=0.0675
c52 5 VSS 0.00154002f $X=0.135 $Y=0.135
c53 2 VSS 0.0604995f $X=0.135 $Y=0.0675
r54 40 41 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.171 $X2=0.297 $Y2=0.18
r55 39 40 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.154 $X2=0.297 $Y2=0.171
r56 38 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.145 $X2=0.297 $Y2=0.154
r57 33 38 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.136 $X2=0.297 $Y2=0.145
r58 31 41 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.18
r59 29 30 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.227
+ $Y=0.198 $X2=0.256 $Y2=0.198
r60 28 29 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.19
+ $Y=0.198 $X2=0.227 $Y2=0.198
r61 27 28 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.163
+ $Y=0.198 $X2=0.19 $Y2=0.198
r62 26 27 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.198 $X2=0.163 $Y2=0.198
r63 25 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.198 $X2=0.297 $Y2=0.189
r64 25 30 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.256 $Y2=0.198
r65 23 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.171 $X2=0.135 $Y2=0.18
r66 20 23 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.171
r67 18 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.189 $X2=0.144 $Y2=0.198
r68 18 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.135 $Y2=0.18
r69 13 33 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.136 $X2=0.297
+ $Y2=0.136
r70 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r71 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r72 5 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.136 $X2=0.135
+ $Y2=0.136
r73 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r74 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI21X1_ASAP7_75T_L%A2 2 7 10 13 15 18 VSS
c27 18 VSS 0.00293381f $X=0.2085 $Y=0.1355
c28 13 VSS 0.00737317f $X=0.243 $Y=0.135
c29 10 VSS 0.0624282f $X=0.243 $Y=0.0675
c30 2 VSS 0.0626776f $X=0.189 $Y=0.0675
r31 18 20 0.797927 $w=4.825e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2085 $Y=0.135 $X2=0.24 $Y2=0.135
r32 13 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.24 $Y=0.136 $X2=0.24
+ $Y2=0.136
r33 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r34 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r35 5 13 46.3636 $w=2.2e-08 $l=5.1e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.24 $Y2=0.135
r36 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r37 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI21X1_ASAP7_75T_L%Y 1 6 11 12 15 16 17 20 24 26 36 42 44 50 51 56
+ 57 63 66 VSS
c26 66 VSS 0.00362882f $X=0.396 $Y=0.036
c27 65 VSS 0.00277971f $X=0.405 $Y=0.036
c28 63 VSS 0.00401496f $X=0.378 $Y=0.036
c29 59 VSS 0.00100946f $X=0.045 $Y=0.036
c30 58 VSS 0.00328948f $X=0.036 $Y=0.036
c31 57 VSS 0.00401379f $X=0.054 $Y=0.036
c32 56 VSS 0.00253697f $X=0.054 $Y=0.036
c33 52 VSS 5.60269e-19 $X=0.405 $Y=0.216
c34 51 VSS 0.00286958f $X=0.405 $Y=0.207
c35 50 VSS 0.00389061f $X=0.405 $Y=0.154
c36 49 VSS 0.00102822f $X=0.405 $Y=0.063
c37 48 VSS 5.29143e-19 $X=0.405 $Y=0.225
c38 46 VSS 0.00208805f $X=0.3825 $Y=0.234
c39 45 VSS 0.0014903f $X=0.369 $Y=0.234
c40 44 VSS 0.00146498f $X=0.36 $Y=0.234
c41 43 VSS 0.00372523f $X=0.342 $Y=0.234
c42 42 VSS 0.0175638f $X=0.306 $Y=0.234
c43 41 VSS 0.00273151f $X=0.126 $Y=0.234
c44 37 VSS 9.61644e-19 $X=0.099 $Y=0.234
c45 36 VSS 0.00142432f $X=0.09 $Y=0.234
c46 35 VSS 0.00155038f $X=0.072 $Y=0.234
c47 34 VSS 0.00383968f $X=0.063 $Y=0.234
c48 30 VSS 0.00340653f $X=0.036 $Y=0.234
c49 29 VSS 0.00521081f $X=0.396 $Y=0.234
c50 28 VSS 3.99179e-19 $X=0.027 $Y=0.207
c51 26 VSS 9.21872e-19 $X=0.027 $Y=0.087
c52 25 VSS 5.7946e-19 $X=0.027 $Y=0.063
c53 24 VSS 0.00514955f $X=0.025 $Y=0.111
c54 22 VSS 0.00108941f $X=0.027 $Y=0.225
c55 20 VSS 0.00760555f $X=0.324 $Y=0.2025
c56 16 VSS 6.5312e-19 $X=0.341 $Y=0.2025
c57 15 VSS 0.00770771f $X=0.108 $Y=0.2025
c58 11 VSS 6.5312e-19 $X=0.125 $Y=0.2025
c59 9 VSS 4.01171e-19 $X=0.376 $Y=0.0675
c60 1 VSS 4.01171e-19 $X=0.071 $Y=0.0675
r61 66 67 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.4005 $Y2=0.036
r62 65 67 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.036 $X2=0.4005 $Y2=0.036
r63 62 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.396 $Y2=0.036
r64 62 63 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r65 58 59 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.045 $Y2=0.036
r66 56 59 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.045 $Y2=0.036
r67 56 57 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r68 53 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.036 $Y2=0.036
r69 51 52 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.207 $X2=0.405 $Y2=0.216
r70 50 51 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.154 $X2=0.405 $Y2=0.207
r71 49 50 6.17901 $w=1.8e-08 $l=9.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.063 $X2=0.405 $Y2=0.154
r72 48 52 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.216
r73 47 65 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.036
r74 47 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.063
r75 45 46 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.369
+ $Y=0.234 $X2=0.3825 $Y2=0.234
r76 44 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.369 $Y2=0.234
r77 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r78 41 42 12.2222 $w=1.8e-08 $l=1.8e-07 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.306 $Y2=0.234
r79 39 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.342 $Y2=0.234
r80 39 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.306 $Y2=0.234
r81 36 37 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.099 $Y2=0.234
r82 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r83 34 35 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.234 $X2=0.072 $Y2=0.234
r84 32 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r85 32 37 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.099 $Y2=0.234
r86 30 34 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.063 $Y2=0.234
r87 29 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r88 29 46 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.3825 $Y2=0.234
r89 27 28 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.2 $X2=0.027 $Y2=0.207
r90 25 26 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.063 $X2=0.027 $Y2=0.087
r91 24 27 6.04321 $w=1.8e-08 $l=8.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.111 $X2=0.027 $Y2=0.2
r92 24 26 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.111 $X2=0.027 $Y2=0.087
r93 22 30 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.225 $X2=0.036 $Y2=0.234
r94 22 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.207
r95 21 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.036
r96 21 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.063
r97 20 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r98 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r99 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r100 15 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r101 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r102 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r103 9 63 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r104 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.376 $Y2=0.0675
r105 4 57 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r106 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./OAI21x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI21x1_ASAP7_75t_L  VSS VDD B A1 A2 Y
* 
* Y	Y
* A2	A2
* A1	A1
* B	B
M0 noxref_6 N_B_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_A1_M1_g noxref_6 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_6 N_A2_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_6 N_A2_M3_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 VSS N_A1_M4_g noxref_6 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_6 N_B_M5_g N_Y_M5_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 N_Y_M6_d N_B_M6_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M7 N_Y_M7_d N_A1_M7_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 noxref_8 N_A2_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 noxref_9 N_A2_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 N_Y_M10_d N_A1_M10_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_Y_M11_d N_B_M11_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "OAI21x1_ASAP7_75t_L.pex.sp.OAI21X1_ASAP7_75T_L.pxi"
* BEGIN of "./OAI21x1_ASAP7_75t_L.pex.sp.OAI21X1_ASAP7_75T_L.pxi"
* File: OAI21x1_ASAP7_75t_L.pex.sp.OAI21X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:52:33 2017
* 
x_PM_OAI21X1_ASAP7_75T_L%B N_B_M0_g N_B_c_3_p N_B_M6_g N_B_M5_g N_B_c_6_p
+ N_B_M11_g B N_B_c_21_p N_B_c_7_p N_B_c_36_p N_B_c_31_p N_B_c_22_p N_B_c_2_p
+ N_B_c_10_p N_B_c_18_p N_B_c_17_p N_B_c_11_p N_B_c_5_p N_B_c_26_p N_B_c_27_p
+ N_B_c_13_p N_B_c_28_p N_B_c_20_p VSS PM_OAI21X1_ASAP7_75T_L%B
x_PM_OAI21X1_ASAP7_75T_L%A1 N_A1_M1_g N_A1_c_41_n N_A1_M7_g N_A1_M4_g
+ N_A1_c_44_n N_A1_M10_g A1 N_A1_c_47_n N_A1_c_74_p N_A1_c_72_p N_A1_c_48_n
+ N_A1_c_49_n N_A1_c_61_p N_A1_c_57_p N_A1_c_50_n N_A1_c_64_p N_A1_c_69_p VSS
+ PM_OAI21X1_ASAP7_75T_L%A1
x_PM_OAI21X1_ASAP7_75T_L%A2 N_A2_M2_g N_A2_M8_g N_A2_M3_g N_A2_c_88_n N_A2_M9_g
+ A2 VSS PM_OAI21X1_ASAP7_75T_L%A2
x_PM_OAI21X1_ASAP7_75T_L%Y N_Y_M0_s N_Y_M5_s N_Y_M7_d N_Y_M6_d N_Y_c_102_n
+ N_Y_M11_d N_Y_M10_d N_Y_c_113_n Y N_Y_c_104_n N_Y_c_105_n N_Y_c_114_n
+ N_Y_c_107_n N_Y_c_109_n N_Y_c_117_n N_Y_c_122_n N_Y_c_110_n N_Y_c_111_n
+ N_Y_c_125_n VSS PM_OAI21X1_ASAP7_75T_L%Y
cc_1 N_B_M0_g N_A1_M1_g 0.00354623f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_B_c_2_p N_A1_M1_g 2.52885e-19 $X=0.163 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_3 N_B_c_3_p N_A1_c_41_n 9.56181e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_B_M5_g N_A1_M4_g 0.00354623f $X=0.351 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_5 N_B_c_5_p N_A1_M4_g 3.05028e-19 $X=0.306 $Y=0.072 $X2=0.297 $Y2=0.0675
cc_6 N_B_c_6_p N_A1_c_44_n 9.56181e-19 $X=0.351 $Y=0.135 $X2=0.297 $Y2=0.135
cc_7 N_B_c_7_p A1 0.00195534f $X=0.081 $Y=0.11725 $X2=0.1345 $Y2=0.1355
cc_8 N_B_c_2_p A1 0.00373908f $X=0.163 $Y=0.072 $X2=0.1345 $Y2=0.1355
cc_9 B N_A1_c_47_n 0.00195534f $X=0.0835 $Y=0.1355 $X2=0.135 $Y2=0.18
cc_10 N_B_c_10_p N_A1_c_48_n 2.44969e-19 $X=0.19 $Y=0.072 $X2=0.163 $Y2=0.198
cc_11 N_B_c_11_p N_A1_c_49_n 2.44969e-19 $X=0.288 $Y=0.072 $X2=0.19 $Y2=0.198
cc_12 N_B_c_5_p N_A1_c_50_n 8.29113e-19 $X=0.306 $Y=0.072 $X2=0.297 $Y2=0.136
cc_13 N_B_c_13_p N_A1_c_50_n 0.00147448f $X=0.351 $Y=0.136 $X2=0.297 $Y2=0.136
cc_14 N_B_M0_g N_A2_M2_g 2.63406e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_15 N_B_c_10_p N_A2_M2_g 2.19803e-19 $X=0.19 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_16 N_B_M5_g N_A2_M3_g 2.63406e-19 $X=0.351 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_17 N_B_c_17_p N_A2_M3_g 3.48794e-19 $X=0.256 $Y=0.072 $X2=0.297 $Y2=0.0675
cc_18 N_B_c_18_p A2 0.00368224f $X=0.227 $Y=0.072 $X2=0.135 $Y2=0.189
cc_19 N_B_c_17_p A2 9.10799e-19 $X=0.256 $Y=0.072 $X2=0.135 $Y2=0.189
cc_20 N_B_c_20_p A2 2.41734e-19 $X=0.351 $Y=0.119 $X2=0.135 $Y2=0.189
cc_21 VSS N_B_c_21_p 5.94525e-19 $X=0.081 $Y=0.099 $X2=0.135 $Y2=0.189
cc_22 VSS N_B_c_22_p 0.0016619f $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.189
cc_23 VSS N_B_c_18_p 0.00191933f $X=0.227 $Y=0.072 $X2=0.135 $Y2=0.136
cc_24 VSS N_B_c_17_p 4.19603e-19 $X=0.256 $Y=0.072 $X2=0.135 $Y2=0.136
cc_25 VSS N_B_c_22_p 0.0195441f $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.18
cc_26 VSS N_B_c_26_p 0.00164678f $X=0.333 $Y=0.072 $X2=0.288 $Y2=0.198
cc_27 VSS N_B_c_27_p 2.08682e-19 $X=0.3375 $Y=0.072 $X2=0.288 $Y2=0.198
cc_28 VSS N_B_c_28_p 6.39016e-19 $X=0.351 $Y=0.099 $X2=0.288 $Y2=0.198
cc_29 B N_Y_c_102_n 0.00114532f $X=0.0835 $Y=0.1355 $X2=0.297 $Y2=0.2025
cc_30 N_B_c_7_p Y 0.00260242f $X=0.081 $Y=0.11725 $X2=0.135 $Y2=0.18
cc_31 N_B_c_31_p N_Y_c_104_n 0.00260242f $X=0.09 $Y=0.072 $X2=0.144 $Y2=0.198
cc_32 N_B_M0_g N_Y_c_105_n 2.56935e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_33 B N_Y_c_105_n 0.00123678f $X=0.0835 $Y=0.1355 $X2=0 $Y2=0
cc_34 N_B_M5_g N_Y_c_107_n 3.7308e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_B_c_13_p N_Y_c_107_n 4.52873e-19 $X=0.351 $Y=0.136 $X2=0 $Y2=0
cc_36 N_B_c_36_p N_Y_c_109_n 0.003707f $X=0.342 $Y=0.072 $X2=0 $Y2=0
cc_37 N_B_c_31_p N_Y_c_110_n 0.00135988f $X=0.09 $Y=0.072 $X2=0 $Y2=0
cc_38 N_B_c_36_p N_Y_c_111_n 0.00135988f $X=0.342 $Y=0.072 $X2=0 $Y2=0
cc_39 N_A1_M1_g N_A2_M2_g 0.0031831f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_40 N_A1_M4_g N_A2_M2_g 2.34385e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_41 N_A1_c_49_n N_A2_M2_g 2.19803e-19 $X=0.19 $Y=0.198 $X2=0.081 $Y2=0.0675
cc_42 N_A1_M1_g N_A2_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_43 N_A1_M4_g N_A2_M3_g 0.0031831f $X=0.297 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_44 N_A1_c_57_p N_A2_M3_g 3.45411e-19 $X=0.256 $Y=0.198 $X2=0.351 $Y2=0.0675
cc_45 N_A1_c_41_n N_A2_c_88_n 0.0010272f $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.135
cc_46 N_A1_c_44_n N_A2_c_88_n 0.00123834f $X=0.297 $Y=0.135 $X2=0.351 $Y2=0.135
cc_47 A1 A2 0.00322057f $X=0.1345 $Y=0.1355 $X2=0.081 $Y2=0.1355
cc_48 N_A1_c_61_p A2 0.00368242f $X=0.227 $Y=0.198 $X2=0.081 $Y2=0.1355
cc_49 N_A1_c_57_p A2 9.58063e-19 $X=0.256 $Y=0.198 $X2=0.081 $Y2=0.1355
cc_50 N_A1_c_50_n A2 0.00105444f $X=0.297 $Y=0.136 $X2=0.081 $Y2=0.1355
cc_51 N_A1_c_64_p A2 7.41132e-19 $X=0.297 $Y=0.154 $X2=0.081 $Y2=0.1355
cc_52 VSS A1 2.75878e-19 $X=0.1345 $Y=0.1355 $X2=0.081 $Y2=0.1355
cc_53 VSS N_A1_M1_g 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_54 VSS N_A1_M4_g 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_55 A1 N_Y_c_102_n 0.00162296f $X=0.1345 $Y=0.1355 $X2=0.351 $Y2=0.2025
cc_56 N_A1_c_69_p N_Y_c_113_n 0.00180096f $X=0.297 $Y=0.171 $X2=0.081 $Y2=0.099
cc_57 N_A1_M1_g N_Y_c_114_n 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0.351 $Y2=0.119
cc_58 N_A1_M4_g N_Y_c_114_n 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0.351 $Y2=0.119
cc_59 N_A1_c_72_p N_Y_c_114_n 0.016421f $X=0.144 $Y=0.198 $X2=0.351 $Y2=0.119
cc_60 N_A1_c_69_p N_Y_c_117_n 4.95573e-19 $X=0.297 $Y=0.171 $X2=0 $Y2=0
cc_61 VSS N_A1_c_74_p 2.44151e-19 $X=0.288 $Y=0.198 $X2=0.081 $Y2=0.0675
cc_62 VSS N_A2_c_88_n 3.51308e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_63 VSS N_A2_c_88_n 7.78051e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.136
cc_64 VSS A2 0.00161796f $X=0.2085 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_65 VSS N_A2_M2_g 2.64781e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_66 VSS N_A2_M3_g 2.64781e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_67 N_A2_M2_g N_Y_c_114_n 2.64781e-19 $X=0.189 $Y=0.0675 $X2=0.351 $Y2=0.119
cc_68 N_A2_M3_g N_Y_c_114_n 2.60867e-19 $X=0.243 $Y=0.0675 $X2=0.351 $Y2=0.119
cc_69 VSS N_Y_c_102_n 0.00122706f $X=0.108 $Y=0.036 $X2=0.351 $Y2=0.2025
cc_70 VSS N_Y_c_113_n 0.00122706f $X=0.324 $Y=0.036 $X2=0.081 $Y2=0.099
cc_71 VSS N_Y_c_122_n 6.57673e-19 $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_72 VSS N_Y_c_110_n 0.00379431f $X=0.108 $Y=0.036 $X2=0 $Y2=0
cc_73 VSS N_Y_c_111_n 0.00363401f $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_74 VSS N_Y_c_125_n 6.57673e-19 $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_75 VSS N_Y_c_114_n 2.33741e-19 $X=0.306 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_76 VSS N_Y_c_114_n 2.33741e-19 $X=0.306 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./OAI21x1_ASAP7_75t_L.pex.sp.OAI21X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI21xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:52:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI21xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI21xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI21xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:52:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI21XP33_ASAP7_75T_L%A1 2 5 7 12 16 VSS
c15 16 VSS 0.00911953f $X=0.064 $Y=0.136
c16 12 VSS 0.00588112f $X=0.065 $Y=0.115
c17 5 VSS 0.00502111f $X=0.081 $Y=0.135
c18 2 VSS 0.06629f $X=0.081 $Y=0.054
r19 16 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.136 $X2=0.064
+ $Y2=0.136
r20 12 16 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.115 $X2=0.064 $Y2=0.136
r21 5 17 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r22 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r23 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI21XP33_ASAP7_75T_L%A2 2 5 7 10 13 VSS
c12 13 VSS 8.0378e-19 $X=0.135 $Y=0.135
c13 10 VSS 4.06577e-19 $X=0.134 $Y=0.121
c14 5 VSS 0.00126471f $X=0.135 $Y=0.135
c15 2 VSS 0.0616076f $X=0.135 $Y=0.054
r16 10 13 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.121 $X2=0.135 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r18 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r19 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI21XP33_ASAP7_75T_L%B 2 5 7 10 VSS
c9 10 VSS 4.01588e-19 $X=0.193 $Y=0.115
c10 5 VSS 0.00170582f $X=0.189 $Y=0.135
c11 2 VSS 0.064013f $X=0.189 $Y=0.054
r12 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI21XP33_ASAP7_75T_L%Y 1 2 5 6 7 10 16 17 19 21 27 28 32 34 36 VSS
c20 36 VSS 0.00171123f $X=0.243 $Y=0.203
c21 34 VSS 6.47494e-19 $X=0.243 $Y=0.1205
c22 33 VSS 0.00129279f $X=0.243 $Y=0.106
c23 32 VSS 0.00229863f $X=0.241 $Y=0.135
c24 30 VSS 0.0011491f $X=0.243 $Y=0.225
c25 28 VSS 0.00146362f $X=0.198 $Y=0.234
c26 27 VSS 0.00370118f $X=0.18 $Y=0.234
c27 22 VSS 0.00921815f $X=0.234 $Y=0.234
c28 21 VSS 5.31938e-19 $X=0.198 $Y=0.072
c29 20 VSS 2.03419e-19 $X=0.18 $Y=0.072
c30 19 VSS 3.19168e-19 $X=0.176 $Y=0.072
c31 18 VSS 1.23838e-19 $X=0.148 $Y=0.072
c32 17 VSS 8.46035e-21 $X=0.144 $Y=0.072
c33 16 VSS 7.23848e-19 $X=0.126 $Y=0.072
c34 11 VSS 0.00714041f $X=0.234 $Y=0.072
c35 10 VSS 0.005984f $X=0.162 $Y=0.216
c36 6 VSS 5.65078e-19 $X=0.179 $Y=0.216
c37 5 VSS 0.00220525f $X=0.108 $Y=0.054
c38 1 VSS 5.98214e-19 $X=0.125 $Y=0.054
r39 35 36 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.171 $X2=0.243 $Y2=0.203
r40 33 34 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.106 $X2=0.243 $Y2=0.1205
r41 32 35 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.171
r42 32 34 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.1205
r43 30 36 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.203
r44 29 33 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.106
r45 27 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r46 24 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r47 22 30 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r48 22 28 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.198 $Y2=0.234
r49 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.072 $X2=0.198 $Y2=0.072
r50 19 20 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.072 $X2=0.18 $Y2=0.072
r51 18 19 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.072 $X2=0.176 $Y2=0.072
r52 17 18 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.148 $Y2=0.072
r53 16 17 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.144 $Y2=0.072
r54 13 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.126 $Y2=0.072
r55 11 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.072 $X2=0.243 $Y2=0.081
r56 11 21 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.198 $Y2=0.072
r57 10 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r58 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.162 $Y2=0.216
r59 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.216 $X2=0.162 $Y2=0.216
r60 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072 $X2=0.108
+ $Y2=0.072
r61 2 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.054 $X2=0.108 $Y2=0.054
r62 1 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.054 $X2=0.108 $Y2=0.054
.ends


* END of "./OAI21xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI21xp33_ASAP7_75t_L  VSS VDD A1 A2 B Y
* 
* Y	Y
* B	B
* A2	A2
* A1	A1
M0 N_Y_M0_d N_A1_M0_g noxref_6 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 noxref_6 N_A2_M1_g N_Y_M1_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 VSS N_B_M2_g noxref_6 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 noxref_8 N_A1_M3_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M4 N_Y_M4_d N_A2_M4_g noxref_8 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M5 VDD N_B_M5_g N_Y_M5_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.189
*
* 
* .include "OAI21xp33_ASAP7_75t_L.pex.sp.OAI21XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI21xp33_ASAP7_75t_L.pex.sp.OAI21XP33_ASAP7_75T_L.pxi"
* File: OAI21xp33_ASAP7_75t_L.pex.sp.OAI21XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:52:56 2017
* 
x_PM_OAI21XP33_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M3_g A1 N_A1_c_15_p VSS
+ PM_OAI21XP33_ASAP7_75T_L%A1
x_PM_OAI21XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_17_n N_A2_M4_g A2 N_A2_c_19_n VSS
+ PM_OAI21XP33_ASAP7_75T_L%A2
x_PM_OAI21XP33_ASAP7_75T_L%B N_B_M2_g N_B_c_30_n N_B_M5_g B VSS
+ PM_OAI21XP33_ASAP7_75T_L%B
x_PM_OAI21XP33_ASAP7_75T_L%Y N_Y_M1_s N_Y_M0_d N_Y_c_37_n N_Y_M5_s N_Y_M4_d
+ N_Y_c_38_n N_Y_c_39_n N_Y_c_42_n N_Y_c_56_n N_Y_c_45_n N_Y_c_40_n N_Y_c_47_n Y
+ N_Y_c_49_n N_Y_c_44_n VSS PM_OAI21XP33_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00361888f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A1_c_2_p N_A2_c_17_n 0.00106637f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A1 A2 0.00161558f $X=0.065 $Y=0.115 $X2=0.134 $Y2=0.121
cc_4 A1 N_A2_c_19_n 0.00161558f $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.135
cc_5 N_A1_M0_g N_B_M2_g 2.98169e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_6 VSS A1 2.8176e-19 $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.054
cc_7 VSS N_A1_c_2_p 2.13815e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_8 VSS A1 0.00297211f $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.135
cc_9 VSS A1 0.003244f $X=0.065 $Y=0.115 $X2=0 $Y2=0
cc_10 VSS N_A1_M0_g 2.39633e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_11 VSS N_A1_c_2_p 3.09341e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_12 A1 N_Y_c_37_n 2.60799e-19 $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.135
cc_13 A1 N_Y_c_38_n 3.19189e-19 $X=0.065 $Y=0.115 $X2=0.134 $Y2=0.121
cc_14 A1 N_Y_c_39_n 0.00129324f $X=0.065 $Y=0.115 $X2=0 $Y2=0
cc_15 N_A1_c_15_p N_Y_c_40_n 5.36322e-19 $X=0.064 $Y=0.136 $X2=0 $Y2=0
cc_16 N_A2_M1_g N_B_M2_g 0.00354623f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_17 N_A2_c_17_n N_B_c_30_n 9.33263e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_18 A2 B 0.00334765f $X=0.134 $Y=0.121 $X2=0 $Y2=0
cc_19 VSS N_A2_M1_g 2.38303e-19 $X=0.135 $Y=0.054 $X2=0.064 $Y2=0.136
cc_20 N_A2_c_19_n N_Y_c_38_n 5.59664e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_21 N_A2_M1_g N_Y_c_42_n 2.76185e-19 $X=0.135 $Y=0.054 $X2=0.064 $Y2=0.136
cc_22 A2 N_Y_c_42_n 0.00123279f $X=0.134 $Y=0.121 $X2=0.064 $Y2=0.136
cc_23 N_A2_c_19_n N_Y_c_44_n 5.00837e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_24 N_B_M2_g N_Y_c_45_n 3.62029e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_25 B N_Y_c_45_n 0.00122403f $X=0.193 $Y=0.115 $X2=0 $Y2=0
cc_26 N_B_M2_g N_Y_c_47_n 3.43731e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_27 B N_Y_c_47_n 6.07428e-19 $X=0.193 $Y=0.115 $X2=0 $Y2=0
cc_28 B N_Y_c_49_n 0.00329908f $X=0.193 $Y=0.115 $X2=0 $Y2=0
cc_29 VSS N_Y_c_37_n 0.00297277f $X=0.056 $Y=0.054 $X2=0.081 $Y2=0.135
cc_30 VSS N_Y_c_37_n 0.00299929f $X=0.162 $Y=0.054 $X2=0.081 $Y2=0.135
cc_31 VSS N_Y_c_37_n 0.00189275f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_32 VSS N_Y_c_37_n 6.2062e-19 $X=0.099 $Y=0.036 $X2=0.081 $Y2=0.135
cc_33 VSS N_Y_c_38_n 4.54531e-19 $X=0.162 $Y=0.054 $X2=0 $Y2=0
cc_34 VSS N_Y_c_39_n 0.00666759f $X=0.162 $Y=0.036 $X2=0.064 $Y2=0.136
cc_35 VSS N_Y_c_56_n 0.00343253f $X=0.162 $Y=0.054 $X2=0 $Y2=0

* END of "./OAI21xp33_ASAP7_75t_L.pex.sp.OAI21XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI21xp5_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:53:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI21xp5_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI21xp5_ASAP7_75t_L.pex.sp.pex"
* File: OAI21xp5_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:53:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI21XP5_ASAP7_75T_L%A1 2 5 7 12 16 VSS
c15 16 VSS 0.00902761f $X=0.064 $Y=0.136
c16 12 VSS 0.00597343f $X=0.065 $Y=0.115
c17 5 VSS 0.00611347f $X=0.081 $Y=0.135
c18 2 VSS 0.06629f $X=0.081 $Y=0.0675
r19 16 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.136 $X2=0.064
+ $Y2=0.136
r20 12 16 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.115 $X2=0.064 $Y2=0.136
r21 5 17 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI21XP5_ASAP7_75T_L%A2 2 5 7 10 13 VSS
c12 13 VSS 6.15402e-19 $X=0.135 $Y=0.135
c13 10 VSS 4.45038e-19 $X=0.134 $Y=0.121
c14 5 VSS 0.00126471f $X=0.135 $Y=0.135
c15 2 VSS 0.0616076f $X=0.135 $Y=0.0675
r16 10 13 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.121 $X2=0.135 $Y2=0.135
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI21XP5_ASAP7_75T_L%B 2 5 7 10 VSS
c10 10 VSS 7.15852e-19 $X=0.193 $Y=0.115
c11 5 VSS 0.00170582f $X=0.189 $Y=0.135
c12 2 VSS 0.064013f $X=0.189 $Y=0.0675
r13 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.115 $X2=0.189 $Y2=0.135
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI21XP5_ASAP7_75T_L%Y 1 2 5 6 7 10 16 17 19 21 27 28 32 34 36 VSS
c22 36 VSS 0.00176181f $X=0.243 $Y=0.203
c23 34 VSS 6.503e-19 $X=0.243 $Y=0.1205
c24 33 VSS 0.0012886f $X=0.243 $Y=0.106
c25 32 VSS 0.00231091f $X=0.241 $Y=0.135
c26 30 VSS 0.00112227f $X=0.243 $Y=0.225
c27 28 VSS 0.00146362f $X=0.198 $Y=0.234
c28 27 VSS 0.00371408f $X=0.18 $Y=0.234
c29 22 VSS 0.00920004f $X=0.234 $Y=0.234
c30 21 VSS 5.31938e-19 $X=0.198 $Y=0.072
c31 20 VSS 2.03419e-19 $X=0.18 $Y=0.072
c32 19 VSS 2.44387e-19 $X=0.176 $Y=0.072
c33 18 VSS 1.23838e-19 $X=0.148 $Y=0.072
c34 17 VSS 8.46035e-21 $X=0.144 $Y=0.072
c35 16 VSS 7.46535e-19 $X=0.126 $Y=0.072
c36 11 VSS 0.0060196f $X=0.234 $Y=0.072
c37 10 VSS 0.00754825f $X=0.162 $Y=0.2025
c38 6 VSS 5.72268e-19 $X=0.179 $Y=0.2025
c39 5 VSS 0.00241636f $X=0.108 $Y=0.0675
c40 1 VSS 6.411e-19 $X=0.125 $Y=0.0675
r41 35 36 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.171 $X2=0.243 $Y2=0.203
r42 33 34 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.106 $X2=0.243 $Y2=0.1205
r43 32 35 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.171
r44 32 34 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.1205
r45 30 36 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.203
r46 29 33 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.106
r47 27 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r48 24 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r49 22 30 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r50 22 28 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.198 $Y2=0.234
r51 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.072 $X2=0.198 $Y2=0.072
r52 19 20 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.072 $X2=0.18 $Y2=0.072
r53 18 19 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.072 $X2=0.176 $Y2=0.072
r54 17 18 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.148 $Y2=0.072
r55 16 17 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.144 $Y2=0.072
r56 13 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.126 $Y2=0.072
r57 11 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.072 $X2=0.243 $Y2=0.081
r58 11 21 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.198 $Y2=0.072
r59 10 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r60 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r61 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r62 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072 $X2=0.108
+ $Y2=0.072
r63 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r64 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OAI21xp5_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI21xp5_ASAP7_75t_L  VSS VDD A1 A2 B Y
* 
* Y	Y
* B	B
* A2	A2
* A1	A1
M0 N_Y_M0_d N_A1_M0_g noxref_6 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_6 N_A2_M1_g N_Y_M1_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_B_M2_g noxref_6 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 noxref_8 N_A1_M3_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M4 N_Y_M4_d N_A2_M4_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M5 VDD N_B_M5_g N_Y_M5_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
*
* 
* .include "OAI21xp5_ASAP7_75t_L.pex.sp.OAI21XP5_ASAP7_75T_L.pxi"
* BEGIN of "./OAI21xp5_ASAP7_75t_L.pex.sp.OAI21XP5_ASAP7_75T_L.pxi"
* File: OAI21xp5_ASAP7_75t_L.pex.sp.OAI21XP5_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:53:18 2017
* 
x_PM_OAI21XP5_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M3_g A1 N_A1_c_15_p VSS
+ PM_OAI21XP5_ASAP7_75T_L%A1
x_PM_OAI21XP5_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_17_n N_A2_M4_g A2 N_A2_c_19_n VSS
+ PM_OAI21XP5_ASAP7_75T_L%A2
x_PM_OAI21XP5_ASAP7_75T_L%B N_B_M2_g N_B_c_30_n N_B_M5_g B VSS
+ PM_OAI21XP5_ASAP7_75T_L%B
x_PM_OAI21XP5_ASAP7_75T_L%Y N_Y_M1_s N_Y_M0_d N_Y_c_38_n N_Y_M5_s N_Y_M4_d
+ N_Y_c_39_n N_Y_c_40_n N_Y_c_43_n N_Y_c_59_n N_Y_c_47_n N_Y_c_41_n N_Y_c_49_n Y
+ N_Y_c_51_n N_Y_c_45_n VSS PM_OAI21XP5_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00361888f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_17_n 0.00106637f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A1 A2 0.00154447f $X=0.065 $Y=0.115 $X2=0.134 $Y2=0.121
cc_4 A1 N_A2_c_19_n 0.00154447f $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.135
cc_5 N_A1_M0_g N_B_M2_g 2.98169e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 VSS A1 2.11432e-19 $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.0675
cc_7 VSS N_A1_c_2_p 4.0003e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_8 VSS A1 0.00353122f $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.135
cc_9 VSS A1 0.00324399f $X=0.065 $Y=0.115 $X2=0 $Y2=0
cc_10 VSS N_A1_M0_g 2.39633e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_11 VSS N_A1_c_2_p 3.09341e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_12 A1 N_Y_c_38_n 7.8712e-19 $X=0.065 $Y=0.115 $X2=0.135 $Y2=0.135
cc_13 A1 N_Y_c_39_n 3.61515e-19 $X=0.065 $Y=0.115 $X2=0.134 $Y2=0.121
cc_14 A1 N_Y_c_40_n 0.00129324f $X=0.065 $Y=0.115 $X2=0 $Y2=0
cc_15 N_A1_c_15_p N_Y_c_41_n 5.36322e-19 $X=0.064 $Y=0.136 $X2=0 $Y2=0
cc_16 N_A2_M1_g N_B_M2_g 0.00354623f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 N_A2_c_17_n N_B_c_30_n 9.33263e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_18 A2 B 0.00307202f $X=0.134 $Y=0.121 $X2=0 $Y2=0
cc_19 VSS N_A2_M1_g 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0.064 $Y2=0.136
cc_20 A2 N_Y_c_39_n 0.00158986f $X=0.134 $Y=0.121 $X2=0 $Y2=0
cc_21 N_A2_M1_g N_Y_c_43_n 2.76185e-19 $X=0.135 $Y=0.0675 $X2=0.064 $Y2=0.136
cc_22 A2 N_Y_c_43_n 0.00123279f $X=0.134 $Y=0.121 $X2=0.064 $Y2=0.136
cc_23 N_A2_c_19_n N_Y_c_45_n 2.44454e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_24 B N_Y_c_39_n 2.71261e-19 $X=0.193 $Y=0.115 $X2=0 $Y2=0
cc_25 N_B_M2_g N_Y_c_47_n 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 B N_Y_c_47_n 0.00122403f $X=0.193 $Y=0.115 $X2=0 $Y2=0
cc_27 N_B_M2_g N_Y_c_49_n 3.43731e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_28 B N_Y_c_49_n 6.07428e-19 $X=0.193 $Y=0.115 $X2=0 $Y2=0
cc_29 B N_Y_c_51_n 0.00303518f $X=0.193 $Y=0.115 $X2=0 $Y2=0
cc_30 VSS N_Y_M1_s 2.09551e-19 $X=0.099 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_31 VSS N_Y_c_38_n 0.00391978f $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.135
cc_32 VSS N_Y_c_38_n 0.00189275f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_33 VSS N_Y_c_38_n 0.0035205f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_34 VSS N_Y_c_38_n 6.2062e-19 $X=0.099 $Y=0.036 $X2=0.081 $Y2=0.135
cc_35 VSS N_Y_c_39_n 0.00138157f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_36 VSS N_Y_c_40_n 0.00666757f $X=0.162 $Y=0.036 $X2=0.064 $Y2=0.136
cc_37 VSS N_Y_c_59_n 0.00233206f $X=0.162 $Y=0.036 $X2=0 $Y2=0

* END of "./OAI21xp5_ASAP7_75t_L.pex.sp.OAI21XP5_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI221xp5_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:53:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI221xp5_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI221xp5_ASAP7_75t_L.pex.sp.pex"
* File: OAI221xp5_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:53:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI221XP5_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c11 10 VSS 6.95749e-19 $X=0.081 $Y=0.135
c12 5 VSS 0.00172166f $X=0.081 $Y=0.135
c13 2 VSS 0.0655264f $X=0.081 $Y=0.0675
r14 10 14 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.148
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI221XP5_ASAP7_75T_L%B2 2 5 7 10 VSS
c11 10 VSS 0.00105185f $X=0.134 $Y=0.109
c12 5 VSS 0.00113686f $X=0.135 $Y=0.135
c13 2 VSS 0.0607967f $X=0.135 $Y=0.0675
r14 10 13 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.109 $X2=0.135 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI221XP5_ASAP7_75T_L%C 2 5 7 10 VSS
c11 10 VSS 0.00138457f $X=0.188 $Y=0.123
c12 5 VSS 0.00120113f $X=0.189 $Y=0.135
c13 2 VSS 0.0599921f $X=0.189 $Y=0.0675
r14 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.123 $X2=0.189 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI221XP5_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c10 10 VSS 0.00122183f $X=0.243 $Y=0.135
c11 5 VSS 0.00124202f $X=0.243 $Y=0.135
c12 2 VSS 0.05968f $X=0.243 $Y=0.0675
r13 10 14 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.169
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI221XP5_ASAP7_75T_L%A2 2 5 7 10 13 VSS
c8 13 VSS 0.00301998f $X=0.297 $Y=0.135
c9 10 VSS 0.00214663f $X=0.295 $Y=0.123
c10 5 VSS 0.00230503f $X=0.297 $Y=0.135
c11 2 VSS 0.0631596f $X=0.297 $Y=0.0675
r12 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.123 $X2=0.297 $Y2=0.135
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OAI221XP5_ASAP7_75T_L%Y 1 2 5 6 9 11 12 15 19 20 21 26 29 30 38 41 44
+ 47 VSS
c25 49 VSS 9.42062e-19 $X=0.2085 $Y=0.234
c26 48 VSS 2.39163e-19 $X=0.201 $Y=0.234
c27 47 VSS 0.00146362f $X=0.198 $Y=0.234
c28 46 VSS 3.78291e-19 $X=0.18 $Y=0.234
c29 45 VSS 0.00558992f $X=0.176 $Y=0.234
c30 44 VSS 0.00142296f $X=0.144 $Y=0.234
c31 43 VSS 3.47945e-19 $X=0.126 $Y=0.234
c32 42 VSS 0.00315399f $X=0.123 $Y=0.234
c33 41 VSS 0.00146362f $X=0.09 $Y=0.234
c34 40 VSS 0.00368249f $X=0.072 $Y=0.234
c35 38 VSS 0.00283822f $X=0.216 $Y=0.234
c36 33 VSS 0.00336615f $X=0.036 $Y=0.234
c37 31 VSS 1.45514e-19 $X=0.099 $Y=0.072
c38 30 VSS 8.46035e-21 $X=0.09 $Y=0.072
c39 29 VSS 3.46932e-19 $X=0.072 $Y=0.072
c40 28 VSS 2.30435e-19 $X=0.04 $Y=0.072
c41 26 VSS 3.3737e-19 $X=0.108 $Y=0.072
c42 24 VSS 0.0019286f $X=0.036 $Y=0.072
c43 23 VSS 5.10117e-19 $X=0.027 $Y=0.2125
c44 21 VSS 0.00149783f $X=0.027 $Y=0.139
c45 20 VSS 0.00112176f $X=0.027 $Y=0.106
c46 19 VSS 0.00273404f $X=0.025 $Y=0.172
c47 17 VSS 6.07272e-19 $X=0.027 $Y=0.225
c48 15 VSS 0.00606778f $X=0.216 $Y=0.216
c49 11 VSS 5.5175e-19 $X=0.233 $Y=0.216
c50 9 VSS 0.00319205f $X=0.056 $Y=0.216
c51 6 VSS 2.6657e-19 $X=0.071 $Y=0.216
c52 5 VSS 0.00233317f $X=0.108 $Y=0.0675
c53 1 VSS 5.68239e-19 $X=0.125 $Y=0.0675
r54 48 49 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.201
+ $Y=0.234 $X2=0.2085 $Y2=0.234
r55 47 48 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.201 $Y2=0.234
r56 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r57 45 46 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.234 $X2=0.18 $Y2=0.234
r58 44 45 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.176 $Y2=0.234
r59 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r60 42 43 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.123
+ $Y=0.234 $X2=0.126 $Y2=0.234
r61 41 42 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.123 $Y2=0.234
r62 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r63 38 49 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.2085 $Y2=0.234
r64 35 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.072 $Y2=0.234
r65 33 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.054 $Y2=0.234
r66 30 31 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.099 $Y2=0.072
r67 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.072 $X2=0.09 $Y2=0.072
r68 28 29 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.072 $X2=0.072 $Y2=0.072
r69 26 31 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.099 $Y2=0.072
r70 24 28 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.072 $X2=0.04 $Y2=0.072
r71 22 23 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.2 $X2=0.027 $Y2=0.2125
r72 20 21 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.106 $X2=0.027 $Y2=0.139
r73 19 22 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.172 $X2=0.027 $Y2=0.2
r74 19 21 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.172 $X2=0.027 $Y2=0.139
r75 17 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.225 $X2=0.036 $Y2=0.234
r76 17 23 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.2125
r77 16 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.081 $X2=0.036 $Y2=0.072
r78 16 20 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.081 $X2=0.027 $Y2=0.106
r79 15 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r80 12 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.216 $X2=0.216 $Y2=0.216
r81 11 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.216 $X2=0.216 $Y2=0.216
r82 9 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r83 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.216 $X2=0.056 $Y2=0.216
r84 5 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072 $X2=0.108
+ $Y2=0.072
r85 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r86 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OAI221xp5_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI221xp5_ASAP7_75t_L  VSS VDD B1 B2 C A1 A2 Y
* 
* Y	Y
* A2	A2
* A1	A1
* C	C
* B2	B2
* B1	B1
M0 N_Y_M0_d N_B1_M0_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_9 N_B2_M1_g N_Y_M1_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_10 N_C_M2_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_A1_M3_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_10 N_A2_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_11 N_B1_M5_g N_Y_M5_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M6 VDD N_B2_M6_g noxref_11 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M7 N_Y_M7_d N_C_M7_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.189
M8 noxref_12 N_A1_M8_g N_Y_M8_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M9 VDD N_A2_M9_g noxref_12 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.189
*
* 
* .include "OAI221xp5_ASAP7_75t_L.pex.sp.OAI221XP5_ASAP7_75T_L.pxi"
* BEGIN of "./OAI221xp5_ASAP7_75t_L.pex.sp.OAI221XP5_ASAP7_75T_L.pxi"
* File: OAI221xp5_ASAP7_75t_L.pex.sp.OAI221XP5_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:53:41 2017
* 
x_PM_OAI221XP5_ASAP7_75T_L%B1 N_B1_M0_g N_B1_c_2_p N_B1_M5_g N_B1_c_3_p B1 VSS
+ PM_OAI221XP5_ASAP7_75T_L%B1
x_PM_OAI221XP5_ASAP7_75T_L%B2 N_B2_M1_g N_B2_c_13_n N_B2_M6_g B2 VSS
+ PM_OAI221XP5_ASAP7_75T_L%B2
x_PM_OAI221XP5_ASAP7_75T_L%C N_C_M2_g N_C_c_25_n N_C_M7_g C VSS
+ PM_OAI221XP5_ASAP7_75T_L%C
x_PM_OAI221XP5_ASAP7_75T_L%A1 N_A1_M3_g N_A1_c_36_n N_A1_M8_g N_A1_c_37_n A1 VSS
+ PM_OAI221XP5_ASAP7_75T_L%A1
x_PM_OAI221XP5_ASAP7_75T_L%A2 N_A2_M4_g N_A2_c_46_n N_A2_M9_g A2 N_A2_c_49_p VSS
+ PM_OAI221XP5_ASAP7_75T_L%A2
x_PM_OAI221XP5_ASAP7_75T_L%Y N_Y_M1_s N_Y_M0_d N_Y_c_67_p N_Y_M5_s N_Y_c_52_n
+ N_Y_M8_s N_Y_M7_d N_Y_c_60_n Y N_Y_c_69_p N_Y_c_53_n N_Y_c_72_p N_Y_c_66_p
+ N_Y_c_54_n N_Y_c_65_n N_Y_c_56_n N_Y_c_58_n N_Y_c_61_n VSS
+ PM_OAI221XP5_ASAP7_75T_L%Y
cc_1 N_B1_M0_g N_B2_M1_g 0.00364065f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_B1_c_2_p N_B2_c_13_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_B1_c_3_p B2 0.00484691f $X=0.081 $Y=0.135 $X2=0.134 $Y2=0.109
cc_4 N_B1_M0_g N_C_M2_g 2.6588e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 N_B1_c_3_p N_Y_c_52_n 3.87865e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.109
cc_6 N_B1_c_3_p N_Y_c_53_n 0.00440946f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_7 N_B1_M0_g N_Y_c_54_n 2.68514e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_8 N_B1_c_3_p N_Y_c_54_n 0.00121543f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_B1_M0_g N_Y_c_56_n 2.64276e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_10 N_B1_c_3_p N_Y_c_56_n 0.00124805f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 VSS N_B1_M0_g 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_12 N_B2_M1_g N_C_M2_g 0.0032267f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_13 N_B2_c_13_n N_C_c_25_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 B2 C 0.00456406f $X=0.134 $Y=0.109 $X2=0.081 $Y2=0.135
cc_15 N_B2_M1_g N_A1_M3_g 2.60137e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_B2_M1_g N_Y_c_58_n 2.56935e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_17 B2 N_Y_c_58_n 0.00123064f $X=0.134 $Y=0.109 $X2=0 $Y2=0
cc_18 VSS N_B2_M1_g 3.47199e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 VSS B2 5.30079e-19 $X=0.134 $Y=0.109 $X2=0 $Y2=0
cc_20 N_C_M2_g N_A1_M3_g 0.00346636f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_21 N_C_c_25_n N_A1_c_36_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 C N_A1_c_37_n 0.00456406f $X=0.188 $Y=0.123 $X2=0.081 $Y2=0.135
cc_23 N_C_M2_g N_A2_M4_g 2.54394e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_24 C N_Y_c_60_n 3.31541e-19 $X=0.188 $Y=0.123 $X2=0 $Y2=0
cc_25 N_C_M2_g N_Y_c_61_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 C N_Y_c_61_n 0.00124805f $X=0.188 $Y=0.123 $X2=0 $Y2=0
cc_27 N_A1_M3_g N_A2_M4_g 0.00310323f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_28 N_A1_c_36_n N_A2_c_46_n 9.33263e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_29 N_A1_c_37_n A2 0.00467338f $X=0.243 $Y=0.135 $X2=0.134 $Y2=0.109
cc_30 N_A1_c_37_n N_Y_c_60_n 3.87865e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 VSS N_A1_M3_g 3.51973e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_32 VSS N_A1_c_37_n 0.00121543f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_33 A2 N_Y_c_60_n 3.94305e-19 $X=0.295 $Y=0.123 $X2=0 $Y2=0
cc_34 N_A2_c_49_p N_Y_c_65_n 4.37254e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_35 VSS N_A2_M4_g 3.51973e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_36 VSS A2 0.00122076f $X=0.295 $Y=0.123 $X2=0 $Y2=0
cc_37 VSS N_Y_c_66_p 2.47657e-19 $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_38 VSS N_Y_c_67_p 0.00371671f $X=0.108 $Y=0.0675 $X2=0.081 $Y2=0.148
cc_39 VSS N_Y_c_52_n 9.98826e-19 $X=0.056 $Y=0.216 $X2=0.081 $Y2=0.148
cc_40 VSS N_Y_c_69_p 3.97918e-19 $X=0.027 $Y=0.106 $X2=0.081 $Y2=0.148
cc_41 VSS N_Y_c_66_p 0.00260156f $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.148
cc_42 VSS N_Y_c_67_p 0.00333582f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_43 VSS N_Y_c_72_p 4.54465e-19 $X=0.108 $Y=0.072 $X2=0 $Y2=0
cc_44 VSS N_Y_c_67_p 0.00250965f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_45 VSS N_Y_c_66_p 0.00714937f $X=0.072 $Y=0.072 $X2=0 $Y2=0
cc_46 VSS N_Y_c_60_n 9.98826e-19 $X=0.216 $Y=0.216 $X2=0.081 $Y2=0.135
cc_47 VSS N_Y_c_72_p 2.95791e-19 $X=0.108 $Y=0.072 $X2=0 $Y2=0

* END of "./OAI221xp5_ASAP7_75t_L.pex.sp.OAI221XP5_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI222xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:54:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI222xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI222xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI222xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:54:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI222XP33_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c11 10 VSS 5.09652e-19 $X=0.081 $Y=0.135
c12 5 VSS 0.00171842f $X=0.081 $Y=0.135
c13 2 VSS 0.066866f $X=0.081 $Y=0.0675
r14 10 14 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.194
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI222XP33_ASAP7_75T_L%A2 2 5 7 10 VSS
c11 10 VSS 0.00167719f $X=0.135 $Y=0.119
c12 5 VSS 0.00113686f $X=0.135 $Y=0.135
c13 2 VSS 0.062389f $X=0.135 $Y=0.0675
r14 10 13 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.119 $X2=0.135 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI222XP33_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c11 10 VSS 0.00167719f $X=0.189 $Y=0.135
c12 5 VSS 0.00113407f $X=0.189 $Y=0.135
c13 2 VSS 0.062389f $X=0.189 $Y=0.0675
r14 10 14 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.172
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI222XP33_ASAP7_75T_L%B1 2 5 7 10 VSS
c11 10 VSS 7.9511e-19 $X=0.243 $Y=0.115
c12 5 VSS 0.00220625f $X=0.243 $Y=0.135
c13 2 VSS 0.0662287f $X=0.243 $Y=0.0675
r14 10 13 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.115 $X2=0.243 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI222XP33_ASAP7_75T_L%C1 2 5 7 10 15 18 VSS
c11 18 VSS 2.57027e-19 $X=0.405 $Y=0.1205
c12 15 VSS 5.34582e-19 $X=0.405 $Y=0.135
c13 10 VSS 0.00156687f $X=0.405 $Y=0.094
c14 5 VSS 0.00228295f $X=0.405 $Y=0.135
c15 2 VSS 0.0640033f $X=0.405 $Y=0.0675
r16 17 18 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.106 $X2=0.405 $Y2=0.1205
r17 15 18 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.1205
r18 10 17 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.094 $X2=0.405 $Y2=0.106
r19 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r20 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r21 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OAI222XP33_ASAP7_75T_L%C2 2 5 7 10 14 VSS
c9 10 VSS 0.00272411f $X=0.459 $Y=0.135
c10 5 VSS 0.00171373f $X=0.459 $Y=0.135
c11 2 VSS 0.0632357f $X=0.459 $Y=0.0675
r12 10 14 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.147
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OAI222XP33_ASAP7_75T_L%Y 1 2 5 6 9 11 14 16 19 23 24 27 30 31 43 44
+ 46 48 50 51 55 56 57 58 59 60 63 VSS
c37 68 VSS 7.78152e-19 $X=0.513 $Y=0.2125
c38 63 VSS 0.00816016f $X=0.516 $Y=0.147
c39 61 VSS 7.47026e-19 $X=0.513 $Y=0.225
c40 60 VSS 0.00146362f $X=0.468 $Y=0.234
c41 59 VSS 0.00346383f $X=0.45 $Y=0.234
c42 58 VSS 0.00146362f $X=0.414 $Y=0.234
c43 57 VSS 0.00271257f $X=0.396 $Y=0.234
c44 56 VSS 9.85989e-19 $X=0.369 $Y=0.234
c45 55 VSS 0.0127088f $X=0.36 $Y=0.234
c46 51 VSS 0.00146362f $X=0.252 $Y=0.234
c47 50 VSS 0.00302652f $X=0.234 $Y=0.234
c48 49 VSS 4.63288e-19 $X=0.202 $Y=0.234
c49 48 VSS 0.00142296f $X=0.198 $Y=0.234
c50 47 VSS 0.00660983f $X=0.18 $Y=0.234
c51 46 VSS 0.00142296f $X=0.144 $Y=0.234
c52 45 VSS 4.63288e-19 $X=0.126 $Y=0.234
c53 44 VSS 0.00287317f $X=0.122 $Y=0.234
c54 43 VSS 0.00146362f $X=0.09 $Y=0.234
c55 42 VSS 0.00454946f $X=0.072 $Y=0.234
c56 35 VSS 0.00327152f $X=0.027 $Y=0.234
c57 34 VSS 0.00920077f $X=0.504 $Y=0.234
c58 32 VSS 1.45514e-19 $X=0.099 $Y=0.072
c59 31 VSS 8.46035e-21 $X=0.09 $Y=0.072
c60 30 VSS 3.8564e-19 $X=0.072 $Y=0.072
c61 29 VSS 0.00112964f $X=0.04 $Y=0.072
c62 27 VSS 3.25827e-19 $X=0.108 $Y=0.072
c63 25 VSS 0.00191981f $X=0.027 $Y=0.072
c64 24 VSS 0.00432139f $X=0.018 $Y=0.2
c65 23 VSS 9.4116e-19 $X=0.018 $Y=0.106
c66 22 VSS 9.4116e-19 $X=0.018 $Y=0.225
c67 19 VSS 0.00470846f $X=0.38 $Y=0.2025
c68 16 VSS 2.69461e-19 $X=0.395 $Y=0.2025
c69 14 VSS 0.00392489f $X=0.268 $Y=0.2025
c70 9 VSS 0.00358217f $X=0.056 $Y=0.2025
c71 6 VSS 2.69461e-19 $X=0.071 $Y=0.2025
c72 5 VSS 0.0023085f $X=0.108 $Y=0.0675
c73 1 VSS 5.76042e-19 $X=0.125 $Y=0.0675
r74 67 68 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.2 $X2=0.513 $Y2=0.2125
r75 63 67 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.147 $X2=0.513 $Y2=0.2
r76 61 68 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.2125
r77 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r78 58 59 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.45 $Y2=0.234
r79 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r80 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.369 $Y2=0.234
r81 53 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r82 53 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.369 $Y2=0.234
r83 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r84 49 50 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.234 $X2=0.234 $Y2=0.234
r85 48 49 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.202 $Y2=0.234
r86 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r87 46 47 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.18 $Y2=0.234
r88 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r89 44 45 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.122
+ $Y=0.234 $X2=0.126 $Y2=0.234
r90 43 44 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.122 $Y2=0.234
r91 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r92 40 55 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.36 $Y2=0.234
r93 40 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.252 $Y2=0.234
r94 37 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.072 $Y2=0.234
r95 35 37 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.054 $Y2=0.234
r96 34 61 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.234 $X2=0.513 $Y2=0.225
r97 34 60 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.468 $Y2=0.234
r98 31 32 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.099 $Y2=0.072
r99 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.072 $X2=0.09 $Y2=0.072
r100 29 30 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.072 $X2=0.072 $Y2=0.072
r101 27 32 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.099 $Y2=0.072
r102 25 29 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.072 $X2=0.04 $Y2=0.072
r103 23 24 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.106 $X2=0.018 $Y2=0.2
r104 22 35 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r105 22 24 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2
r106 21 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.081 $X2=0.027 $Y2=0.072
r107 21 23 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.106
r108 19 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r109 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.38 $Y2=0.2025
r110 14 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r111 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.268 $Y2=0.2025
r112 9 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r113 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r114 5 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072 $X2=0.108
+ $Y2=0.072
r115 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r116 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OAI222xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI222xp33_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 C1 C2 Y
* 
* Y	Y
* C2	C2
* C1	C1
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 N_Y_M0_d N_A1_M0_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_9 N_A2_M1_g N_Y_M1_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_10 N_B2_M2_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_9 N_B1_M3_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_10 N_C1_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 VSS N_C2_M5_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 noxref_12 N_A1_M6_g N_Y_M6_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 VDD N_A2_M7_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 noxref_13 N_B2_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 N_Y_M9_d N_B1_M9_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 noxref_14 N_C1_M10_g N_Y_M10_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M11 VDD N_C2_M11_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "OAI222xp33_ASAP7_75t_L.pex.sp.OAI222XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI222xp33_ASAP7_75t_L.pex.sp.OAI222XP33_ASAP7_75T_L.pxi"
* File: OAI222xp33_ASAP7_75t_L.pex.sp.OAI222XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:54:03 2017
* 
x_PM_OAI222XP33_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M6_g N_A1_c_3_p A1 VSS
+ PM_OAI222XP33_ASAP7_75T_L%A1
x_PM_OAI222XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_13_n N_A2_M7_g A2 VSS
+ PM_OAI222XP33_ASAP7_75T_L%A2
x_PM_OAI222XP33_ASAP7_75T_L%B2 N_B2_M2_g N_B2_c_25_n N_B2_M8_g N_B2_c_26_n B2
+ VSS PM_OAI222XP33_ASAP7_75T_L%B2
x_PM_OAI222XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_36_n N_B1_M9_g B1 VSS
+ PM_OAI222XP33_ASAP7_75T_L%B1
x_PM_OAI222XP33_ASAP7_75T_L%C1 N_C1_M4_g N_C1_c_47_p N_C1_M10_g C1 N_C1_c_53_p
+ N_C1_c_45_n VSS PM_OAI222XP33_ASAP7_75T_L%C1
x_PM_OAI222XP33_ASAP7_75T_L%C2 N_C2_M5_g N_C2_c_57_n N_C2_M11_g N_C2_c_58_n C2
+ VSS PM_OAI222XP33_ASAP7_75T_L%C2
x_PM_OAI222XP33_ASAP7_75T_L%Y N_Y_M1_s N_Y_M0_d N_Y_c_84_n N_Y_M6_s N_Y_c_65_n
+ N_Y_M9_d N_Y_c_75_n N_Y_M10_s N_Y_c_78_n N_Y_c_89_n N_Y_c_66_n N_Y_c_90_n
+ N_Y_c_91_n N_Y_c_67_n N_Y_c_69_n N_Y_c_99_p N_Y_c_71_n N_Y_c_73_n N_Y_c_95_n
+ N_Y_c_76_n N_Y_c_96_n N_Y_c_97_n N_Y_c_98_n N_Y_c_79_n N_Y_c_101_p N_Y_c_81_n
+ Y VSS PM_OAI222XP33_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00372052f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_13_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p A2 0.00477924f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.119
cc_4 N_A1_M0_g N_B2_M2_g 2.74891e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 VSS N_A1_M0_g 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_6 N_A1_c_3_p N_Y_c_65_n 0.00141058f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.119
cc_7 N_A1_c_3_p N_Y_c_66_n 0.00311007f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_8 N_A1_M0_g N_Y_c_67_n 2.68514e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_9 N_A1_c_3_p N_Y_c_67_n 0.00121543f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_10 N_A1_M0_g N_Y_c_69_n 2.64276e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_11 N_A1_c_3_p N_Y_c_69_n 0.00124805f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_12 N_A2_M1_g N_B2_M2_g 0.00335739f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_13 N_A2_c_13_n N_B2_c_25_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 A2 N_B2_c_26_n 0.00406615f $X=0.135 $Y=0.119 $X2=0.081 $Y2=0.135
cc_15 N_A2_M1_g N_B1_M3_g 2.74891e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 VSS N_A2_M1_g 3.47199e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_17 VSS A2 5.30079e-19 $X=0.135 $Y=0.119 $X2=0 $Y2=0
cc_18 N_A2_M1_g N_Y_c_71_n 2.56935e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 A2 N_Y_c_71_n 0.00123064f $X=0.135 $Y=0.119 $X2=0 $Y2=0
cc_20 N_B2_M2_g N_B1_M3_g 0.00372052f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_21 N_B2_c_25_n N_B1_c_36_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 N_B2_c_26_n B1 0.00477924f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 VSS N_B2_M2_g 3.57119e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 VSS N_B2_c_26_n 5.37372e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_25 N_B2_M2_g N_Y_c_73_n 2.56935e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_B2_c_26_n N_Y_c_73_n 0.00123064f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_27 B1 N_C1_c_45_n 5.26533e-19 $X=0.243 $Y=0.115 $X2=0 $Y2=0
cc_28 VSS N_B1_M3_g 2.08515e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_29 VSS N_B1_M3_g 2.76185e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_30 VSS B1 0.0012322f $X=0.243 $Y=0.115 $X2=0 $Y2=0
cc_31 B1 N_Y_c_75_n 0.00153032f $X=0.243 $Y=0.115 $X2=0.135 $Y2=0.135
cc_32 N_B1_M3_g N_Y_c_76_n 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_33 B1 N_Y_c_76_n 0.00124805f $X=0.243 $Y=0.115 $X2=0 $Y2=0
cc_34 N_C1_M4_g N_C2_M5_g 0.00347357f $X=0.405 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_35 N_C1_c_47_p N_C2_c_57_n 9.79748e-19 $X=0.405 $Y=0.135 $X2=0.243 $Y2=0.135
cc_36 C1 N_C2_c_58_n 0.00575328f $X=0.405 $Y=0.094 $X2=0.243 $Y2=0.115
cc_37 VSS C1 4.64783e-19 $X=0.405 $Y=0.094 $X2=0 $Y2=0
cc_38 VSS C1 0.00112518f $X=0.405 $Y=0.094 $X2=0 $Y2=0
cc_39 VSS N_C1_M4_g 2.64276e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_40 VSS C1 0.00125352f $X=0.405 $Y=0.094 $X2=0 $Y2=0
cc_41 N_C1_c_53_p N_Y_c_78_n 0.00153032f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_42 N_C1_M4_g N_Y_c_79_n 2.64276e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_C1_c_53_p N_Y_c_79_n 0.00125352f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_44 VSS N_C2_M5_g 2.7596e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_45 VSS N_C2_c_58_n 0.00125352f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_46 VSS N_C2_c_58_n 0.00114532f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_47 N_C2_M5_g N_Y_c_81_n 2.64276e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_48 N_C2_c_58_n N_Y_c_81_n 0.00125352f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_49 N_C2_c_58_n Y 0.00496438f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_50 VSS N_Y_c_84_n 0.00359992f $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.135
cc_51 VSS N_Y_c_84_n 0.00333673f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_52 VSS N_Y_c_84_n 0.00250965f $X=0.122 $Y=0.036 $X2=0.081 $Y2=0.135
cc_53 VSS N_Y_c_65_n 0.00138157f $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.135
cc_54 VSS N_Y_c_75_n 0.00138157f $X=0.27 $Y=0.036 $X2=0.081 $Y2=0.194
cc_55 VSS N_Y_c_89_n 3.56073e-19 $X=0.054 $Y=0.036 $X2=0 $Y2=0
cc_56 VSS N_Y_c_90_n 4.46493e-19 $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_57 VSS N_Y_c_91_n 2.63376e-19 $X=0.071 $Y=0.0675 $X2=0 $Y2=0
cc_58 VSS N_Y_c_91_n 0.00256253f $X=0.054 $Y=0.036 $X2=0 $Y2=0
cc_59 VSS N_Y_c_91_n 0.00707171f $X=0.122 $Y=0.036 $X2=0 $Y2=0
cc_60 VSS N_Y_c_90_n 2.90501e-19 $X=0.234 $Y=0.072 $X2=0 $Y2=0
cc_61 VSS N_Y_c_95_n 8.02788e-19 $X=0.234 $Y=0.072 $X2=0 $Y2=0
cc_62 VSS N_Y_c_96_n 8.02788e-19 $X=0.313 $Y=0.072 $X2=0 $Y2=0
cc_63 VSS N_Y_c_97_n 2.14558e-19 $X=0.396 $Y=0.036 $X2=0 $Y2=0
cc_64 VSS N_Y_c_98_n 2.14558e-19 $X=0.432 $Y=0.036 $X2=0 $Y2=0
cc_65 VSS N_Y_c_99_p 3.16424e-19 $X=0.122 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_66 VSS N_Y_c_95_n 3.16424e-19 $X=0.234 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_67 VSS N_Y_c_101_p 3.56327e-19 $X=0.45 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./OAI222xp33_ASAP7_75t_L.pex.sp.OAI222XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI22x1_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:54:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI22x1_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI22x1_ASAP7_75t_L.pex.sp.pex"
* File: OAI22x1_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:54:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI22X1_ASAP7_75T_L%B2 2 5 7 10 13 15 20 25 27 28 29 30 32 34 VSS
c32 40 VSS 1.80714e-19 $X=0.24 $Y=0.18
c33 34 VSS 2.04312e-19 $X=0.24 $Y=0.135
c34 32 VSS 1.70674e-19 $X=0.24 $Y=0.189
c35 31 VSS 5.67196e-19 $X=0.213 $Y=0.198
c36 30 VSS 0.00158425f $X=0.195 $Y=0.198
c37 29 VSS 0.00207482f $X=0.158 $Y=0.198
c38 28 VSS 1.5733e-19 $X=0.106 $Y=0.198
c39 27 VSS 4.68273e-20 $X=0.087 $Y=0.198
c40 26 VSS 1.94766e-19 $X=0.231 $Y=0.198
c41 25 VSS 3.54309e-19 $X=0.078 $Y=0.171
c42 20 VSS 0.00335953f $X=0.078 $Y=0.118
c43 18 VSS 3.51388e-19 $X=0.078 $Y=0.189
c44 13 VSS 9.94291e-19 $X=0.24 $Y=0.135
c45 10 VSS 0.0596118f $X=0.24 $Y=0.0675
c46 5 VSS 0.00251826f $X=0.078 $Y=0.135
c47 2 VSS 0.0640836f $X=0.078 $Y=0.0675
r48 39 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.24
+ $Y=0.171 $X2=0.24 $Y2=0.18
r49 34 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.24
+ $Y=0.135 $X2=0.24 $Y2=0.171
r50 32 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.24
+ $Y=0.189 $X2=0.24 $Y2=0.18
r51 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.195
+ $Y=0.198 $X2=0.213 $Y2=0.198
r52 29 30 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.158
+ $Y=0.198 $X2=0.195 $Y2=0.198
r53 28 29 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.106
+ $Y=0.198 $X2=0.158 $Y2=0.198
r54 27 28 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.087
+ $Y=0.198 $X2=0.106 $Y2=0.198
r55 26 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.231 $Y=0.198 $X2=0.24 $Y2=0.189
r56 26 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.231
+ $Y=0.198 $X2=0.213 $Y2=0.198
r57 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.153 $X2=0.078 $Y2=0.171
r58 22 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.135 $X2=0.078 $Y2=0.153
r59 20 22 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.118 $X2=0.078 $Y2=0.135
r60 18 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.078 $Y=0.189 $X2=0.087 $Y2=0.198
r61 18 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.189 $X2=0.078 $Y2=0.171
r62 13 34 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.24 $Y=0.135 $X2=0.24
+ $Y2=0.135
r63 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.24
+ $Y=0.135 $X2=0.24 $Y2=0.2025
r64 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.24
+ $Y=0.0675 $X2=0.24 $Y2=0.135
r65 5 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.078 $Y=0.135 $X2=0.078
+ $Y2=0.135
r66 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.078
+ $Y=0.135 $X2=0.078 $Y2=0.2025
r67 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.078
+ $Y=0.0675 $X2=0.078 $Y2=0.135
.ends

.subckt PM_OAI22X1_ASAP7_75T_L%B1 2 7 10 13 15 20 24 27 VSS
c24 27 VSS 1.30273e-19 $X=0.186 $Y=0.1255
c25 24 VSS 0.00136973f $X=0.186 $Y=0.135
c26 20 VSS 0.00274692f $X=0.18 $Y=0.108
c27 13 VSS 0.00532127f $X=0.186 $Y=0.135
c28 10 VSS 0.0613446f $X=0.186 $Y=0.0675
c29 2 VSS 0.0619872f $X=0.132 $Y=0.0675
r30 26 27 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.186
+ $Y=0.116 $X2=0.186 $Y2=0.1255
r31 24 27 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.186
+ $Y=0.135 $X2=0.186 $Y2=0.1255
r32 20 26 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.186
+ $Y=0.108 $X2=0.186 $Y2=0.116
r33 13 24 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.186 $Y=0.135 $X2=0.186
+ $Y2=0.135
r34 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.186
+ $Y=0.135 $X2=0.186 $Y2=0.2025
r35 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.186
+ $Y=0.0675 $X2=0.186 $Y2=0.135
r36 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.132
+ $Y=0.135 $X2=0.186 $Y2=0.135
r37 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.132
+ $Y=0.135 $X2=0.132 $Y2=0.2025
r38 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.132
+ $Y=0.0675 $X2=0.132 $Y2=0.135
.ends

.subckt PM_OAI22X1_ASAP7_75T_L%A2 2 5 7 10 13 15 17 19 23 27 28 29 33 36 38 VSS
c36 36 VSS 2.00449e-19 $X=0.456 $Y=0.171
c37 33 VSS 7.84621e-19 $X=0.456 $Y=0.135
c38 31 VSS 3.51388e-19 $X=0.456 $Y=0.189
c39 29 VSS 0.00192557f $X=0.428 $Y=0.198
c40 28 VSS 0.00158425f $X=0.376 $Y=0.198
c41 27 VSS 3.27558e-19 $X=0.339 $Y=0.198
c42 26 VSS 2.02211e-20 $X=0.306 $Y=0.198
c43 24 VSS 1.49134e-19 $X=0.447 $Y=0.198
c44 23 VSS 1.80714e-19 $X=0.294 $Y=0.18
c45 19 VSS 1.97602e-19 $X=0.294 $Y=0.135
c46 17 VSS 2.17415e-19 $X=0.294 $Y=0.189
c47 13 VSS 0.00128452f $X=0.456 $Y=0.135
c48 10 VSS 0.065901f $X=0.456 $Y=0.0675
c49 5 VSS 0.00150858f $X=0.294 $Y=0.135
c50 2 VSS 0.0607338f $X=0.294 $Y=0.0675
r51 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.456
+ $Y=0.153 $X2=0.456 $Y2=0.171
r52 33 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.456
+ $Y=0.135 $X2=0.456 $Y2=0.153
r53 31 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.456
+ $Y=0.189 $X2=0.456 $Y2=0.171
r54 28 29 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.376
+ $Y=0.198 $X2=0.428 $Y2=0.198
r55 27 28 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.339
+ $Y=0.198 $X2=0.376 $Y2=0.198
r56 26 27 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.198 $X2=0.339 $Y2=0.198
r57 25 38 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.303
+ $Y=0.198 $X2=0.294 $Y2=0.198
r58 25 26 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.303
+ $Y=0.198 $X2=0.306 $Y2=0.198
r59 24 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.447 $Y=0.198 $X2=0.456 $Y2=0.189
r60 24 29 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.198 $X2=0.428 $Y2=0.198
r61 22 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.294
+ $Y=0.171 $X2=0.294 $Y2=0.18
r62 19 22 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.294
+ $Y=0.135 $X2=0.294 $Y2=0.171
r63 17 38 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.294
+ $Y=0.189 $X2=0.294 $Y2=0.198
r64 17 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.294
+ $Y=0.189 $X2=0.294 $Y2=0.18
r65 13 33 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.456 $Y=0.135 $X2=0.456
+ $Y2=0.135
r66 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.456
+ $Y=0.135 $X2=0.456 $Y2=0.2025
r67 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.456
+ $Y=0.0675 $X2=0.456 $Y2=0.135
r68 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.294 $Y=0.135 $X2=0.294
+ $Y2=0.135
r69 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.294
+ $Y=0.135 $X2=0.294 $Y2=0.2025
r70 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.294
+ $Y=0.0675 $X2=0.294 $Y2=0.135
.ends

.subckt PM_OAI22X1_ASAP7_75T_L%A1 2 7 10 13 15 18 20 30 VSS
c26 20 VSS 6.50194e-19 $X=0.348 $Y=0.135
c27 18 VSS 0.00119149f $X=0.348 $Y=0.153
c28 13 VSS 0.00513876f $X=0.402 $Y=0.135
c29 10 VSS 0.0637989f $X=0.402 $Y=0.0675
c30 2 VSS 0.0626674f $X=0.348 $Y=0.0675
r31 18 30 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.348
+ $Y=0.1575 $X2=0.356 $Y2=0.1575
r32 18 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.348
+ $Y=0.153 $X2=0.348 $Y2=0.135
r33 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.402
+ $Y=0.135 $X2=0.402 $Y2=0.2025
r34 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.402
+ $Y=0.0675 $X2=0.402 $Y2=0.135
r35 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.348
+ $Y=0.135 $X2=0.402 $Y2=0.135
r36 5 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.348 $Y=0.135 $X2=0.348
+ $Y2=0.135
r37 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.348
+ $Y=0.135 $X2=0.348 $Y2=0.2025
r38 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.348
+ $Y=0.0675 $X2=0.348 $Y2=0.135
.ends

.subckt PM_OAI22X1_ASAP7_75T_L%Y 1 2 5 6 7 10 11 14 16 17 20 21 24 37 42 51 52
+ 53 55 56 60 62 VSS
c47 64 VSS 4.55454e-19 $X=0.51 $Y=0.216
c48 62 VSS 0.00123172f $X=0.51 $Y=0.1275
c49 61 VSS 8.85605e-19 $X=0.51 $Y=0.099
c50 60 VSS 0.00333801f $X=0.51 $Y=0.156
c51 58 VSS 4.30151e-19 $X=0.51 $Y=0.225
c52 56 VSS 3.46932e-19 $X=0.497 $Y=0.072
c53 55 VSS 8.46035e-21 $X=0.465 $Y=0.072
c54 53 VSS 3.69675e-19 $X=0.428 $Y=0.072
c55 52 VSS 5.76352e-20 $X=0.376 $Y=0.072
c56 51 VSS 5.76656e-19 $X=0.339 $Y=0.072
c57 43 VSS 0.0021974f $X=0.501 $Y=0.072
c58 42 VSS 0.0176071f $X=0.465 $Y=0.234
c59 41 VSS 0.00359728f $X=0.285 $Y=0.234
c60 37 VSS 0.0176042f $X=0.249 $Y=0.234
c61 36 VSS 0.00257895f $X=0.069 $Y=0.234
c62 28 VSS 0.00223184f $X=0.051 $Y=0.234
c63 26 VSS 0.00709337f $X=0.501 $Y=0.234
c64 24 VSS 0.00381938f $X=0.481 $Y=0.2025
c65 20 VSS 0.00480088f $X=0.267 $Y=0.2025
c66 16 VSS 5.38922e-19 $X=0.284 $Y=0.2025
c67 14 VSS 0.00359039f $X=0.053 $Y=0.2025
c68 11 VSS 2.69461e-19 $X=0.068 $Y=0.2025
c69 10 VSS 0.00215645f $X=0.429 $Y=0.0675
c70 6 VSS 7.35996e-19 $X=0.446 $Y=0.0675
c71 5 VSS 0.0025205f $X=0.321 $Y=0.0675
c72 1 VSS 6.53507e-19 $X=0.338 $Y=0.0675
r73 63 64 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.51
+ $Y=0.207 $X2=0.51 $Y2=0.216
r74 61 62 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.51
+ $Y=0.099 $X2=0.51 $Y2=0.1275
r75 60 63 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.51
+ $Y=0.156 $X2=0.51 $Y2=0.207
r76 60 62 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.51
+ $Y=0.156 $X2=0.51 $Y2=0.1275
r77 58 64 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.51
+ $Y=0.225 $X2=0.51 $Y2=0.216
r78 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.51
+ $Y=0.081 $X2=0.51 $Y2=0.099
r79 55 56 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.465
+ $Y=0.072 $X2=0.497 $Y2=0.072
r80 53 54 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.428
+ $Y=0.072 $X2=0.4285 $Y2=0.072
r81 52 53 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.376
+ $Y=0.072 $X2=0.428 $Y2=0.072
r82 51 52 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.339
+ $Y=0.072 $X2=0.376 $Y2=0.072
r83 49 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.429
+ $Y=0.072 $X2=0.465 $Y2=0.072
r84 49 54 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.429
+ $Y=0.072 $X2=0.4285 $Y2=0.072
r85 45 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.321
+ $Y=0.072 $X2=0.339 $Y2=0.072
r86 43 57 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.501 $Y=0.072 $X2=0.51 $Y2=0.081
r87 43 56 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.501
+ $Y=0.072 $X2=0.497 $Y2=0.072
r88 41 42 12.2222 $w=1.8e-08 $l=1.8e-07 $layer=M1 $thickness=3.6e-08 $X=0.285
+ $Y=0.234 $X2=0.465 $Y2=0.234
r89 39 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.483
+ $Y=0.234 $X2=0.465 $Y2=0.234
r90 36 37 12.2222 $w=1.8e-08 $l=1.8e-07 $layer=M1 $thickness=3.6e-08 $X=0.069
+ $Y=0.234 $X2=0.249 $Y2=0.234
r91 34 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.267
+ $Y=0.234 $X2=0.285 $Y2=0.234
r92 34 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.267
+ $Y=0.234 $X2=0.249 $Y2=0.234
r93 28 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.051
+ $Y=0.234 $X2=0.069 $Y2=0.234
r94 26 58 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.501 $Y=0.234 $X2=0.51 $Y2=0.225
r95 26 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.501
+ $Y=0.234 $X2=0.483 $Y2=0.234
r96 24 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.483 $Y=0.234 $X2=0.483
+ $Y2=0.234
r97 21 24 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.466 $Y=0.2025 $X2=0.481 $Y2=0.2025
r98 20 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.267 $Y=0.234 $X2=0.267
+ $Y2=0.234
r99 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.25 $Y=0.2025 $X2=0.267 $Y2=0.2025
r100 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.284 $Y=0.2025 $X2=0.267 $Y2=0.2025
r101 14 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.051 $Y=0.234
+ $X2=0.051 $Y2=0.234
r102 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.068 $Y=0.2025 $X2=0.053 $Y2=0.2025
r103 10 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.429 $Y=0.072
+ $X2=0.429 $Y2=0.072
r104 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.412 $Y=0.0675 $X2=0.429 $Y2=0.0675
r105 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.446 $Y=0.0675 $X2=0.429 $Y2=0.0675
r106 5 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.321 $Y=0.072 $X2=0.321
+ $Y2=0.072
r107 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.304 $Y=0.0675 $X2=0.321 $Y2=0.0675
r108 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.338 $Y=0.0675 $X2=0.321 $Y2=0.0675
.ends


* END of "./OAI22x1_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI22x1_ASAP7_75t_L  VSS VDD B2 B1 A2 A1 Y
* 
* Y	Y
* A1	A1
* A2	A2
* B1	B1
* B2	B2
M0 VSS N_B2_M0_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.068
+ $Y=0.027
M1 noxref_7 N_B1_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.122
+ $Y=0.027
M2 noxref_7 N_B1_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.176
+ $Y=0.027
M3 VSS N_B2_M3_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.23 $Y=0.027
M4 N_Y_M4_d N_A2_M4_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.284
+ $Y=0.027
M5 noxref_7 N_A1_M5_g N_Y_M5_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.338
+ $Y=0.027
M6 noxref_7 N_A1_M6_g N_Y_M6_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.392
+ $Y=0.027
M7 N_Y_M7_d N_A2_M7_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.446
+ $Y=0.027
M8 N_Y_M8_d N_B2_M8_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.068
+ $Y=0.162
M9 noxref_9 N_B1_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.122
+ $Y=0.162
M10 noxref_10 N_B1_M10_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.176
+ $Y=0.162
M11 N_Y_M11_d N_B2_M11_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.23
+ $Y=0.162
M12 N_Y_M12_d N_A2_M12_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.284 $Y=0.162
M13 noxref_11 N_A1_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.338
+ $Y=0.162
M14 noxref_12 N_A1_M14_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.392
+ $Y=0.162
M15 N_Y_M15_d N_A2_M15_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.446 $Y=0.162
*
* 
* .include "OAI22x1_ASAP7_75t_L.pex.sp.OAI22X1_ASAP7_75T_L.pxi"
* BEGIN of "./OAI22x1_ASAP7_75t_L.pex.sp.OAI22X1_ASAP7_75T_L.pxi"
* File: OAI22x1_ASAP7_75t_L.pex.sp.OAI22X1_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:54:25 2017
* 
x_PM_OAI22X1_ASAP7_75T_L%B2 N_B2_M0_g N_B2_c_7_p N_B2_M8_g N_B2_M3_g N_B2_c_8_p
+ N_B2_M11_g B2 N_B2_c_11_p N_B2_c_32_p N_B2_c_24_p N_B2_c_3_p N_B2_c_6_p
+ N_B2_c_17_p N_B2_c_13_p VSS PM_OAI22X1_ASAP7_75T_L%B2
x_PM_OAI22X1_ASAP7_75T_L%B1 N_B1_M1_g N_B1_M9_g N_B1_M2_g N_B1_c_39_n N_B1_M10_g
+ B1 N_B1_c_43_n N_B1_c_46_n VSS PM_OAI22X1_ASAP7_75T_L%B1
x_PM_OAI22X1_ASAP7_75T_L%A2 N_A2_M4_g N_A2_c_58_n N_A2_M12_g N_A2_M7_g
+ N_A2_c_70_p N_A2_M15_g N_A2_c_59_n N_A2_c_60_n N_A2_c_61_n N_A2_c_86_p
+ N_A2_c_65_p N_A2_c_68_p N_A2_c_75_p N_A2_c_73_p A2 VSS
+ PM_OAI22X1_ASAP7_75T_L%A2
x_PM_OAI22X1_ASAP7_75T_L%A1 N_A1_M5_g N_A1_M13_g N_A1_M6_g N_A1_c_100_n
+ N_A1_M14_g N_A1_c_103_n N_A1_c_105_n A1 VSS PM_OAI22X1_ASAP7_75T_L%A1
x_PM_OAI22X1_ASAP7_75T_L%Y N_Y_M5_s N_Y_M4_d N_Y_c_138_n N_Y_M7_d N_Y_M6_s
+ N_Y_c_126_n N_Y_M8_d N_Y_c_119_n N_Y_M12_d N_Y_M11_d N_Y_c_120_n N_Y_M15_d
+ N_Y_c_128_n N_Y_c_121_n N_Y_c_129_n N_Y_c_132_n N_Y_c_141_n N_Y_c_133_n
+ N_Y_c_134_n N_Y_c_159_n Y N_Y_c_137_n VSS PM_OAI22X1_ASAP7_75T_L%Y
cc_1 N_B2_M0_g N_B1_M1_g 0.00315405f $X=0.078 $Y=0.0675 $X2=0.132 $Y2=0.0675
cc_2 N_B2_M3_g N_B1_M1_g 2.25374e-19 $X=0.24 $Y=0.0675 $X2=0.132 $Y2=0.0675
cc_3 N_B2_c_3_p N_B1_M1_g 3.97719e-19 $X=0.158 $Y=0.198 $X2=0.132 $Y2=0.0675
cc_4 N_B2_M0_g N_B1_M2_g 2.25374e-19 $X=0.078 $Y=0.0675 $X2=0.186 $Y2=0.0675
cc_5 N_B2_M3_g N_B1_M2_g 0.00315405f $X=0.24 $Y=0.0675 $X2=0.186 $Y2=0.0675
cc_6 N_B2_c_6_p N_B1_M2_g 2.52885e-19 $X=0.195 $Y=0.198 $X2=0.186 $Y2=0.0675
cc_7 N_B2_c_7_p N_B1_c_39_n 0.00130109f $X=0.078 $Y=0.135 $X2=0.186 $Y2=0.135
cc_8 N_B2_c_8_p N_B1_c_39_n 9.59209e-19 $X=0.24 $Y=0.135 $X2=0.186 $Y2=0.135
cc_9 N_B2_c_3_p N_B1_c_39_n 7.25985e-19 $X=0.158 $Y=0.198 $X2=0.186 $Y2=0.135
cc_10 B2 B1 0.00124427f $X=0.078 $Y=0.118 $X2=0.18 $Y2=0.108
cc_11 N_B2_c_11_p N_B1_c_43_n 4.40275e-19 $X=0.078 $Y=0.171 $X2=0.186 $Y2=0.135
cc_12 N_B2_c_6_p N_B1_c_43_n 0.00373189f $X=0.195 $Y=0.198 $X2=0.186 $Y2=0.135
cc_13 N_B2_c_13_p N_B1_c_43_n 0.00165391f $X=0.24 $Y=0.135 $X2=0.186 $Y2=0.135
cc_14 N_B2_c_13_p N_B1_c_46_n 8.26953e-19 $X=0.24 $Y=0.135 $X2=0.186 $Y2=0.1255
cc_15 N_B2_M3_g N_A2_M4_g 0.00353901f $X=0.24 $Y=0.0675 $X2=0.132 $Y2=0.0675
cc_16 N_B2_c_8_p N_A2_c_58_n 8.87978e-19 $X=0.24 $Y=0.135 $X2=0.132 $Y2=0.135
cc_17 N_B2_c_17_p N_A2_c_59_n 0.00127963f $X=0.24 $Y=0.189 $X2=0 $Y2=0
cc_18 N_B2_c_13_p N_A2_c_60_n 0.00127963f $X=0.24 $Y=0.135 $X2=0.186 $Y2=0.108
cc_19 N_B2_c_13_p N_A2_c_61_n 0.00127963f $X=0.24 $Y=0.135 $X2=0.186 $Y2=0.135
cc_20 N_B2_M3_g N_A1_M5_g 2.949e-19 $X=0.24 $Y=0.0675 $X2=0.132 $Y2=0.0675
cc_21 VSS B2 8.25153e-19 $X=0.078 $Y=0.118 $X2=0 $Y2=0
cc_22 VSS N_B2_M0_g 2.38303e-19 $X=0.078 $Y=0.0675 $X2=0.186 $Y2=0.135
cc_23 VSS B2 0.00377207f $X=0.078 $Y=0.118 $X2=0.186 $Y2=0.135
cc_24 VSS N_B2_c_24_p 2.48779e-19 $X=0.106 $Y=0.198 $X2=0 $Y2=0
cc_25 VSS N_B2_c_3_p 2.48779e-19 $X=0.158 $Y=0.198 $X2=0 $Y2=0
cc_26 VSS N_B2_M3_g 3.62717e-19 $X=0.24 $Y=0.0675 $X2=0 $Y2=0
cc_27 VSS N_B2_c_13_p 4.46831e-19 $X=0.24 $Y=0.135 $X2=0 $Y2=0
cc_28 N_B2_c_11_p N_Y_c_119_n 0.0010499f $X=0.078 $Y=0.171 $X2=0.186 $Y2=0.2025
cc_29 N_B2_c_13_p N_Y_c_120_n 0.00158846f $X=0.24 $Y=0.135 $X2=0.18 $Y2=0.108
cc_30 N_B2_M0_g N_Y_c_121_n 2.38303e-19 $X=0.078 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_B2_M3_g N_Y_c_121_n 2.38303e-19 $X=0.24 $Y=0.0675 $X2=0 $Y2=0
cc_32 N_B2_c_32_p N_Y_c_121_n 0.016433f $X=0.087 $Y=0.198 $X2=0 $Y2=0
cc_33 N_B1_M2_g N_A2_M4_g 2.60137e-19 $X=0.186 $Y=0.0675 $X2=0.078 $Y2=0.0675
cc_34 VSS N_B1_c_39_n 3.80455e-19 $X=0.186 $Y=0.135 $X2=0.078 $Y2=0.2025
cc_35 VSS N_B1_c_39_n 8.00061e-19 $X=0.186 $Y=0.135 $X2=0.24 $Y2=0.189
cc_36 VSS B1 0.002048f $X=0.18 $Y=0.108 $X2=0.24 $Y2=0.189
cc_37 VSS N_B1_M1_g 4.62717e-19 $X=0.132 $Y=0.0675 $X2=0.24 $Y2=0.135
cc_38 VSS N_B1_c_39_n 3.50613e-19 $X=0.186 $Y=0.135 $X2=0.24 $Y2=0.135
cc_39 VSS N_B1_M2_g 2.34993e-19 $X=0.186 $Y=0.0675 $X2=0.24 $Y2=0.18
cc_40 VSS B1 0.00368948f $X=0.18 $Y=0.108 $X2=0.24 $Y2=0.18
cc_41 N_B1_M1_g N_Y_c_121_n 2.64781e-19 $X=0.132 $Y=0.0675 $X2=0 $Y2=0
cc_42 N_B1_M2_g N_Y_c_121_n 2.38303e-19 $X=0.186 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_A2_M4_g N_A1_M5_g 0.00358983f $X=0.294 $Y=0.0675 $X2=0.078 $Y2=0.0675
cc_44 N_A2_M7_g N_A1_M5_g 2.6588e-19 $X=0.456 $Y=0.0675 $X2=0.078 $Y2=0.0675
cc_45 N_A2_c_65_p N_A1_M5_g 2.52885e-19 $X=0.376 $Y=0.198 $X2=0.078 $Y2=0.0675
cc_46 N_A2_M4_g N_A1_M6_g 2.6588e-19 $X=0.294 $Y=0.0675 $X2=0.24 $Y2=0.0675
cc_47 N_A2_M7_g N_A1_M6_g 0.00364065f $X=0.456 $Y=0.0675 $X2=0.24 $Y2=0.0675
cc_48 N_A2_c_68_p N_A1_M6_g 3.99641e-19 $X=0.428 $Y=0.198 $X2=0.24 $Y2=0.0675
cc_49 N_A2_c_58_n N_A1_c_100_n 9.81317e-19 $X=0.294 $Y=0.135 $X2=0.24 $Y2=0.135
cc_50 N_A2_c_70_p N_A1_c_100_n 0.00129593f $X=0.456 $Y=0.135 $X2=0.24 $Y2=0.135
cc_51 N_A2_c_68_p N_A1_c_100_n 6.92083e-19 $X=0.428 $Y=0.198 $X2=0.24 $Y2=0.135
cc_52 N_A2_c_65_p N_A1_c_103_n 0.00371882f $X=0.376 $Y=0.198 $X2=0.078 $Y2=0.189
cc_53 N_A2_c_73_p N_A1_c_103_n 4.25941e-19 $X=0.456 $Y=0.171 $X2=0.078 $Y2=0.189
cc_54 N_A2_c_60_n N_A1_c_105_n 0.00239031f $X=0.294 $Y=0.135 $X2=0.078 $Y2=0.118
cc_55 N_A2_c_75_p N_A1_c_105_n 0.00101781f $X=0.456 $Y=0.135 $X2=0.078 $Y2=0.118
cc_56 VSS N_A2_M4_g 3.75866e-19 $X=0.294 $Y=0.0675 $X2=0 $Y2=0
cc_57 VSS N_A2_c_60_n 4.38244e-19 $X=0.294 $Y=0.135 $X2=0 $Y2=0
cc_58 VSS N_A2_M7_g 2.38303e-19 $X=0.456 $Y=0.0675 $X2=0 $Y2=0
cc_59 VSS N_A2_c_75_p 2.73699e-19 $X=0.456 $Y=0.135 $X2=0 $Y2=0
cc_60 N_A2_c_75_p N_Y_c_126_n 0.0313705f $X=0.456 $Y=0.135 $X2=0.24 $Y2=0.0675
cc_61 N_A2_c_60_n N_Y_c_120_n 0.00158846f $X=0.294 $Y=0.135 $X2=0.078 $Y2=0.118
cc_62 N_A2_c_73_p N_Y_c_128_n 0.00158881f $X=0.456 $Y=0.171 $X2=0.078 $Y2=0.153
cc_63 N_A2_M4_g N_Y_c_129_n 2.38303e-19 $X=0.294 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_A2_M7_g N_Y_c_129_n 2.38303e-19 $X=0.456 $Y=0.0675 $X2=0 $Y2=0
cc_65 N_A2_c_59_n N_Y_c_129_n 0.0164209f $X=0.294 $Y=0.189 $X2=0 $Y2=0
cc_66 N_A2_c_86_p N_Y_c_132_n 3.65124e-19 $X=0.339 $Y=0.198 $X2=0 $Y2=0
cc_67 N_A2_c_68_p N_Y_c_133_n 3.65124e-19 $X=0.428 $Y=0.198 $X2=0 $Y2=0
cc_68 N_A2_M7_g N_Y_c_134_n 2.52885e-19 $X=0.456 $Y=0.0675 $X2=0 $Y2=0
cc_69 N_A2_c_75_p N_Y_c_134_n 0.00371986f $X=0.456 $Y=0.135 $X2=0 $Y2=0
cc_70 N_A2_c_73_p Y 0.00218788f $X=0.456 $Y=0.171 $X2=0 $Y2=0
cc_71 N_A2_c_75_p N_Y_c_137_n 0.00218788f $X=0.456 $Y=0.135 $X2=0 $Y2=0
cc_72 VSS N_A2_c_86_p 2.54007e-19 $X=0.339 $Y=0.198 $X2=0.078 $Y2=0.0675
cc_73 VSS N_A1_c_100_n 3.78279e-19 $X=0.402 $Y=0.135 $X2=0 $Y2=0
cc_74 VSS N_A1_c_100_n 8.00061e-19 $X=0.402 $Y=0.135 $X2=0 $Y2=0
cc_75 VSS N_A1_c_105_n 8.76024e-19 $X=0.348 $Y=0.135 $X2=0 $Y2=0
cc_76 VSS N_A1_M5_g 2.15135e-19 $X=0.348 $Y=0.0675 $X2=0 $Y2=0
cc_77 VSS N_A1_M6_g 2.64781e-19 $X=0.402 $Y=0.0675 $X2=0 $Y2=0
cc_78 N_A1_c_105_n N_Y_c_138_n 3.21662e-19 $X=0.348 $Y=0.135 $X2=0.078 $Y2=0.135
cc_79 N_A1_M5_g N_Y_c_129_n 2.38303e-19 $X=0.348 $Y=0.0675 $X2=0 $Y2=0
cc_80 N_A1_M6_g N_Y_c_129_n 2.64781e-19 $X=0.402 $Y=0.0675 $X2=0 $Y2=0
cc_81 N_A1_M5_g N_Y_c_141_n 2.56447e-19 $X=0.348 $Y=0.0675 $X2=0 $Y2=0
cc_82 N_A1_c_105_n N_Y_c_141_n 0.00373962f $X=0.348 $Y=0.135 $X2=0 $Y2=0
cc_83 N_A1_M6_g N_Y_c_133_n 3.99641e-19 $X=0.402 $Y=0.0675 $X2=0 $Y2=0
cc_84 N_A1_c_100_n N_Y_c_133_n 5.37025e-19 $X=0.402 $Y=0.135 $X2=0 $Y2=0
cc_85 VSS N_Y_c_138_n 0.00339475f $X=0.267 $Y=0.036 $X2=0.078 $Y2=0.135
cc_86 VSS N_Y_c_138_n 0.0036466f $X=0.375 $Y=0.036 $X2=0.078 $Y2=0.135
cc_87 VSS N_Y_c_138_n 0.00250965f $X=0.3405 $Y=0.036 $X2=0.078 $Y2=0.135
cc_88 VSS N_Y_c_126_n 0.00372512f $X=0.375 $Y=0.036 $X2=0.24 $Y2=0.0675
cc_89 VSS N_Y_c_126_n 0.00251378f $X=0.483 $Y=0.036 $X2=0.24 $Y2=0.0675
cc_90 VSS N_Y_c_126_n 0.00384465f $X=0.483 $Y=0.036 $X2=0.24 $Y2=0.0675
cc_91 VSS N_Y_c_119_n 0.00107252f $X=0.051 $Y=0.036 $X2=0.24 $Y2=0.2025
cc_92 VSS N_Y_c_120_n 0.00107252f $X=0.267 $Y=0.036 $X2=0.078 $Y2=0.118
cc_93 VSS N_Y_c_128_n 0.00138157f $X=0.483 $Y=0.036 $X2=0.078 $Y2=0.153
cc_94 VSS N_Y_c_132_n 5.00406e-19 $X=0.267 $Y=0.036 $X2=0 $Y2=0
cc_95 VSS N_Y_c_132_n 0.00796074f $X=0.3405 $Y=0.036 $X2=0 $Y2=0
cc_96 VSS N_Y_c_141_n 0.00128262f $X=0.375 $Y=0.036 $X2=0 $Y2=0
cc_97 VSS N_Y_c_133_n 0.00107804f $X=0.375 $Y=0.036 $X2=0 $Y2=0
cc_98 VSS N_Y_c_133_n 0.00796074f $X=0.483 $Y=0.036 $X2=0 $Y2=0
cc_99 VSS N_Y_c_159_n 2.47657e-19 $X=0.481 $Y=0.0675 $X2=0 $Y2=0
cc_100 VSS N_Y_c_159_n 0.00260156f $X=0.483 $Y=0.036 $X2=0 $Y2=0
cc_101 VSS N_Y_c_137_n 2.86097e-19 $X=0.483 $Y=0.036 $X2=0 $Y2=0
cc_102 VSS N_Y_c_121_n 2.27254e-19 $X=0.249 $Y=0.234 $X2=0.078 $Y2=0.0675
cc_103 VSS N_Y_c_121_n 2.21722e-19 $X=0.249 $Y=0.234 $X2=0.078 $Y2=0.0675
cc_104 VSS N_Y_c_129_n 2.27254e-19 $X=0.465 $Y=0.234 $X2=0.078 $Y2=0.0675
cc_105 VSS N_Y_c_129_n 2.27254e-19 $X=0.465 $Y=0.234 $X2=0.078 $Y2=0.0675

* END of "./OAI22x1_ASAP7_75t_L.pex.sp.OAI22X1_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI22xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:54:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI22xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI22xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI22xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:54:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI22XP33_ASAP7_75T_L%A1 2 5 7 13 VSS
c10 13 VSS 0.00108961f $X=0.081 $Y=0.137
c11 5 VSS 0.00171842f $X=0.081 $Y=0.135
c12 2 VSS 0.0655219f $X=0.081 $Y=0.054
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI22XP33_ASAP7_75T_L%A2 2 5 7 13 VSS
c12 13 VSS 7.1352e-19 $X=0.134 $Y=0.137
c13 5 VSS 0.00113686f $X=0.135 $Y=0.135
c14 2 VSS 0.0617048f $X=0.135 $Y=0.054
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI22XP33_ASAP7_75T_L%B2 2 5 7 15 VSS
c11 15 VSS 0.00249308f $X=0.189 $Y=0.138
c12 5 VSS 0.00123188f $X=0.189 $Y=0.135
c13 2 VSS 0.0612814f $X=0.189 $Y=0.054
r14 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI22XP33_ASAP7_75T_L%B1 2 5 7 14 VSS
c9 14 VSS 0.0119502f $X=0.242 $Y=0.138
c10 5 VSS 0.00227588f $X=0.243 $Y=0.135
c11 2 VSS 0.064914f $X=0.243 $Y=0.054
r12 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r13 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r14 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI22XP33_ASAP7_75T_L%Y 1 2 5 6 7 10 14 15 16 24 25 30 33 36 VSS
c20 37 VSS 9.61186e-19 $X=0.153 $Y=0.234
c21 36 VSS 0.00142296f $X=0.144 $Y=0.234
c22 35 VSS 9.49502e-19 $X=0.126 $Y=0.234
c23 34 VSS 0.0025752f $X=0.117 $Y=0.234
c24 33 VSS 0.00146362f $X=0.09 $Y=0.234
c25 32 VSS 0.00758013f $X=0.072 $Y=0.234
c26 30 VSS 0.00290871f $X=0.162 $Y=0.234
c27 28 VSS 0.00321443f $X=0.027 $Y=0.234
c28 26 VSS 1.49741e-19 $X=0.099 $Y=0.072
c29 25 VSS 8.46035e-21 $X=0.09 $Y=0.072
c30 24 VSS 5.00007e-19 $X=0.072 $Y=0.072
c31 23 VSS 9.77732e-19 $X=0.04 $Y=0.072
c32 21 VSS 4.62191e-19 $X=0.108 $Y=0.072
c33 19 VSS 0.00191766f $X=0.027 $Y=0.072
c34 18 VSS 7.00744e-19 $X=0.018 $Y=0.2125
c35 16 VSS 4.27371e-19 $X=0.018 $Y=0.115
c36 15 VSS 0.00112063f $X=0.018 $Y=0.106
c37 14 VSS 0.00410446f $X=0.02 $Y=0.124
c38 12 VSS 5.68738e-19 $X=0.018 $Y=0.225
c39 10 VSS 0.00410355f $X=0.162 $Y=0.216
c40 6 VSS 5.65078e-19 $X=0.179 $Y=0.216
c41 5 VSS 0.00282776f $X=0.108 $Y=0.054
c42 1 VSS 5.83614e-19 $X=0.125 $Y=0.054
r43 36 37 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.153 $Y2=0.234
r44 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r45 34 35 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.234 $X2=0.126 $Y2=0.234
r46 33 34 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.117 $Y2=0.234
r47 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r48 30 37 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.153 $Y2=0.234
r49 28 32 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.072 $Y2=0.234
r50 25 26 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.099 $Y2=0.072
r51 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.072 $X2=0.09 $Y2=0.072
r52 23 24 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.072 $X2=0.072 $Y2=0.072
r53 21 26 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.099 $Y2=0.072
r54 19 23 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.072 $X2=0.04 $Y2=0.072
r55 17 18 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r56 15 16 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.106 $X2=0.018 $Y2=0.115
r57 14 17 5.16049 $w=1.8e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.124 $X2=0.018 $Y2=0.2
r58 14 16 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.124 $X2=0.018 $Y2=0.115
r59 12 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r60 12 18 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r61 11 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.081 $X2=0.027 $Y2=0.072
r62 11 15 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.106
r63 10 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r64 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.162 $Y2=0.216
r65 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.216 $X2=0.162 $Y2=0.216
r66 5 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072 $X2=0.108
+ $Y2=0.072
r67 2 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.054 $X2=0.108 $Y2=0.054
r68 1 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.054 $X2=0.108 $Y2=0.054
.ends


* END of "./OAI22xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI22xp33_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 Y
* 
* Y	Y
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 N_Y_M0_d N_A1_M0_g noxref_8 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 noxref_8 N_A2_M1_g N_Y_M1_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 VSS N_B2_M2_g noxref_8 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.027
M3 noxref_8 N_B1_M3_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 noxref_9 N_A1_M4_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M5 N_Y_M5_d N_A2_M5_g noxref_9 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M6 noxref_10 N_B2_M6_g N_Y_M6_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M7 VDD N_B1_M7_g noxref_10 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
*
* 
* .include "OAI22xp33_ASAP7_75t_L.pex.sp.OAI22XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI22xp33_ASAP7_75t_L.pex.sp.OAI22XP33_ASAP7_75T_L.pxi"
* File: OAI22xp33_ASAP7_75t_L.pex.sp.OAI22XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:54:48 2017
* 
x_PM_OAI22XP33_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M4_g A1 VSS
+ PM_OAI22XP33_ASAP7_75T_L%A1
x_PM_OAI22XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_12_n N_A2_M5_g A2 VSS
+ PM_OAI22XP33_ASAP7_75T_L%A2
x_PM_OAI22XP33_ASAP7_75T_L%B2 N_B2_M2_g N_B2_c_25_n N_B2_M6_g B2 VSS
+ PM_OAI22XP33_ASAP7_75T_L%B2
x_PM_OAI22XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_36_n N_B1_M7_g B1 VSS
+ PM_OAI22XP33_ASAP7_75T_L%B1
x_PM_OAI22XP33_ASAP7_75T_L%Y N_Y_M1_s N_Y_M0_d N_Y_c_55_p N_Y_M6_s N_Y_M5_d
+ N_Y_c_48_n Y N_Y_c_56_p N_Y_c_43_n N_Y_c_54_p N_Y_c_44_n N_Y_c_53_n N_Y_c_46_n
+ N_Y_c_49_n VSS PM_OAI22XP33_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.0036697f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A1_c_2_p N_A2_c_12_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A1 A2 0.00484691f $X=0.081 $Y=0.137 $X2=0.134 $Y2=0.137
cc_4 N_A1_M0_g N_B2_M2_g 3.03912e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 A1 N_Y_c_43_n 0.00356618f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_6 N_A1_M0_g N_Y_c_44_n 2.68514e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_7 A1 N_Y_c_44_n 0.00121543f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_8 N_A1_M0_g N_Y_c_46_n 2.64276e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_9 A1 N_Y_c_46_n 0.00124805f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_10 VSS N_A1_M0_g 2.38303e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_11 N_A2_M1_g N_B2_M2_g 0.00361888f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_12 N_A2_c_12_n N_B2_c_25_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_13 A2 B2 0.00439547f $X=0.134 $Y=0.137 $X2=0 $Y2=0
cc_14 N_A2_M1_g N_B1_M3_g 2.69148e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_15 A2 N_Y_c_48_n 3.87865e-19 $X=0.134 $Y=0.137 $X2=0.081 $Y2=0.135
cc_16 N_A2_M1_g N_Y_c_49_n 2.56935e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_17 A2 N_Y_c_49_n 0.00123064f $X=0.134 $Y=0.137 $X2=0 $Y2=0
cc_18 VSS N_A2_M1_g 3.47199e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_19 VSS A2 5.30079e-19 $X=0.134 $Y=0.137 $X2=0 $Y2=0
cc_20 N_B2_M2_g N_B1_M3_g 0.00323392f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_21 N_B2_c_25_n N_B1_c_36_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 B2 B1 0.00565996f $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_23 B2 N_Y_c_48_n 3.87865e-19 $X=0.189 $Y=0.138 $X2=0.081 $Y2=0.135
cc_24 VSS B2 9.95856e-19 $X=0.189 $Y=0.138 $X2=0.081 $Y2=0.135
cc_25 VSS N_B2_M2_g 2.56935e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_26 VSS B2 0.00123604f $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_27 B1 N_Y_c_48_n 3.8851e-19 $X=0.242 $Y=0.138 $X2=0.135 $Y2=0.135
cc_28 B1 N_Y_c_53_n 7.09702e-19 $X=0.242 $Y=0.138 $X2=0 $Y2=0
cc_29 VSS B1 6.98375e-19 $X=0.242 $Y=0.138 $X2=0 $Y2=0
cc_30 VSS N_B1_M3_g 2.56935e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_31 VSS B1 0.00123969f $X=0.242 $Y=0.138 $X2=0 $Y2=0
cc_32 VSS N_Y_c_54_p 2.69772e-19 $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.054
cc_33 VSS N_Y_c_55_p 0.00359978f $X=0.108 $Y=0.054 $X2=0.081 $Y2=0.135
cc_34 VSS N_Y_c_56_p 2.98193e-19 $X=0.018 $Y=0.106 $X2=0.081 $Y2=0.135
cc_35 VSS N_Y_c_54_p 0.00255467f $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.135
cc_36 VSS N_Y_c_55_p 0.00356866f $X=0.108 $Y=0.054 $X2=0.081 $Y2=0.135
cc_37 VSS N_Y_c_48_n 9.28287e-19 $X=0.162 $Y=0.216 $X2=0.081 $Y2=0.135
cc_38 VSS N_Y_c_55_p 0.00189275f $X=0.108 $Y=0.054 $X2=0 $Y2=0
cc_39 VSS N_Y_c_54_p 0.00670034f $X=0.072 $Y=0.072 $X2=0 $Y2=0
cc_40 VSS N_Y_c_55_p 6.35113e-19 $X=0.108 $Y=0.054 $X2=0 $Y2=0

* END of "./OAI22xp33_ASAP7_75t_L.pex.sp.OAI22XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI22xp5_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:55:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI22xp5_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI22xp5_ASAP7_75t_L.pex.sp.pex"
* File: OAI22xp5_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:55:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI22XP5_ASAP7_75T_L%A1 2 5 7 13 VSS
c10 13 VSS 0.00178342f $X=0.081 $Y=0.137
c11 5 VSS 0.00171842f $X=0.081 $Y=0.135
c12 2 VSS 0.0655219f $X=0.081 $Y=0.0675
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI22XP5_ASAP7_75T_L%A2 2 5 7 14 VSS
c13 14 VSS 0.00122494f $X=0.134 $Y=0.137
c14 5 VSS 0.00110459f $X=0.135 $Y=0.135
c15 2 VSS 0.0618838f $X=0.135 $Y=0.0675
r16 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI22XP5_ASAP7_75T_L%B2 2 5 7 15 VSS
c11 15 VSS 0.00285149f $X=0.189 $Y=0.138
c12 5 VSS 0.00119608f $X=0.189 $Y=0.135
c13 2 VSS 0.0615532f $X=0.189 $Y=0.0675
r14 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI22XP5_ASAP7_75T_L%B1 2 5 7 14 VSS
c10 14 VSS 0.0127247f $X=0.242 $Y=0.138
c11 5 VSS 0.00227588f $X=0.243 $Y=0.135
c12 2 VSS 0.064914f $X=0.243 $Y=0.0675
r13 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI22XP5_ASAP7_75T_L%Y 1 2 5 6 7 10 14 15 16 21 24 25 30 33 34 VSS
c21 35 VSS 9.60848e-19 $X=0.126 $Y=0.234
c22 34 VSS 0.00242114f $X=0.117 $Y=0.234
c23 33 VSS 0.00146362f $X=0.09 $Y=0.234
c24 32 VSS 0.00797257f $X=0.072 $Y=0.234
c25 30 VSS 0.00471725f $X=0.162 $Y=0.234
c26 28 VSS 0.00321443f $X=0.027 $Y=0.234
c27 26 VSS 1.51286e-19 $X=0.099 $Y=0.072
c28 25 VSS 8.46035e-21 $X=0.09 $Y=0.072
c29 24 VSS 5.33412e-19 $X=0.072 $Y=0.072
c30 23 VSS 9.77732e-19 $X=0.04 $Y=0.072
c31 21 VSS 2.63908e-19 $X=0.108 $Y=0.072
c32 19 VSS 0.00191766f $X=0.027 $Y=0.072
c33 18 VSS 4.28499e-19 $X=0.018 $Y=0.207
c34 16 VSS 4.27371e-19 $X=0.018 $Y=0.115
c35 15 VSS 0.00112034f $X=0.018 $Y=0.106
c36 14 VSS 0.00402652f $X=0.02 $Y=0.124
c37 12 VSS 8.29409e-19 $X=0.018 $Y=0.225
c38 10 VSS 0.00485022f $X=0.162 $Y=0.2025
c39 6 VSS 6.12285e-19 $X=0.179 $Y=0.2025
c40 5 VSS 0.00256112f $X=0.108 $Y=0.0675
c41 1 VSS 6.7534e-19 $X=0.125 $Y=0.0675
r42 34 35 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.234 $X2=0.126 $Y2=0.234
r43 33 34 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.117 $Y2=0.234
r44 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r45 30 35 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.126 $Y2=0.234
r46 28 32 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.072 $Y2=0.234
r47 25 26 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.099 $Y2=0.072
r48 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.072 $X2=0.09 $Y2=0.072
r49 23 24 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.072 $X2=0.072 $Y2=0.072
r50 21 26 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.099 $Y2=0.072
r51 19 23 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.072 $X2=0.04 $Y2=0.072
r52 17 18 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.207
r53 15 16 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.106 $X2=0.018 $Y2=0.115
r54 14 17 5.16049 $w=1.8e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.124 $X2=0.018 $Y2=0.2
r55 14 16 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.124 $X2=0.018 $Y2=0.115
r56 12 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r57 12 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.207
r58 11 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.081 $X2=0.027 $Y2=0.072
r59 11 15 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.106
r60 10 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r61 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r62 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r63 5 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072 $X2=0.108
+ $Y2=0.072
r64 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r65 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./OAI22xp5_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI22xp5_ASAP7_75t_L  VSS VDD A1 A2 B2 B1 Y
* 
* Y	Y
* B1	B1
* B2	B2
* A2	A2
* A1	A1
M0 N_Y_M0_d N_A1_M0_g noxref_8 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_8 N_A2_M1_g N_Y_M1_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_B2_M2_g noxref_8 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_8 N_B1_M3_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_9 N_A1_M4_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 N_Y_M5_d N_A2_M5_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 noxref_10 N_B2_M6_g N_Y_M6_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M7 VDD N_B1_M7_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
*
* 
* .include "OAI22xp5_ASAP7_75t_L.pex.sp.OAI22XP5_ASAP7_75T_L.pxi"
* BEGIN of "./OAI22xp5_ASAP7_75t_L.pex.sp.OAI22XP5_ASAP7_75T_L.pxi"
* File: OAI22xp5_ASAP7_75t_L.pex.sp.OAI22XP5_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:55:10 2017
* 
x_PM_OAI22XP5_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M4_g A1 VSS
+ PM_OAI22XP5_ASAP7_75T_L%A1
x_PM_OAI22XP5_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_12_n N_A2_M5_g A2 VSS
+ PM_OAI22XP5_ASAP7_75T_L%A2
x_PM_OAI22XP5_ASAP7_75T_L%B2 N_B2_M2_g N_B2_c_26_n N_B2_M6_g B2 VSS
+ PM_OAI22XP5_ASAP7_75T_L%B2
x_PM_OAI22XP5_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_38_n N_B1_M7_g B1 VSS
+ PM_OAI22XP5_ASAP7_75T_L%B1
x_PM_OAI22XP5_ASAP7_75T_L%Y N_Y_M1_s N_Y_M0_d N_Y_c_57_p N_Y_M6_s N_Y_M5_d
+ N_Y_c_50_n Y N_Y_c_58_p N_Y_c_45_n N_Y_c_53_n N_Y_c_56_p N_Y_c_46_n N_Y_c_51_n
+ N_Y_c_48_n N_Y_c_65_p VSS PM_OAI22XP5_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.0036697f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A1_c_2_p N_A2_c_12_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A1 A2 0.00468131f $X=0.081 $Y=0.137 $X2=0.134 $Y2=0.137
cc_4 N_A1_M0_g N_B2_M2_g 3.03912e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 A1 N_Y_c_45_n 0.0031019f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_6 N_A1_M0_g N_Y_c_46_n 2.68514e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_7 A1 N_Y_c_46_n 0.00121543f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_8 N_A1_M0_g N_Y_c_48_n 2.64276e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_9 A1 N_Y_c_48_n 0.00124805f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_10 VSS N_A1_M0_g 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_11 N_A2_M1_g N_B2_M2_g 0.00361888f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_12 N_A2_c_12_n N_B2_c_26_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_13 A2 B2 0.00240077f $X=0.134 $Y=0.137 $X2=0 $Y2=0
cc_14 N_A2_M1_g N_B1_M3_g 2.69148e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_15 A2 B1 6.34014e-19 $X=0.134 $Y=0.137 $X2=0 $Y2=0
cc_16 A2 N_Y_c_50_n 0.00261703f $X=0.134 $Y=0.137 $X2=0.081 $Y2=0.135
cc_17 N_A2_M1_g N_Y_c_51_n 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_18 A2 N_Y_c_51_n 0.00404783f $X=0.134 $Y=0.137 $X2=0 $Y2=0
cc_19 VSS N_A2_M1_g 3.47199e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_20 VSS A2 5.3065e-19 $X=0.134 $Y=0.137 $X2=0 $Y2=0
cc_21 N_B2_M2_g N_B1_M3_g 0.00323392f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_22 N_B2_c_26_n N_B1_c_38_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 B2 B1 0.00385905f $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_24 B2 N_Y_c_53_n 6.89204e-19 $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_25 VSS B2 0.00233505f $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_26 VSS N_B2_M2_g 2.34993e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_27 VSS B2 0.00455569f $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_28 B1 N_Y_c_50_n 8.23902e-19 $X=0.242 $Y=0.138 $X2=0 $Y2=0
cc_29 B1 N_Y_c_51_n 7.09702e-19 $X=0.242 $Y=0.138 $X2=0 $Y2=0
cc_30 VSS B1 6.98375e-19 $X=0.242 $Y=0.138 $X2=0 $Y2=0
cc_31 VSS N_B1_M3_g 2.56935e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_32 VSS B1 0.00123969f $X=0.242 $Y=0.138 $X2=0 $Y2=0
cc_33 VSS N_Y_c_56_p 2.6846e-19 $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_34 VSS N_Y_c_57_p 0.00359978f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_35 VSS N_Y_c_58_p 2.98193e-19 $X=0.018 $Y=0.106 $X2=0 $Y2=0
cc_36 VSS N_Y_c_56_p 0.00255467f $X=0.072 $Y=0.072 $X2=0 $Y2=0
cc_37 VSS N_Y_c_57_p 0.00362239f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_38 VSS N_Y_c_50_n 0.00158656f $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_39 VSS N_Y_c_57_p 0.00189275f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_40 VSS N_Y_c_56_p 0.00678908f $X=0.072 $Y=0.072 $X2=0 $Y2=0
cc_41 VSS N_Y_c_57_p 6.35113e-19 $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_42 VSS N_Y_c_65_p 2.65006e-19 $X=0.117 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./OAI22xp5_ASAP7_75t_L.pex.sp.OAI22XP5_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI311xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:55:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI311xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI311xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI311xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:55:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI311XP33_ASAP7_75T_L%A3 2 5 7 17 VSS
c5 17 VSS 0.0181247f $X=0.08 $Y=0.136
c6 5 VSS 0.00275452f $X=0.081 $Y=0.135
c7 2 VSS 0.0643308f $X=0.081 $Y=0.0675
r8 5 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r9 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r10 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI311XP33_ASAP7_75T_L%A2 2 5 7 15 VSS
c12 15 VSS 0.00402403f $X=0.134 $Y=0.136
c13 5 VSS 0.00131688f $X=0.135 $Y=0.135
c14 2 VSS 0.059793f $X=0.135 $Y=0.0675
r15 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI311XP33_ASAP7_75T_L%A1 2 5 7 13 VSS
c13 13 VSS 0.0021029f $X=0.196 $Y=0.136
c14 5 VSS 0.00118479f $X=0.189 $Y=0.135
c15 2 VSS 0.060496f $X=0.189 $Y=0.0675
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI311XP33_ASAP7_75T_L%B1 2 5 7 13 VSS
c11 13 VSS 0.00135757f $X=0.247 $Y=0.134
c12 5 VSS 0.00123712f $X=0.243 $Y=0.135
c13 2 VSS 0.0620388f $X=0.243 $Y=0.0675
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI311XP33_ASAP7_75T_L%C1 2 5 7 10 VSS
c9 10 VSS 0.00137012f $X=0.297 $Y=0.134
c10 5 VSS 0.00179274f $X=0.297 $Y=0.135
c11 2 VSS 0.0660696f $X=0.297 $Y=0.0675
r12 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r13 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OAI311XP33_ASAP7_75T_L%Y 1 7 8 10 13 19 26 27 28 34 39 42 45 VSS
c14 45 VSS 0.00384059f $X=0.342 $Y=0.036
c15 44 VSS 0.00278493f $X=0.351 $Y=0.036
c16 42 VSS 0.00232427f $X=0.324 $Y=0.036
c17 39 VSS 0.00565612f $X=0.351 $Y=0.2
c18 38 VSS 0.00126f $X=0.351 $Y=0.07
c19 37 VSS 9.04094e-19 $X=0.351 $Y=0.225
c20 35 VSS 4.19362e-19 $X=0.31 $Y=0.234
c21 34 VSS 0.00142296f $X=0.306 $Y=0.234
c22 33 VSS 0.00632503f $X=0.288 $Y=0.234
c23 32 VSS 0.00100794f $X=0.252 $Y=0.234
c24 28 VSS 6.7196e-19 $X=0.241 $Y=0.234
c25 27 VSS 0.00434692f $X=0.234 $Y=0.234
c26 20 VSS 0.00657518f $X=0.342 $Y=0.234
c27 19 VSS 0.00474875f $X=0.216 $Y=0.2025
c28 13 VSS 0.00574947f $X=0.322 $Y=0.216
c29 9 VSS 5.36031e-19 $X=0.216 $Y=0.2245
c30 4 VSS 3.02808e-19 $X=0.322 $Y=0.0675
r31 45 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.3465 $Y2=0.036
r32 44 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.036 $X2=0.3465 $Y2=0.036
r33 41 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r34 41 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r35 38 39 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.07 $X2=0.351 $Y2=0.2
r36 37 39 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.2
r37 36 44 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.036
r38 36 38 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.07
r39 34 35 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.31 $Y2=0.234
r40 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r41 32 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.288 $Y2=0.234
r42 30 35 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.31 $Y2=0.234
r43 27 28 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.241 $Y2=0.234
r44 26 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.234 $X2=0.252 $Y2=0.234
r45 26 28 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.234 $X2=0.241 $Y2=0.234
r46 22 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.234 $Y2=0.234
r47 20 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.234 $X2=0.351 $Y2=0.225
r48 20 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.324 $Y2=0.234
r49 19 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r50 13 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r51 10 13 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.216 $X2=0.322 $Y2=0.216
r52 8 9 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.2245 $X2=0.216 $Y2=0.2245
r53 7 9 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2245 $X2=0.216 $Y2=0.2245
r54 6 19 3.12934 $w=6.1e-08 $l=5.18073e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.216 $Y=0.206 $X2=0.199 $Y2=0.162
r55 6 9 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.216 $Y=0.206 $X2=0.216 $Y2=0.2245
r56 4 42 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r57 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends


* END of "./OAI311xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI311xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 C1 Y
* 
* Y	Y
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 noxref_8 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_A2_M1_g noxref_8 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_8 N_A1_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_10 N_B1_M3_g noxref_8 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_C1_M4_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_11 N_A3_M5_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M6 noxref_12 N_A2_M6_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 N_Y_M7_d N_A1_M7_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M8 VDD N_B1_M8_g N_Y_M8_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M9 N_Y_M9_d N_C1_M9_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.189
*
* 
* .include "OAI311xp33_ASAP7_75t_L.pex.sp.OAI311XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI311xp33_ASAP7_75t_L.pex.sp.OAI311XP33_ASAP7_75T_L.pxi"
* File: OAI311xp33_ASAP7_75t_L.pex.sp.OAI311XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:55:33 2017
* 
x_PM_OAI311XP33_ASAP7_75T_L%A3 N_A3_M0_g N_A3_c_2_p N_A3_M5_g A3 VSS
+ PM_OAI311XP33_ASAP7_75T_L%A3
x_PM_OAI311XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_7_n N_A2_M6_g A2 VSS
+ PM_OAI311XP33_ASAP7_75T_L%A2
x_PM_OAI311XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_20_n N_A1_M7_g A1 VSS
+ PM_OAI311XP33_ASAP7_75T_L%A1
x_PM_OAI311XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_33_n N_B1_M8_g B1 VSS
+ PM_OAI311XP33_ASAP7_75T_L%B1
x_PM_OAI311XP33_ASAP7_75T_L%C1 N_C1_M4_g N_C1_c_44_n N_C1_M9_g C1 VSS
+ PM_OAI311XP33_ASAP7_75T_L%C1
x_PM_OAI311XP33_ASAP7_75T_L%Y N_Y_M4_d N_Y_M8_s N_Y_M7_d N_Y_M9_d N_Y_c_57_n
+ N_Y_c_51_n Y N_Y_c_52_n N_Y_c_56_n N_Y_c_58_n N_Y_c_60_n N_Y_c_61_n N_Y_c_64_n
+ VSS PM_OAI311XP33_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_A2_M1_g 0.00347357f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A3_c_2_p N_A2_c_7_n 0.00120426f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A3 A2 0.0026877f $X=0.08 $Y=0.136 $X2=0.134 $Y2=0.136
cc_4 N_A3_M0_g N_A1_M2_g 2.69148e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 VSS A3 2.10206e-19 $X=0.08 $Y=0.136 $X2=0 $Y2=0
cc_6 N_A2_M1_g N_A1_M2_g 0.00325575f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_7 N_A2_c_7_n N_A1_c_20_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_8 A2 A1 0.00565033f $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_9 N_A2_M1_g N_B1_M3_g 2.69148e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_10 VSS A2 0.00132451f $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_11 VSS N_A2_M1_g 2.64276e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_12 VSS A2 0.00125674f $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_13 A2 N_Y_c_51_n 7.83333e-19 $X=0.134 $Y=0.136 $X2=0.081 $Y2=0.135
cc_14 A2 N_Y_c_52_n 4.82846e-19 $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_15 N_A1_M2_g N_B1_M3_g 0.00359705f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_A1_c_20_n N_B1_c_33_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_17 A1 B1 0.00506253f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_18 N_A1_M2_g N_C1_M4_g 2.69148e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_19 VSS A1 0.00114532f $X=0.196 $Y=0.136 $X2=0.081 $Y2=0.135
cc_20 VSS N_A1_M2_g 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_21 VSS A1 0.00125352f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_22 A1 N_Y_c_51_n 0.0013295f $X=0.196 $Y=0.136 $X2=0.081 $Y2=0.135
cc_23 N_A1_M2_g N_Y_c_52_n 2.80442e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 N_B1_M3_g N_C1_M4_g 0.00330657f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_25 N_B1_c_33_n N_C1_c_44_n 9.33263e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_26 B1 C1 0.00624003f $X=0.247 $Y=0.134 $X2=0.135 $Y2=0.135
cc_27 VSS N_B1_M3_g 3.06796e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_28 VSS B1 0.0013399f $X=0.247 $Y=0.134 $X2=0 $Y2=0
cc_29 B1 N_Y_c_51_n 0.00127618f $X=0.247 $Y=0.134 $X2=0 $Y2=0
cc_30 B1 N_Y_c_56_n 0.00123604f $X=0.247 $Y=0.134 $X2=0 $Y2=0
cc_31 C1 N_Y_c_57_n 3.31541e-19 $X=0.297 $Y=0.134 $X2=0.196 $Y2=0.136
cc_32 N_C1_M4_g N_Y_c_58_n 2.56935e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_33 C1 N_Y_c_58_n 0.00123604f $X=0.297 $Y=0.134 $X2=0 $Y2=0
cc_34 C1 N_Y_c_60_n 0.00546796f $X=0.297 $Y=0.134 $X2=0 $Y2=0
cc_35 C1 N_Y_c_61_n 0.0013399f $X=0.297 $Y=0.134 $X2=0 $Y2=0
cc_36 VSS N_Y_c_51_n 0.00107252f $X=0.216 $Y=0.036 $X2=0.081 $Y2=0.135
cc_37 VSS N_Y_c_61_n 0.00147748f $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_38 VSS N_Y_c_64_n 4.51619e-19 $X=0.216 $Y=0.036 $X2=0 $Y2=0

* END of "./OAI311xp33_ASAP7_75t_L.pex.sp.OAI311XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI31xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:55:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI31xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI31xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI31xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:55:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI31XP33_ASAP7_75T_L%A3 2 5 7 13 VSS
c5 13 VSS 0.00742663f $X=0.0855 $Y=0.1355
c6 5 VSS 0.00298625f $X=0.081 $Y=0.135
c7 2 VSS 0.0631569f $X=0.081 $Y=0.054
r8 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.136 $X2=0.081
+ $Y2=0.136
r9 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r10 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI31XP33_ASAP7_75T_L%A2 2 5 7 10 VSS
c12 10 VSS 0.00230441f $X=0.1355 $Y=0.1355
c13 5 VSS 0.00178389f $X=0.135 $Y=0.135
c14 2 VSS 0.059793f $X=0.135 $Y=0.054
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.136 $X2=0.135
+ $Y2=0.136
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI31XP33_ASAP7_75T_L%A1 2 5 7 10 VSS
c13 10 VSS 0.00151062f $X=0.1895 $Y=0.1355
c14 5 VSS 0.00178389f $X=0.189 $Y=0.135
c15 2 VSS 0.0607616f $X=0.189 $Y=0.054
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.136 $X2=0.189
+ $Y2=0.136
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI31XP33_ASAP7_75T_L%B 2 5 7 10 VSS
c8 10 VSS 0.00118636f $X=0.2405 $Y=0.1355
c9 5 VSS 0.00234817f $X=0.243 $Y=0.135
c10 2 VSS 0.0654963f $X=0.243 $Y=0.054
r11 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.136 $X2=0.243
+ $Y2=0.136
r12 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r13 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI31XP33_ASAP7_75T_L%Y 1 4 7 8 11 20 22 27 28 29 37 VSS
c13 37 VSS 0.00203647f $X=0.288 $Y=0.072
c14 36 VSS 0.00163204f $X=0.297 $Y=0.072
c15 31 VSS 7.84313e-19 $X=0.297 $Y=0.2125
c16 29 VSS 9.30571e-20 $X=0.297 $Y=0.1085
c17 28 VSS 0.00131632f $X=0.297 $Y=0.106
c18 27 VSS 0.00408956f $X=0.299 $Y=0.111
c19 25 VSS 6.45213e-19 $X=0.297 $Y=0.225
c20 23 VSS 3.86697e-19 $X=0.256 $Y=0.234
c21 22 VSS 0.00142432f $X=0.252 $Y=0.234
c22 21 VSS 4.1452e-19 $X=0.234 $Y=0.234
c23 20 VSS 0.0039184f $X=0.23 $Y=0.234
c24 15 VSS 0.0088253f $X=0.288 $Y=0.234
c25 11 VSS 0.00531813f $X=0.205 $Y=0.163
c26 4 VSS 0.00174116f $X=0.268 $Y=0.054
r27 37 38 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.2925 $Y2=0.072
r28 36 38 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.072 $X2=0.2925 $Y2=0.072
r29 33 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.072 $X2=0.288 $Y2=0.072
r30 30 31 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.2 $X2=0.297 $Y2=0.2125
r31 28 29 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.1085
r32 27 30 6.04321 $w=1.8e-08 $l=8.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.111 $X2=0.297 $Y2=0.2
r33 27 29 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.111 $X2=0.297 $Y2=0.1085
r34 25 31 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.2125
r35 24 36 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.081 $X2=0.297 $Y2=0.072
r36 24 28 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.081 $X2=0.297 $Y2=0.106
r37 22 23 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.256 $Y2=0.234
r38 21 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r39 20 21 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.234 $X2=0.234 $Y2=0.234
r40 17 20 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.23 $Y2=0.234
r41 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r42 15 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.234 $X2=0.297 $Y2=0.225
r43 15 23 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.256 $Y2=0.234
r44 11 18 61.2798 $w=2.4e-08 $l=7.1e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.163 $X2=0.216 $Y2=0.234
r45 8 11 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2245 $X2=0.216 $Y2=0.2245
r46 7 11 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2245 $X2=0.216 $Y2=0.2245
r47 4 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.072 $X2=0.27
+ $Y2=0.072
r48 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.054 $X2=0.268 $Y2=0.054
.ends


* END of "./OAI31xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI31xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 B Y
* 
* Y	Y
* B	B
* A1	A1
* A2	A2
* A3	A3
M0 noxref_7 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 VSS N_A2_M1_g noxref_7 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 noxref_7 N_A1_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.027
M3 N_Y_M3_d N_B_M3_g noxref_7 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 noxref_9 N_A3_M4_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 noxref_10 N_A2_M5_g noxref_9 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 N_Y_M6_d N_A1_M6_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M7 VDD N_B_M7_g N_Y_M7_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.189
*
* 
* .include "OAI31xp33_ASAP7_75t_L.pex.sp.OAI31XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI31xp33_ASAP7_75t_L.pex.sp.OAI31XP33_ASAP7_75T_L.pxi"
* File: OAI31xp33_ASAP7_75t_L.pex.sp.OAI31XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:55:55 2017
* 
x_PM_OAI31XP33_ASAP7_75T_L%A3 N_A3_M0_g N_A3_c_2_p N_A3_M4_g A3 VSS
+ PM_OAI31XP33_ASAP7_75T_L%A3
x_PM_OAI31XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_7_n N_A2_M5_g A2 VSS
+ PM_OAI31XP33_ASAP7_75T_L%A2
x_PM_OAI31XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_20_n N_A1_M6_g A1 VSS
+ PM_OAI31XP33_ASAP7_75T_L%A1
x_PM_OAI31XP33_ASAP7_75T_L%B N_B_M3_g N_B_c_33_n N_B_M7_g B VSS
+ PM_OAI31XP33_ASAP7_75T_L%B
x_PM_OAI31XP33_ASAP7_75T_L%Y N_Y_M3_d N_Y_c_48_n N_Y_M7_s N_Y_M6_d N_Y_c_39_n
+ N_Y_c_40_n N_Y_c_45_n Y N_Y_c_42_n N_Y_c_47_n N_Y_c_43_n VSS
+ PM_OAI31XP33_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_A2_M1_g 0.00347357f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A3_c_2_p N_A2_c_7_n 9.56181e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A3 A2 0.00802362f $X=0.0855 $Y=0.1355 $X2=0.1355 $Y2=0.1355
cc_4 N_A3_M0_g N_A1_M2_g 2.69148e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 VSS A3 3.31541e-19 $X=0.0855 $Y=0.1355 $X2=0.135 $Y2=0.135
cc_6 N_A2_M1_g N_A1_M2_g 0.00325575f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_7 N_A2_c_7_n N_A1_c_20_n 9.07968e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_8 A2 A1 0.00613955f $X=0.1355 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_9 N_A2_M1_g N_B_M3_g 2.69148e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_10 VSS A2 3.31541e-19 $X=0.1355 $Y=0.1355 $X2=0.081 $Y2=0.135
cc_11 VSS N_A2_M1_g 2.64276e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_12 VSS A2 0.00125674f $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_13 A2 N_Y_c_39_n 7.56932e-19 $X=0.1355 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_14 A2 N_Y_c_40_n 4.56622e-19 $X=0.1355 $Y=0.1355 $X2=0 $Y2=0
cc_15 N_A1_M2_g N_B_M3_g 0.00359705f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_16 N_A1_c_20_n N_B_c_33_n 9.56181e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_17 A1 B 0.00393834f $X=0.1895 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_18 VSS A1 3.61412e-19 $X=0.1895 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_19 VSS N_A1_M2_g 2.64276e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_20 VSS A1 0.00125352f $X=0.1895 $Y=0.1355 $X2=0 $Y2=0
cc_21 A1 N_Y_c_39_n 0.0013295f $X=0.1895 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_22 A1 N_Y_c_42_n 5.26804e-19 $X=0.1895 $Y=0.1355 $X2=0 $Y2=0
cc_23 A1 N_Y_c_43_n 2.59217e-19 $X=0.1895 $Y=0.1355 $X2=0 $Y2=0
cc_24 B N_Y_c_39_n 0.00127618f $X=0.2405 $Y=0.1355 $X2=0 $Y2=0
cc_25 N_B_M3_g N_Y_c_45_n 2.56935e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_26 B N_Y_c_45_n 0.00123064f $X=0.2405 $Y=0.1355 $X2=0 $Y2=0
cc_27 B N_Y_c_47_n 0.00441984f $X=0.2405 $Y=0.1355 $X2=0 $Y2=0
cc_28 VSS N_Y_c_48_n 0.002591f $X=0.216 $Y=0.054 $X2=0.081 $Y2=0.135
cc_29 VSS N_Y_c_48_n 3.09692e-19 $X=0.216 $Y=0.036 $X2=0.081 $Y2=0.135
cc_30 VSS N_Y_c_39_n 9.28287e-19 $X=0.216 $Y=0.054 $X2=0.081 $Y2=0.136
cc_31 VSS N_Y_c_43_n 3.59474e-19 $X=0.216 $Y=0.054 $X2=0 $Y2=0

* END of "./OAI31xp33_ASAP7_75t_L.pex.sp.OAI31XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI31xp67_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:56:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI31xp67_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI31xp67_ASAP7_75t_L.pex.sp.pex"
* File: OAI31xp67_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:56:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI31XP67_ASAP7_75T_L%A3 2 7 10 13 15 28 30 33 VSS
c18 33 VSS 9.55459e-19 $X=0.0605 $Y=0.135
c19 32 VSS 0.00132257f $X=0.04 $Y=0.135
c20 30 VSS 8.29931e-19 $X=0.081 $Y=0.135
c21 28 VSS 0.0115557f $X=0.039 $Y=0.134
c22 13 VSS 0.00776257f $X=0.135 $Y=0.135
c23 10 VSS 0.0623753f $X=0.135 $Y=0.0675
c24 2 VSS 0.0670913f $X=0.081 $Y=0.0675
r25 32 33 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.135 $X2=0.0605 $Y2=0.135
r26 30 33 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0605 $Y2=0.135
r27 28 32 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.039
+ $Y=0.135 $X2=0.04 $Y2=0.135
r28 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r29 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r30 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r31 5 30 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r32 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r33 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI31XP67_ASAP7_75T_L%B 2 7 10 13 24 26 VSS
c35 26 VSS 0.00100406f $X=0.189 $Y=0.135
c36 24 VSS 0.00350472f $X=0.162 $Y=0.131
c37 13 VSS 0.00389607f $X=0.243 $Y=0.135
c38 10 VSS 0.0684522f $X=0.243 $Y=0.0675
c39 2 VSS 0.0623453f $X=0.189 $Y=0.0675
r40 24 26 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.135 $X2=0.189 $Y2=0.135
r41 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r42 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r43 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r44 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r45 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI31XP67_ASAP7_75T_L%A2 2 7 10 13 15 22 26 27 VSS
c28 27 VSS 3.35447e-19 $X=0.3845 $Y=0.135
c29 26 VSS 0.00205662f $X=0.364 $Y=0.135
c30 24 VSS 3.90789e-19 $X=0.405 $Y=0.135
c31 22 VSS 0.00200239f $X=0.331 $Y=0.137
c32 13 VSS 0.00421199f $X=0.459 $Y=0.135
c33 10 VSS 0.0631881f $X=0.459 $Y=0.0675
c34 2 VSS 0.0665455f $X=0.405 $Y=0.0675
r35 26 27 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.364
+ $Y=0.135 $X2=0.3845 $Y2=0.135
r36 24 27 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.3845 $Y2=0.135
r37 22 26 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.331
+ $Y=0.135 $X2=0.364 $Y2=0.135
r38 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r39 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r40 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r41 5 24 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r42 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r43 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OAI31XP67_ASAP7_75T_L%A1 2 7 10 13 15 23 24 25 VSS
c25 25 VSS 7.52043e-19 $X=0.6225 $Y=0.135
c26 24 VSS 7.53212e-19 $X=0.608 $Y=0.135
c27 23 VSS 0.00533219f $X=0.637 $Y=0.134
c28 13 VSS 0.00454174f $X=0.567 $Y=0.135
c29 10 VSS 0.0666959f $X=0.567 $Y=0.0675
c30 2 VSS 0.0631881f $X=0.513 $Y=0.0675
r31 24 25 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.608
+ $Y=0.135 $X2=0.6225 $Y2=0.135
r32 23 25 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.637
+ $Y=0.135 $X2=0.6225 $Y2=0.135
r33 19 24 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.608 $Y2=0.135
r34 13 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r35 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r36 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r37 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r38 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r39 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OAI31XP67_ASAP7_75T_L%Y 1 2 5 6 9 11 12 15 17 18 19 20 22 23 24 25 26
+ 28 29 36 38 39 42 51 56 VSS
c63 57 VSS 2.67452e-19 $X=0.234 $Y=0.198
c64 56 VSS 4.09224e-19 $X=0.243 $Y=0.198
c65 51 VSS 5.91473e-19 $X=0.216 $Y=0.198
c66 48 VSS 1.77025e-19 $X=0.234 $Y=0.072
c67 42 VSS 5.8316e-20 $X=0.216 $Y=0.072
c68 39 VSS 0.00213769f $X=0.6285 $Y=0.234
c69 38 VSS 0.00692832f $X=0.608 $Y=0.234
c70 36 VSS 0.00387584f $X=0.649 $Y=0.234
c71 29 VSS 0.0543395f $X=0.649 $Y=0.072
c72 28 VSS 0.00761484f $X=0.649 $Y=0.072
c73 26 VSS 4.40637e-21 $X=0.554 $Y=0.072
c74 25 VSS 0.00305119f $X=0.553 $Y=0.072
c75 24 VSS 0.00457695f $X=0.419 $Y=0.072
c76 23 VSS 4.75287e-19 $X=0.288 $Y=0.072
c77 20 VSS 1.43629e-19 $X=0.252 $Y=0.072
c78 18 VSS 4.28707e-19 $X=0.243 $Y=0.126
c79 17 VSS 3.66662e-19 $X=0.243 $Y=0.189
c80 15 VSS 0.00283143f $X=0.54 $Y=0.2025
c81 11 VSS 6.03275e-19 $X=0.557 $Y=0.2025
c82 9 VSS 0.00583269f $X=0.214 $Y=0.216
c83 5 VSS 0.00296627f $X=0.216 $Y=0.0675
c84 1 VSS 5.61665e-19 $X=0.233 $Y=0.0675
r85 57 58 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.2385 $Y2=0.198
r86 56 58 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.198 $X2=0.2385 $Y2=0.198
r87 51 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.234 $Y2=0.198
r88 48 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.2385 $Y2=0.072
r89 47 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.072 $X2=0.2385 $Y2=0.072
r90 42 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.072 $X2=0.234 $Y2=0.072
r91 38 39 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.608
+ $Y=0.234 $X2=0.6285 $Y2=0.234
r92 36 39 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.649
+ $Y=0.234 $X2=0.6285 $Y2=0.234
r93 36 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.649 $Y=0.234 $X2=0.649
+ $Y2=0.234
r94 32 38 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.608 $Y2=0.234
r95 29 37 139.821 $w=2.4e-08 $l=1.62e-07 $layer=LISD $thickness=2.8e-08 $X=0.649
+ $Y=0.072 $X2=0.649 $Y2=0.234
r96 28 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.649 $Y=0.072 $X2=0.649
+ $Y2=0.072
r97 25 26 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.553
+ $Y=0.072 $X2=0.554 $Y2=0.072
r98 24 25 9.09877 $w=1.8e-08 $l=1.34e-07 $layer=M1 $thickness=3.6e-08 $X=0.419
+ $Y=0.072 $X2=0.553 $Y2=0.072
r99 23 24 8.89506 $w=1.8e-08 $l=1.31e-07 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.419 $Y2=0.072
r100 22 28 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.619
+ $Y=0.072 $X2=0.649 $Y2=0.072
r101 22 26 4.41358 $w=1.8e-08 $l=6.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.619
+ $Y=0.072 $X2=0.554 $Y2=0.072
r102 20 47 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.072 $X2=0.243 $Y2=0.072
r103 20 23 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.072 $X2=0.288 $Y2=0.072
r104 18 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.144
r105 17 56 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.198
r106 17 19 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.144
r107 16 47 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.072
r108 16 18 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.126
r109 15 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r110 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r111 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r112 9 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r113 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.216 $X2=0.214 $Y2=0.216
r114 5 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072 $X2=0.216
+ $Y2=0.072
r115 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r116 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./OAI31xp67_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI31xp67_ASAP7_75t_L  VSS VDD A3 B A2 A1 Y
* 
* Y	Y
* A1	A1
* A2	A2
* B	B
* A3	A3
M0 VSS N_A3_M0_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_A3_M1_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_B_M2_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_Y_M3_d N_B_M3_g noxref_7 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_7 N_A2_M4_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 noxref_7 N_A2_M5_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 noxref_7 N_A1_M6_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M7 noxref_7 N_A1_M7_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M8 noxref_8 N_A3_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M9 noxref_8 N_A3_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M10 N_Y_M10_d N_B_M10_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M11 noxref_8 N_A2_M11_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M12 noxref_8 N_A2_M12_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M13 N_Y_M13_d N_A1_M13_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
M14 N_Y_M14_d N_A1_M14_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
*
* 
* .include "OAI31xp67_ASAP7_75t_L.pex.sp.OAI31XP67_ASAP7_75T_L.pxi"
* BEGIN of "./OAI31xp67_ASAP7_75t_L.pex.sp.OAI31XP67_ASAP7_75T_L.pxi"
* File: OAI31xp67_ASAP7_75t_L.pex.sp.OAI31XP67_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:56:18 2017
* 
x_PM_OAI31XP67_ASAP7_75T_L%A3 N_A3_M0_g N_A3_M8_g N_A3_M1_g N_A3_c_4_p N_A3_M9_g
+ A3 N_A3_c_8_p N_A3_c_13_p VSS PM_OAI31XP67_ASAP7_75T_L%A3
x_PM_OAI31XP67_ASAP7_75T_L%B N_B_M2_g N_B_M10_g N_B_M3_g N_B_c_22_n B N_B_c_27_n
+ VSS PM_OAI31XP67_ASAP7_75T_L%B
x_PM_OAI31XP67_ASAP7_75T_L%A2 N_A2_M4_g N_A2_M11_g N_A2_M5_g N_A2_c_57_p
+ N_A2_M12_g A2 N_A2_c_62_p N_A2_c_68_p VSS PM_OAI31XP67_ASAP7_75T_L%A2
x_PM_OAI31XP67_ASAP7_75T_L%A1 N_A1_M6_g N_A1_M13_g N_A1_M7_g N_A1_c_85_n
+ N_A1_M14_g A1 N_A1_c_93_p N_A1_c_95_p VSS PM_OAI31XP67_ASAP7_75T_L%A1
x_PM_OAI31XP67_ASAP7_75T_L%Y N_Y_M3_d N_Y_M2_d N_Y_c_108_n N_Y_M10_d N_Y_c_109_n
+ N_Y_M14_d N_Y_M13_d N_Y_c_130_n N_Y_c_110_n N_Y_c_113_n N_Y_c_116_n
+ N_Y_c_147_n Y N_Y_c_148_n N_Y_c_124_n N_Y_c_127_n N_Y_c_133_n N_Y_c_134_n
+ N_Y_c_136_n N_Y_c_138_n N_Y_c_139_n N_Y_c_141_n N_Y_c_118_n N_Y_c_120_n
+ N_Y_c_128_n VSS PM_OAI31XP67_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_B_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_A3_M1_g N_B_M2_g 0.00323392f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A3_M1_g N_B_M3_g 2.69148e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_4 N_A3_c_4_p N_B_c_22_n 0.00149358f $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_5 N_A3_M1_g B 0.00143821f $X=0.135 $Y=0.0675 $X2=0.162 $Y2=0.131
cc_6 N_A3_c_4_p B 0.00199657f $X=0.135 $Y=0.135 $X2=0.162 $Y2=0.131
cc_7 A3 B 0.00112126f $X=0.039 $Y=0.134 $X2=0.162 $Y2=0.131
cc_8 N_A3_c_8_p B 9.16541e-19 $X=0.081 $Y=0.135 $X2=0.162 $Y2=0.131
cc_9 N_A3_c_4_p N_B_c_27_n 4.61613e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_10 VSS A3 0.00142719f $X=0.039 $Y=0.134 $X2=0 $Y2=0
cc_11 VSS N_A3_M0_g 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_12 VSS N_A3_c_4_p 6.39404e-19 $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_13 VSS N_A3_c_13_p 0.00103581f $X=0.0605 $Y=0.135 $X2=0.243 $Y2=0.135
cc_14 VSS N_A3_M1_g 2.56935e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 VSS N_A3_c_4_p 3.80485e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_16 VSS N_A3_c_4_p 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_17 VSS N_A3_c_4_p 3.22497e-19 $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_18 VSS N_A3_M1_g 2.64276e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 VSS B 0.00129462f $X=0.162 $Y=0.131 $X2=0.04 $Y2=0.135
cc_20 VSS B 0.00123604f $X=0.162 $Y=0.131 $X2=0 $Y2=0
cc_21 VSS N_B_c_27_n 5.19988e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_22 VSS N_B_M2_g 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_23 VSS N_B_c_27_n 5.19988e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_24 VSS N_B_M3_g 2.08515e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_25 VSS B 0.00132102f $X=0.162 $Y=0.131 $X2=0.081 $Y2=0.135
cc_26 VSS B 0.00125352f $X=0.162 $Y=0.131 $X2=0 $Y2=0
cc_27 VSS N_B_M2_g 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_28 VSS N_B_c_27_n 0.00103934f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_29 VSS N_B_M3_g 2.38303e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_B_c_22_n N_Y_M3_d 3.8028e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_31 N_B_c_22_n N_Y_c_108_n 9.18375e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_32 N_B_c_22_n N_Y_c_109_n 3.82299e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_33 N_B_M3_g N_Y_c_110_n 2.67951e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_34 N_B_c_22_n N_Y_c_110_n 4.86057e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_35 B N_Y_c_110_n 6.4382e-19 $X=0.162 $Y=0.131 $X2=0 $Y2=0
cc_36 N_B_M3_g N_Y_c_113_n 2.57919e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_B_c_22_n N_Y_c_113_n 4.68063e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_38 B N_Y_c_113_n 5.38082e-19 $X=0.162 $Y=0.131 $X2=0 $Y2=0
cc_39 N_B_c_22_n N_Y_c_116_n 0.00127415f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_40 N_B_c_27_n N_Y_c_116_n 8.41056e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_41 N_B_c_22_n N_Y_c_118_n 4.39606e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_42 B N_Y_c_118_n 2.11326e-19 $X=0.162 $Y=0.131 $X2=0 $Y2=0
cc_43 N_B_c_22_n N_Y_c_120_n 4.02804e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_44 B N_Y_c_120_n 2.08234e-19 $X=0.162 $Y=0.131 $X2=0 $Y2=0
cc_45 N_A2_M4_g N_A1_M6_g 2.74891e-19 $X=0.405 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_46 N_A2_M5_g N_A1_M6_g 0.00335739f $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_47 N_A2_M5_g N_A1_M7_g 2.74891e-19 $X=0.459 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_48 N_A2_c_57_p N_A1_c_85_n 0.00170501f $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.135
cc_49 VSS N_A2_c_57_p 3.80413e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_50 VSS N_A2_c_57_p 8.00061e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_51 VSS N_A2_M4_g 2.64781e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_52 VSS N_A2_M5_g 2.64781e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_53 VSS N_A2_c_62_p 3.34398e-19 $X=0.364 $Y=0.135 $X2=0 $Y2=0
cc_54 VSS N_A2_c_57_p 3.80413e-19 $X=0.459 $Y=0.135 $X2=0.189 $Y2=0.216
cc_55 VSS N_A2_c_57_p 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_56 VSS N_A2_M4_g 2.21754e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_57 VSS A2 0.00124544f $X=0.331 $Y=0.137 $X2=0.189 $Y2=0.135
cc_58 VSS N_A2_c_62_p 7.18834e-19 $X=0.364 $Y=0.135 $X2=0.189 $Y2=0.135
cc_59 VSS N_A2_c_68_p 7.18834e-19 $X=0.3845 $Y=0.135 $X2=0.189 $Y2=0.135
cc_60 A2 N_Y_c_110_n 0.001255f $X=0.331 $Y=0.137 $X2=0 $Y2=0
cc_61 A2 N_Y_c_116_n 0.001255f $X=0.331 $Y=0.137 $X2=0 $Y2=0
cc_62 N_A2_M4_g N_Y_c_124_n 3.31725e-19 $X=0.405 $Y=0.0675 $X2=0.162 $Y2=0.131
cc_63 N_A2_c_57_p N_Y_c_124_n 7.97733e-19 $X=0.459 $Y=0.135 $X2=0.162 $Y2=0.131
cc_64 A2 N_Y_c_124_n 0.00511299f $X=0.331 $Y=0.137 $X2=0.162 $Y2=0.131
cc_65 N_A2_M5_g N_Y_c_127_n 3.99641e-19 $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_66 A2 N_Y_c_128_n 0.001255f $X=0.331 $Y=0.137 $X2=0 $Y2=0
cc_67 VSS A2 6.31608e-19 $X=0.331 $Y=0.137 $X2=0.189 $Y2=0.135
cc_68 VSS N_A2_M4_g 3.31725e-19 $X=0.405 $Y=0.0675 $X2=0.162 $Y2=0.135
cc_69 VSS N_A2_c_57_p 7.90552e-19 $X=0.459 $Y=0.135 $X2=0.162 $Y2=0.135
cc_70 VSS A2 3.52753e-19 $X=0.331 $Y=0.137 $X2=0.162 $Y2=0.135
cc_71 VSS N_A2_c_68_p 0.00189591f $X=0.3845 $Y=0.135 $X2=0.162 $Y2=0.135
cc_72 VSS N_A2_M5_g 4.95023e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_73 VSS N_A1_c_85_n 3.80413e-19 $X=0.567 $Y=0.135 $X2=0.331 $Y2=0.135
cc_74 VSS N_A1_M6_g 2.64781e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_75 VSS N_A1_c_85_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_76 N_A1_c_85_n N_Y_M14_d 3.80413e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_77 N_A1_c_85_n N_Y_c_130_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0.459 $Y2=0.2025
cc_78 N_A1_M6_g N_Y_c_127_n 3.99641e-19 $X=0.513 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_79 N_A1_c_85_n N_Y_c_127_n 8.21544e-19 $X=0.567 $Y=0.135 $X2=0.405 $Y2=0.135
cc_80 N_A1_c_93_p N_Y_c_133_n 0.00192512f $X=0.608 $Y=0.135 $X2=0.364 $Y2=0.135
cc_81 N_A1_M7_g N_Y_c_134_n 4.27107e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_82 N_A1_c_95_p N_Y_c_134_n 0.00192512f $X=0.6225 $Y=0.135 $X2=0 $Y2=0
cc_83 N_A1_c_85_n N_Y_c_136_n 8.89529e-19 $X=0.567 $Y=0.135 $X2=0.405 $Y2=0.135
cc_84 A1 N_Y_c_136_n 0.00624991f $X=0.637 $Y=0.134 $X2=0.405 $Y2=0.135
cc_85 A1 N_Y_c_138_n 3.98708e-19 $X=0.637 $Y=0.134 $X2=0 $Y2=0
cc_86 N_A1_M7_g N_Y_c_139_n 2.64781e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_87 N_A1_c_93_p N_Y_c_139_n 3.98708e-19 $X=0.608 $Y=0.135 $X2=0 $Y2=0
cc_88 N_A1_c_95_p N_Y_c_141_n 3.98708e-19 $X=0.6225 $Y=0.135 $X2=0 $Y2=0
cc_89 VSS N_A1_M7_g 3.31725e-19 $X=0.567 $Y=0.0675 $X2=0.364 $Y2=0.135
cc_90 VSS A1 2.46082e-19 $X=0.637 $Y=0.134 $X2=0.364 $Y2=0.135
cc_91 VSS N_A1_c_93_p 0.00188722f $X=0.608 $Y=0.135 $X2=0.364 $Y2=0.135
cc_92 VSS N_A1_M6_g 4.95023e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_93 VSS N_A1_c_85_n 8.17112e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_94 VSS N_Y_c_108_n 0.0038699f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_95 VSS N_Y_c_108_n 0.0034183f $X=0.27 $Y=0.036 $X2=0.081 $Y2=0.135
cc_96 VSS N_Y_c_108_n 0.00249183f $X=0.236 $Y=0.036 $X2=0.081 $Y2=0.135
cc_97 VSS N_Y_c_130_n 0.00169333f $X=0.54 $Y=0.036 $X2=0.135 $Y2=0.2025
cc_98 VSS N_Y_c_113_n 4.92442e-19 $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_99 VSS N_Y_c_147_n 0.0145014f $X=0.54 $Y=0.036 $X2=0 $Y2=0
cc_100 VSS N_Y_c_148_n 3.27573e-19 $X=0.268 $Y=0.0675 $X2=0 $Y2=0
cc_101 VSS N_Y_c_148_n 0.00262229f $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_102 VSS N_Y_c_127_n 0.00226064f $X=0.432 $Y=0.036 $X2=0 $Y2=0
cc_103 VSS N_Y_c_127_n 0.00226064f $X=0.54 $Y=0.036 $X2=0 $Y2=0
cc_104 VSS N_Y_c_118_n 4.4805e-19 $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_105 VSS N_Y_c_118_n 0.0145014f $X=0.236 $Y=0.036 $X2=0 $Y2=0
cc_106 VSS N_Y_c_109_n 0.00319086f $X=0.252 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_107 VSS N_Y_c_148_n 2.71189e-19 $X=0.288 $Y=0.234 $X2=0 $Y2=0
cc_108 VSS N_Y_c_124_n 2.71189e-19 $X=0.364 $Y=0.234 $X2=0 $Y2=0
cc_109 VSS N_Y_c_139_n 3.08222e-19 $X=0.432 $Y=0.234 $X2=0 $Y2=0
cc_110 VSS N_Y_c_120_n 0.00464705f $X=0.252 $Y=0.234 $X2=0 $Y2=0
cc_111 VSS N_Y_c_130_n 0.00318647f $X=0.54 $Y=0.2025 $X2=0.135 $Y2=0.0675
cc_112 VSS N_Y_c_139_n 4.47473e-19 $X=0.608 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_113 VSS N_Y_c_130_n 0.00350507f $X=0.54 $Y=0.2025 $X2=0.135 $Y2=0.2025
cc_114 VSS N_Y_c_136_n 0.00464962f $X=0.649 $Y=0.072 $X2=0.135 $Y2=0.2025
cc_115 VSS N_Y_c_139_n 0.00251885f $X=0.608 $Y=0.234 $X2=0.135 $Y2=0.2025
cc_116 VSS N_Y_c_124_n 3.52391e-19 $X=0.419 $Y=0.072 $X2=0 $Y2=0
cc_117 VSS N_Y_c_127_n 3.52391e-19 $X=0.553 $Y=0.072 $X2=0 $Y2=0
cc_118 VSS N_Y_c_136_n 2.23682e-19 $X=0.649 $Y=0.072 $X2=0 $Y2=0
cc_119 VSS N_Y_c_130_n 0.00226064f $X=0.54 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_120 VSS N_Y_c_134_n 3.52391e-19 $X=0.649 $Y=0.072 $X2=0.081 $Y2=0.135
cc_121 VSS N_Y_c_139_n 0.00705122f $X=0.608 $Y=0.234 $X2=0.081 $Y2=0.135

* END of "./OAI31xp67_ASAP7_75t_L.pex.sp.OAI31XP67_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI321xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:56:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI321xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI321xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI321xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:56:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI321XP33_ASAP7_75T_L%A3 2 5 7 19 VSS
c5 19 VSS 0.0184885f $X=0.08 $Y=0.136
c6 5 VSS 0.00275452f $X=0.081 $Y=0.135
c7 2 VSS 0.0643308f $X=0.081 $Y=0.0675
r8 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r9 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r10 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI321XP33_ASAP7_75T_L%A2 2 5 7 15 VSS
c11 15 VSS 0.00290906f $X=0.134 $Y=0.136
c12 5 VSS 0.00132829f $X=0.135 $Y=0.135
c13 2 VSS 0.0599284f $X=0.135 $Y=0.0675
r14 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI321XP33_ASAP7_75T_L%A1 2 5 7 13 VSS
c12 13 VSS 0.00103414f $X=0.196 $Y=0.136
c13 5 VSS 0.00119626f $X=0.189 $Y=0.135
c14 2 VSS 0.0606313f $X=0.189 $Y=0.0675
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI321XP33_ASAP7_75T_L%C 2 5 7 10 VSS
c11 10 VSS 0.00128201f $X=0.243 $Y=0.134
c12 5 VSS 0.00120688f $X=0.243 $Y=0.135
c13 2 VSS 0.061622f $X=0.243 $Y=0.0675
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI321XP33_ASAP7_75T_L%B1 2 5 7 10 VSS
c11 10 VSS 9.49292e-19 $X=0.296 $Y=0.134
c12 5 VSS 0.00113128f $X=0.297 $Y=0.135
c13 2 VSS 0.0619691f $X=0.297 $Y=0.0675
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OAI321XP33_ASAP7_75T_L%B2 2 5 7 10 VSS
c11 10 VSS 5.93188e-19 $X=0.348 $Y=0.134
c12 5 VSS 0.00170643f $X=0.351 $Y=0.135
c13 2 VSS 0.066866f $X=0.351 $Y=0.0675
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.216
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OAI321XP33_ASAP7_75T_L%Y 1 2 5 7 8 10 13 19 26 27 32 35 38 40 45 46
+ 49 50 VSS
c28 50 VSS 0.00423691f $X=0.405 $Y=0.2
c29 49 VSS 0.00112176f $X=0.405 $Y=0.106
c30 48 VSS 0.00112176f $X=0.405 $Y=0.225
c31 46 VSS 8.46035e-21 $X=0.36 $Y=0.072
c32 45 VSS 4.59335e-19 $X=0.342 $Y=0.072
c33 40 VSS 0.00240073f $X=0.396 $Y=0.072
c34 39 VSS 8.90106e-19 $X=0.369 $Y=0.234
c35 38 VSS 0.00142296f $X=0.36 $Y=0.234
c36 37 VSS 0.00310342f $X=0.342 $Y=0.234
c37 36 VSS 4.3113e-19 $X=0.31 $Y=0.234
c38 35 VSS 0.00146362f $X=0.306 $Y=0.234
c39 34 VSS 0.00554947f $X=0.288 $Y=0.234
c40 33 VSS 4.31197e-19 $X=0.256 $Y=0.234
c41 32 VSS 0.00142296f $X=0.252 $Y=0.234
c42 28 VSS 4.19362e-19 $X=0.234 $Y=0.234
c43 27 VSS 0.00376122f $X=0.23 $Y=0.234
c44 20 VSS 0.00614869f $X=0.396 $Y=0.234
c45 19 VSS 0.00474306f $X=0.216 $Y=0.2025
c46 13 VSS 0.00345731f $X=0.376 $Y=0.216
c47 9 VSS 5.22702e-19 $X=0.216 $Y=0.2245
c48 5 VSS 0.00233317f $X=0.324 $Y=0.0675
c49 1 VSS 5.75997e-19 $X=0.341 $Y=0.0675
r50 49 50 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.106 $X2=0.405 $Y2=0.2
r51 48 50 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.2
r52 47 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.081 $X2=0.405 $Y2=0.106
r53 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.072 $X2=0.36 $Y2=0.072
r54 42 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.072 $X2=0.342 $Y2=0.072
r55 40 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.072 $X2=0.405 $Y2=0.081
r56 40 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.072 $X2=0.36 $Y2=0.072
r57 38 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.369 $Y2=0.234
r58 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r59 36 37 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.31
+ $Y=0.234 $X2=0.342 $Y2=0.234
r60 35 36 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.31 $Y2=0.234
r61 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r62 33 34 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.234 $X2=0.288 $Y2=0.234
r63 32 33 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.256 $Y2=0.234
r64 30 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.369 $Y2=0.234
r65 27 28 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.234 $X2=0.234 $Y2=0.234
r66 26 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.234 $X2=0.252 $Y2=0.234
r67 26 28 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.234 $X2=0.234 $Y2=0.234
r68 22 27 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.23 $Y2=0.234
r69 20 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r70 20 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.378 $Y2=0.234
r71 19 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r72 13 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r73 10 13 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.216 $X2=0.376 $Y2=0.216
r74 8 9 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.2245 $X2=0.216 $Y2=0.2245
r75 7 9 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2245 $X2=0.216 $Y2=0.2245
r76 6 19 3.12934 $w=6.1e-08 $l=5.18073e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.216 $Y=0.206 $X2=0.199 $Y2=0.162
r77 6 9 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.216 $Y=0.206 $X2=0.216 $Y2=0.2245
r78 5 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.072 $X2=0.324
+ $Y2=0.072
r79 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.324 $Y2=0.0675
r80 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.0675 $X2=0.324 $Y2=0.0675
.ends


* END of "./OAI321xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI321xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 C B1 B2 Y
* 
* Y	Y
* B2	B2
* B1	B1
* C	C
* A1	A1
* A2	A2
* A3	A3
M0 noxref_9 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_A2_M1_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_9 N_A1_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_10 N_C_M3_g noxref_9 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_B1_M4_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_10 N_B2_M5_g N_Y_M5_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_12 N_A3_M6_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 noxref_13 N_A2_M7_g noxref_12 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 N_Y_M8_d N_A1_M8_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 VDD N_C_M9_g N_Y_M9_s VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.189
M10 noxref_14 N_B1_M10_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.189
M11 N_Y_M11_d N_B2_M11_g noxref_14 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.341 $Y=0.189
*
* 
* .include "OAI321xp33_ASAP7_75t_L.pex.sp.OAI321XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI321xp33_ASAP7_75t_L.pex.sp.OAI321XP33_ASAP7_75T_L.pxi"
* File: OAI321xp33_ASAP7_75t_L.pex.sp.OAI321XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:56:41 2017
* 
x_PM_OAI321XP33_ASAP7_75T_L%A3 N_A3_M0_g N_A3_c_2_p N_A3_M6_g A3 VSS
+ PM_OAI321XP33_ASAP7_75T_L%A3
x_PM_OAI321XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_7_n N_A2_M7_g A2 VSS
+ PM_OAI321XP33_ASAP7_75T_L%A2
x_PM_OAI321XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_19_n N_A1_M8_g A1 VSS
+ PM_OAI321XP33_ASAP7_75T_L%A1
x_PM_OAI321XP33_ASAP7_75T_L%C N_C_M3_g N_C_c_31_n N_C_M9_g C VSS
+ PM_OAI321XP33_ASAP7_75T_L%C
x_PM_OAI321XP33_ASAP7_75T_L%B1 N_B1_M4_g N_B1_c_42_n N_B1_M10_g B1 VSS
+ PM_OAI321XP33_ASAP7_75T_L%B1
x_PM_OAI321XP33_ASAP7_75T_L%B2 N_B2_M5_g N_B2_c_53_n N_B2_M11_g B2 VSS
+ PM_OAI321XP33_ASAP7_75T_L%B2
x_PM_OAI321XP33_ASAP7_75T_L%Y N_Y_M5_s N_Y_M4_d N_Y_c_80_n N_Y_M9_s N_Y_M8_d
+ N_Y_M11_d N_Y_c_71_n N_Y_c_62_n Y N_Y_c_63_n N_Y_c_67_n N_Y_c_69_n N_Y_c_72_n
+ N_Y_c_84_n N_Y_c_79_n N_Y_c_74_n N_Y_c_89_n N_Y_c_76_n VSS
+ PM_OAI321XP33_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_A2_M1_g 0.00347357f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A3_c_2_p N_A2_c_7_n 0.00120426f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A3 A2 0.00247926f $X=0.08 $Y=0.136 $X2=0.134 $Y2=0.136
cc_4 N_A3_M0_g N_A1_M2_g 2.69148e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 VSS A3 3.43147e-19 $X=0.08 $Y=0.136 $X2=0 $Y2=0
cc_6 N_A2_M1_g N_A1_M2_g 0.00325575f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_7 N_A2_c_7_n N_A1_c_19_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_8 A2 A1 0.00465395f $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_9 N_A2_M1_g N_C_M3_g 2.69148e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_10 VSS N_A2_M1_g 3.62029e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_11 VSS A2 0.0012376f $X=0.134 $Y=0.136 $X2=0.081 $Y2=0.135
cc_12 A2 N_Y_c_62_n 6.82426e-19 $X=0.134 $Y=0.136 $X2=0.08 $Y2=0.136
cc_13 A2 N_Y_c_63_n 4.83329e-19 $X=0.134 $Y=0.136 $X2=0 $Y2=0
cc_14 N_A1_M2_g N_C_M3_g 0.00359705f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_15 N_A1_c_19_n N_C_c_31_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_16 A1 C 0.00406615f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_17 N_A1_M2_g N_B1_M4_g 2.69148e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_18 VSS N_A1_M2_g 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_19 VSS A1 0.0012322f $X=0.196 $Y=0.136 $X2=0 $Y2=0
cc_20 A1 N_Y_c_62_n 0.0013295f $X=0.196 $Y=0.136 $X2=0.08 $Y2=0.136
cc_21 N_A1_M2_g N_Y_c_63_n 2.84579e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_22 N_C_M3_g N_B1_M4_g 0.00330657f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_23 N_C_c_31_n N_B1_c_42_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_24 C B1 0.00453023f $X=0.243 $Y=0.134 $X2=0.135 $Y2=0.135
cc_25 N_C_M3_g N_B2_M5_g 2.74891e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_26 C N_Y_c_62_n 0.00127618f $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_27 N_C_M3_g N_Y_c_67_n 2.56935e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_28 C N_Y_c_67_n 0.00123064f $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_29 N_B1_M4_g N_B2_M5_g 0.00372052f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_30 N_B1_c_42_n N_B2_c_53_n 9.33263e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_31 B1 B2 0.00484406f $X=0.296 $Y=0.134 $X2=0.189 $Y2=0.135
cc_32 VSS N_B1_M4_g 3.57119e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_33 VSS B1 5.37372e-19 $X=0.296 $Y=0.134 $X2=0 $Y2=0
cc_34 N_B1_M4_g N_Y_c_69_n 2.64276e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_35 B1 N_Y_c_69_n 0.00124805f $X=0.296 $Y=0.134 $X2=0 $Y2=0
cc_36 VSS N_B2_M5_g 2.08515e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_37 B2 N_Y_c_71_n 3.87865e-19 $X=0.348 $Y=0.134 $X2=0.243 $Y2=0.135
cc_38 N_B2_M5_g N_Y_c_72_n 2.56935e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_39 B2 N_Y_c_72_n 0.00123064f $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_40 N_B2_M5_g N_Y_c_74_n 2.76185e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_41 B2 N_Y_c_74_n 0.0012322f $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_42 B2 N_Y_c_76_n 0.00441847f $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_43 VSS N_Y_c_62_n 0.00138157f $X=0.216 $Y=0.0675 $X2=0.08 $Y2=0.136
cc_44 VSS N_Y_c_63_n 2.10682e-19 $X=0.216 $Y=0.072 $X2=0 $Y2=0
cc_45 VSS N_Y_c_79_n 2.88175e-19 $X=0.216 $Y=0.072 $X2=0 $Y2=0
cc_46 VSS N_Y_c_80_n 0.0033367f $X=0.27 $Y=0.036 $X2=0.243 $Y2=0.135
cc_47 VSS N_Y_c_80_n 0.00371671f $X=0.378 $Y=0.036 $X2=0.243 $Y2=0.135
cc_48 VSS N_Y_c_80_n 0.00250965f $X=0.344 $Y=0.036 $X2=0.243 $Y2=0.135
cc_49 VSS N_Y_c_71_n 9.98826e-19 $X=0.378 $Y=0.036 $X2=0.243 $Y2=0.135
cc_50 VSS N_Y_c_84_n 2.47657e-19 $X=0.376 $Y=0.0675 $X2=0 $Y2=0
cc_51 VSS N_Y_c_84_n 0.00260156f $X=0.378 $Y=0.036 $X2=0 $Y2=0
cc_52 VSS N_Y_c_79_n 4.49388e-19 $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_53 VSS N_Y_c_79_n 0.00369159f $X=0.344 $Y=0.036 $X2=0 $Y2=0
cc_54 VSS N_Y_c_74_n 0.00369159f $X=0.378 $Y=0.036 $X2=0 $Y2=0
cc_55 VSS N_Y_c_89_n 3.97918e-19 $X=0.378 $Y=0.036 $X2=0 $Y2=0

* END of "./OAI321xp33_ASAP7_75t_L.pex.sp.OAI321XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI322xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:57:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI322xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI322xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI322xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:57:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI322XP33_ASAP7_75T_L%B2 2 5 7 10 VSS
c8 10 VSS 0.00502923f $X=0.075 $Y=0.134
c9 5 VSS 0.00230059f $X=0.081 $Y=0.135
c10 2 VSS 0.0649001f $X=0.081 $Y=0.0675
r11 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r12 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r13 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI322XP33_ASAP7_75T_L%B1 2 5 7 10 VSS
c10 10 VSS 0.00111927f $X=0.131 $Y=0.134
c11 5 VSS 0.00123757f $X=0.135 $Y=0.135
c12 2 VSS 0.0618833f $X=0.135 $Y=0.0675
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI322XP33_ASAP7_75T_L%A1 2 5 7 10 VSS
c13 10 VSS 4.81053e-19 $X=0.187 $Y=0.136
c14 5 VSS 0.00111823f $X=0.189 $Y=0.135
c15 2 VSS 0.0618966f $X=0.189 $Y=0.0675
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI322XP33_ASAP7_75T_L%A2 2 5 7 13 VSS
c13 13 VSS 4.81053e-19 $X=0.247 $Y=0.136
c14 5 VSS 0.00112315f $X=0.243 $Y=0.135
c15 2 VSS 0.0623167f $X=0.243 $Y=0.0675
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI322XP33_ASAP7_75T_L%A3 2 5 7 15 VSS
c12 15 VSS 7.63284e-19 $X=0.296 $Y=0.136
c13 5 VSS 0.00110907f $X=0.297 $Y=0.135
c14 2 VSS 0.0620676f $X=0.297 $Y=0.0675
r15 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OAI322XP33_ASAP7_75T_L%C2 2 5 7 10 VSS
c11 10 VSS 0.00117666f $X=0.348 $Y=0.134
c12 5 VSS 0.00113128f $X=0.351 $Y=0.135
c13 2 VSS 0.062389f $X=0.351 $Y=0.0675
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.216
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OAI322XP33_ASAP7_75T_L%C1 2 5 7 10 VSS
c11 10 VSS 5.93188e-19 $X=0.405 $Y=0.134
c12 5 VSS 0.00170643f $X=0.405 $Y=0.135
c13 2 VSS 0.066866f $X=0.405 $Y=0.0675
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r15 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.216
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OAI322XP33_ASAP7_75T_L%Y 1 2 5 7 8 10 13 19 26 27 28 29 30 34 35 37
+ 39 42 44 49 50 53 55 VSS
c35 56 VSS 5.10117e-19 $X=0.459 $Y=0.2125
c36 55 VSS 0.00416781f $X=0.459 $Y=0.2
c37 54 VSS 9.06404e-21 $X=0.459 $Y=0.106
c38 53 VSS 0.00108865f $X=0.459 $Y=0.105
c39 52 VSS 6.07272e-19 $X=0.459 $Y=0.225
c40 50 VSS 8.46035e-21 $X=0.414 $Y=0.072
c41 49 VSS 4.59335e-19 $X=0.396 $Y=0.072
c42 44 VSS 0.00240073f $X=0.45 $Y=0.072
c43 43 VSS 8.90106e-19 $X=0.423 $Y=0.234
c44 42 VSS 0.00142296f $X=0.414 $Y=0.234
c45 41 VSS 0.00310342f $X=0.396 $Y=0.234
c46 40 VSS 4.17449e-19 $X=0.364 $Y=0.234
c47 39 VSS 0.00146362f $X=0.36 $Y=0.234
c48 38 VSS 0.00666605f $X=0.342 $Y=0.234
c49 37 VSS 0.00146362f $X=0.306 $Y=0.234
c50 36 VSS 4.17449e-19 $X=0.288 $Y=0.234
c51 35 VSS 0.00307159f $X=0.284 $Y=0.234
c52 34 VSS 8.53778e-19 $X=0.252 $Y=0.234
c53 30 VSS 7.04757e-19 $X=0.241 $Y=0.234
c54 29 VSS 0.00340162f $X=0.234 $Y=0.234
c55 28 VSS 0.00146362f $X=0.198 $Y=0.234
c56 27 VSS 0.0039381f $X=0.18 $Y=0.234
c57 20 VSS 0.00615748f $X=0.45 $Y=0.234
c58 19 VSS 0.00305925f $X=0.162 $Y=0.2025
c59 13 VSS 0.00345731f $X=0.43 $Y=0.216
c60 9 VSS 5.57323e-19 $X=0.162 $Y=0.2245
c61 5 VSS 0.00234286f $X=0.378 $Y=0.0675
c62 1 VSS 5.75997e-19 $X=0.395 $Y=0.0675
r63 55 56 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.2 $X2=0.459 $Y2=0.2125
r64 54 55 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.106 $X2=0.459 $Y2=0.2
r65 53 54 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.105 $X2=0.459 $Y2=0.106
r66 52 56 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.2125
r67 51 53 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.105
r68 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.072 $X2=0.414 $Y2=0.072
r69 46 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.396 $Y2=0.072
r70 44 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.072 $X2=0.459 $Y2=0.081
r71 44 50 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.072 $X2=0.414 $Y2=0.072
r72 42 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.423 $Y2=0.234
r73 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r74 40 41 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.364
+ $Y=0.234 $X2=0.396 $Y2=0.234
r75 39 40 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.364 $Y2=0.234
r76 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r77 37 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.342 $Y2=0.234
r78 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r79 35 36 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.234 $X2=0.288 $Y2=0.234
r80 34 35 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.284 $Y2=0.234
r81 32 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.423 $Y2=0.234
r82 29 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.241 $Y2=0.234
r83 28 29 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.234 $Y2=0.234
r84 27 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r85 26 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.234 $X2=0.252 $Y2=0.234
r86 26 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.234 $X2=0.241 $Y2=0.234
r87 22 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r88 20 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r89 20 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.432 $Y2=0.234
r90 19 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r91 13 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r92 10 13 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.216 $X2=0.43 $Y2=0.216
r93 8 9 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.2245 $X2=0.162 $Y2=0.2245
r94 7 9 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2245 $X2=0.162 $Y2=0.2245
r95 6 19 3.12934 $w=6.1e-08 $l=2.40416e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.162 $Y=0.206 $X2=0.145 $Y2=0.189
r96 6 9 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.162 $Y=0.206 $X2=0.162 $Y2=0.2245
r97 5 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.072 $X2=0.378
+ $Y2=0.072
r98 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.0675 $X2=0.378 $Y2=0.0675
r99 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.378 $Y2=0.0675
.ends


* END of "./OAI322xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI322xp33_ASAP7_75t_L  VSS VDD B2 B1 A1 A2 A3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
M0 VSS N_B2_M0_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 noxref_10 N_B1_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_11 N_A1_M2_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_10 N_A2_M3_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_11 N_A3_M4_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 N_Y_M5_d N_C2_M5_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 noxref_11 N_C1_M6_g N_Y_M6_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_13 N_B2_M7_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M8 N_Y_M8_d N_B1_M8_g noxref_13 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M9 noxref_14 N_A1_M9_g N_Y_M9_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M10 noxref_15 N_A2_M10_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M11 VDD N_A3_M11_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M12 noxref_16 N_C2_M12_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341
+ $Y=0.189
M13 N_Y_M13_d N_C1_M13_g noxref_16 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.395 $Y=0.189
*
* 
* .include "OAI322xp33_ASAP7_75t_L.pex.sp.OAI322XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI322xp33_ASAP7_75t_L.pex.sp.OAI322XP33_ASAP7_75T_L.pxi"
* File: OAI322xp33_ASAP7_75t_L.pex.sp.OAI322XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:57:03 2017
* 
x_PM_OAI322XP33_ASAP7_75T_L%B2 N_B2_M0_g N_B2_c_2_p N_B2_M7_g B2 VSS
+ PM_OAI322XP33_ASAP7_75T_L%B2
x_PM_OAI322XP33_ASAP7_75T_L%B1 N_B1_M1_g N_B1_c_10_n N_B1_M8_g B1 VSS
+ PM_OAI322XP33_ASAP7_75T_L%B1
x_PM_OAI322XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_21_n N_A1_M9_g A1 VSS
+ PM_OAI322XP33_ASAP7_75T_L%A1
x_PM_OAI322XP33_ASAP7_75T_L%A2 N_A2_M3_g N_A2_c_34_n N_A2_M10_g A2 VSS
+ PM_OAI322XP33_ASAP7_75T_L%A2
x_PM_OAI322XP33_ASAP7_75T_L%A3 N_A3_M4_g N_A3_c_47_n N_A3_M11_g A3 VSS
+ PM_OAI322XP33_ASAP7_75T_L%A3
x_PM_OAI322XP33_ASAP7_75T_L%C2 N_C2_M5_g N_C2_c_59_n N_C2_M12_g C2 VSS
+ PM_OAI322XP33_ASAP7_75T_L%C2
x_PM_OAI322XP33_ASAP7_75T_L%C1 N_C1_M6_g N_C1_c_70_n N_C1_M13_g C1 VSS
+ PM_OAI322XP33_ASAP7_75T_L%C1
x_PM_OAI322XP33_ASAP7_75T_L%Y N_Y_M6_s N_Y_M5_d N_Y_c_102_n N_Y_M9_s N_Y_M8_d
+ N_Y_M13_d N_Y_c_91_n N_Y_c_79_n Y N_Y_c_80_n N_Y_c_83_n N_Y_c_99_n N_Y_c_85_n
+ N_Y_c_86_n N_Y_c_100_n N_Y_c_87_n N_Y_c_89_n N_Y_c_92_n N_Y_c_106_n
+ N_Y_c_101_n N_Y_c_94_n N_Y_c_111_n N_Y_c_96_n VSS PM_OAI322XP33_ASAP7_75T_L%Y
cc_1 N_B2_M0_g N_B1_M1_g 0.00323392f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_B2_c_2_p N_B1_c_10_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 B2 B1 0.00464555f $X=0.075 $Y=0.134 $X2=0.131 $Y2=0.134
cc_4 N_B2_M0_g N_A1_M2_g 2.69148e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 VSS N_B2_M0_g 3.62029e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_6 VSS B2 0.0012376f $X=0.075 $Y=0.134 $X2=0 $Y2=0
cc_7 B2 N_Y_c_79_n 4.85822e-19 $X=0.075 $Y=0.134 $X2=0 $Y2=0
cc_8 B2 N_Y_c_80_n 4.5241e-19 $X=0.075 $Y=0.134 $X2=0 $Y2=0
cc_9 N_B1_M1_g N_A1_M2_g 0.0036697f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_10 N_B1_c_10_n N_A1_c_21_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_11 B1 A1 0.00406615f $X=0.131 $Y=0.134 $X2=0.075 $Y2=0.134
cc_12 N_B1_M1_g N_A2_M3_g 3.09654e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_13 VSS N_B1_M1_g 3.62029e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_14 VSS B1 0.0012322f $X=0.131 $Y=0.134 $X2=0 $Y2=0
cc_15 B1 N_Y_c_79_n 0.00133251f $X=0.131 $Y=0.134 $X2=0 $Y2=0
cc_16 N_A1_M2_g N_A2_M3_g 0.00374235f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 N_A1_c_21_n N_A2_c_34_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_18 A1 A2 0.00483372f $X=0.187 $Y=0.136 $X2=0.081 $Y2=0.135
cc_19 N_A1_M2_g N_A3_M4_g 3.09654e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_20 VSS N_A1_M2_g 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_21 VSS A1 0.0012322f $X=0.187 $Y=0.136 $X2=0 $Y2=0
cc_22 A1 N_Y_c_79_n 0.0013295f $X=0.187 $Y=0.136 $X2=0 $Y2=0
cc_23 N_A1_M2_g N_Y_c_83_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 A1 N_Y_c_83_n 0.00124805f $X=0.187 $Y=0.136 $X2=0 $Y2=0
cc_25 N_A2_M3_g N_A3_M4_g 0.00372052f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_26 N_A2_c_34_n N_A3_c_47_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_27 A2 A3 0.00481191f $X=0.247 $Y=0.136 $X2=0 $Y2=0
cc_28 N_A2_M3_g N_C2_M5_g 2.74891e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_29 VSS N_A2_M3_g 2.68514e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_30 VSS A2 0.00121543f $X=0.247 $Y=0.136 $X2=0 $Y2=0
cc_31 VSS N_A2_M3_g 2.38303e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_32 A2 N_Y_c_85_n 0.00123064f $X=0.247 $Y=0.136 $X2=0 $Y2=0
cc_33 N_A2_M3_g N_Y_c_86_n 2.03357e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_34 N_A3_M4_g N_C2_M5_g 0.00335739f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_35 N_A3_c_47_n N_C2_c_59_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_36 A3 C2 0.00407268f $X=0.296 $Y=0.136 $X2=0.187 $Y2=0.136
cc_37 N_A3_M4_g N_C1_M6_g 2.74891e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_38 VSS N_A3_M4_g 3.45454e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_39 VSS A3 5.39731e-19 $X=0.296 $Y=0.136 $X2=0 $Y2=0
cc_40 N_A3_M4_g N_Y_c_87_n 2.64276e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_41 A3 N_Y_c_87_n 0.00124825f $X=0.296 $Y=0.136 $X2=0 $Y2=0
cc_42 N_C2_M5_g N_C1_M6_g 0.00372052f $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_43 N_C2_c_59_n N_C1_c_70_n 9.33263e-19 $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_44 C2 C1 0.00479746f $X=0.348 $Y=0.134 $X2=0.243 $Y2=0.135
cc_45 VSS N_C2_M5_g 3.55324e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_46 VSS C2 5.47169e-19 $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_47 N_C2_M5_g N_Y_c_89_n 2.64276e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_48 C2 N_Y_c_89_n 0.00124825f $X=0.348 $Y=0.134 $X2=0 $Y2=0
cc_49 VSS N_C1_M6_g 2.08515e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_50 C1 N_Y_c_91_n 3.87865e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_51 N_C1_M6_g N_Y_c_92_n 2.56935e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_52 C1 N_Y_c_92_n 0.00123064f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_53 N_C1_M6_g N_Y_c_94_n 2.76185e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_54 C1 N_Y_c_94_n 0.0012322f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_55 C1 N_Y_c_96_n 0.00440796f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_56 VSS N_Y_c_79_n 0.00139129f $X=0.162 $Y=0.0675 $X2=0 $Y2=0
cc_57 VSS N_Y_c_80_n 2.83966e-19 $X=0.1545 $Y=0.072 $X2=0 $Y2=0
cc_58 VSS N_Y_c_99_n 2.83966e-19 $X=0.202 $Y=0.072 $X2=0 $Y2=0
cc_59 VSS N_Y_c_100_n 2.83966e-19 $X=0.261 $Y=0.072 $X2=0 $Y2=0
cc_60 VSS N_Y_c_101_n 2.91395e-19 $X=0.27 $Y=0.072 $X2=0 $Y2=0
cc_61 VSS N_Y_c_102_n 0.00334511f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.135
cc_62 VSS N_Y_c_102_n 0.00373054f $X=0.432 $Y=0.036 $X2=0.189 $Y2=0.135
cc_63 VSS N_Y_c_102_n 0.00250965f $X=0.398 $Y=0.036 $X2=0.189 $Y2=0.135
cc_64 VSS N_Y_c_91_n 9.98826e-19 $X=0.432 $Y=0.036 $X2=0.189 $Y2=0.135
cc_65 VSS N_Y_c_106_n 2.47657e-19 $X=0.43 $Y=0.0675 $X2=0 $Y2=0
cc_66 VSS N_Y_c_106_n 0.00260156f $X=0.432 $Y=0.036 $X2=0 $Y2=0
cc_67 VSS N_Y_c_101_n 4.49388e-19 $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_68 VSS N_Y_c_101_n 0.00369159f $X=0.398 $Y=0.036 $X2=0 $Y2=0
cc_69 VSS N_Y_c_94_n 0.00369159f $X=0.432 $Y=0.036 $X2=0 $Y2=0
cc_70 VSS N_Y_c_111_n 3.84257e-19 $X=0.432 $Y=0.036 $X2=0 $Y2=0
cc_71 VSS N_Y_c_99_n 3.48201e-19 $X=0.234 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_72 VSS N_Y_c_100_n 3.19955e-19 $X=0.284 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./OAI322xp33_ASAP7_75t_L.pex.sp.OAI322XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI32xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:57:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI32xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI32xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI32xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:57:26 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI32XP33_ASAP7_75T_L%A1 2 5 7 12 15 17 VSS
c14 17 VSS 0.00717332f $X=0.066 $Y=0.0355
c15 15 VSS 0.00138151f $X=0.064 $Y=0.081
c16 14 VSS 8.66832e-19 $X=0.064 $Y=0.063
c17 12 VSS 0.00396218f $X=0.064 $Y=0.135
c18 5 VSS 0.00499815f $X=0.081 $Y=0.135
c19 2 VSS 0.0653824f $X=0.081 $Y=0.054
r20 17 19 0.528714 $w=4e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.053
+ $Y=0.0355 $X2=0.053 $Y2=0.045
r21 14 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.063 $X2=0.064 $Y2=0.081
r22 14 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.063 $X2=0.064 $Y2=0.045
r23 12 15 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.135 $X2=0.064 $Y2=0.081
r24 12 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r25 5 13 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r27 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI32XP33_ASAP7_75T_L%A2 2 5 7 10 12 20 VSS
c18 20 VSS 5.21467e-19 $X=0.135 $Y=0.1915
c19 12 VSS 8.8977e-19 $X=0.135 $Y=0.135
c20 10 VSS 5.14523e-19 $X=0.135 $Y=0.189
c21 5 VSS 0.00108083f $X=0.135 $Y=0.135
c22 2 VSS 0.0606055f $X=0.135 $Y=0.054
r23 10 20 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.135 $Y2=0.198
r24 10 12 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.135 $Y2=0.135
r25 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r27 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI32XP33_ASAP7_75T_L%A3 2 5 7 11 13 14 17 VSS
c16 17 VSS 0.001236f $X=0.187 $Y=0.0755
c17 14 VSS 1.11188e-19 $X=0.189 $Y=0.1205
c18 13 VSS 6.45073e-19 $X=0.189 $Y=0.106
c19 11 VSS 4.45217e-19 $X=0.189 $Y=0.135
c20 5 VSS 0.00107802f $X=0.189 $Y=0.135
c21 2 VSS 0.0604511f $X=0.189 $Y=0.054
r22 17 19 0.447408 $w=4.2e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.201
+ $Y=0.0755 $X2=0.201 $Y2=0.081
r23 13 14 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.106 $X2=0.189 $Y2=0.1205
r24 13 19 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.106 $X2=0.189 $Y2=0.081
r25 11 14 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.1205
r26 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r27 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI32XP33_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c11 10 VSS 9.97444e-19 $X=0.243 $Y=0.135
c12 5 VSS 0.00113686f $X=0.243 $Y=0.135
c13 2 VSS 0.0617155f $X=0.243 $Y=0.054
r14 10 14 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.1505
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI32XP33_ASAP7_75T_L%B2 2 5 7 10 VSS
c11 10 VSS 4.87963e-19 $X=0.298 $Y=0.1165
c12 5 VSS 0.00170409f $X=0.297 $Y=0.135
c13 2 VSS 0.066446f $X=0.297 $Y=0.054
r14 10 13 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1165 $X2=0.297 $Y2=0.135
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OAI32XP33_ASAP7_75T_L%Y 1 2 5 6 9 11 14 24 25 27 28 29 32 35 41 42 43
+ 48 52 VSS
c29 50 VSS 4.55454e-19 $X=0.351 $Y=0.216
c30 49 VSS 2.4939e-19 $X=0.351 $Y=0.207
c31 48 VSS 0.00419284f $X=0.351 $Y=0.2
c32 47 VSS 0.00132122f $X=0.351 $Y=0.106
c33 46 VSS 0.00381964f $X=0.351 $Y=0.225
c34 44 VSS 1.42799e-19 $X=0.34 $Y=0.072
c35 43 VSS 3.90732e-19 $X=0.338 $Y=0.072
c36 42 VSS 8.46035e-21 $X=0.306 $Y=0.072
c37 41 VSS 5.02599e-19 $X=0.288 $Y=0.072
c38 36 VSS 0.00199921f $X=0.342 $Y=0.072
c39 35 VSS 0.00146362f $X=0.306 $Y=0.234
c40 34 VSS 0.0030651f $X=0.288 $Y=0.234
c41 33 VSS 4.89341e-19 $X=0.256 $Y=0.234
c42 32 VSS 0.00142296f $X=0.252 $Y=0.234
c43 31 VSS 0.0024156f $X=0.234 $Y=0.234
c44 30 VSS 0.00455239f $X=0.222 $Y=0.234
c45 29 VSS 0.00146362f $X=0.198 $Y=0.234
c46 28 VSS 0.00338401f $X=0.18 $Y=0.234
c47 27 VSS 0.00340784f $X=0.144 $Y=0.234
c48 26 VSS 5.69744e-19 $X=0.104 $Y=0.234
c49 25 VSS 0.00236146f $X=0.099 $Y=0.234
c50 24 VSS 0.00373945f $X=0.073 $Y=0.234
c51 16 VSS 0.00364982f $X=0.342 $Y=0.234
c52 14 VSS 0.00345862f $X=0.322 $Y=0.216
c53 9 VSS 0.00346338f $X=0.056 $Y=0.2025
c54 6 VSS 5.01571e-19 $X=0.071 $Y=0.2025
c55 5 VSS 0.00220204f $X=0.27 $Y=0.054
c56 1 VSS 5.70405e-19 $X=0.287 $Y=0.054
r57 49 50 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.207 $X2=0.351 $Y2=0.216
r58 48 49 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.2 $X2=0.351 $Y2=0.207
r59 47 48 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.106 $X2=0.351 $Y2=0.2
r60 46 52 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.234
r61 46 50 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.216
r62 45 47 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.106
r63 43 44 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.072 $X2=0.34 $Y2=0.072
r64 42 43 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.072 $X2=0.338 $Y2=0.072
r65 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.306 $Y2=0.072
r66 38 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.072 $X2=0.288 $Y2=0.072
r67 36 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.072 $X2=0.351 $Y2=0.081
r68 36 44 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.072 $X2=0.34 $Y2=0.072
r69 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r70 33 34 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.234 $X2=0.288 $Y2=0.234
r71 32 33 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.256 $Y2=0.234
r72 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r73 30 31 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.222
+ $Y=0.234 $X2=0.234 $Y2=0.234
r74 29 30 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.222 $Y2=0.234
r75 28 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r76 27 28 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.18 $Y2=0.234
r77 26 27 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.104
+ $Y=0.234 $X2=0.144 $Y2=0.234
r78 25 26 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.234 $X2=0.104 $Y2=0.234
r79 24 25 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.073
+ $Y=0.234 $X2=0.099 $Y2=0.234
r80 22 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.306 $Y2=0.234
r81 18 24 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.073 $Y2=0.234
r82 16 52 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.351 $Y2=0.234
r83 16 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.324 $Y2=0.234
r84 14 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r85 11 14 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.216 $X2=0.322 $Y2=0.216
r86 9 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r87 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
r88 5 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.072 $X2=0.27
+ $Y2=0.072
r89 2 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.054 $X2=0.27 $Y2=0.054
r90 1 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.054 $X2=0.27 $Y2=0.054
.ends


* END of "./OAI32xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI32xp33_ASAP7_75t_L  VSS VDD A1 A2 A3 B1 B2 Y
* 
* Y	Y
* B2	B2
* B1	B1
* A3	A3
* A2	A2
* A1	A1
M0 noxref_8 N_A1_M0_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 VSS N_A2_M1_g noxref_8 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 noxref_8 N_A3_M2_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.027
M3 N_Y_M3_d N_B1_M3_g noxref_8 VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 noxref_8 N_B2_M4_g N_Y_M4_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.027
M5 noxref_10 N_A1_M5_g N_Y_M5_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M6 noxref_11 N_A2_M6_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 VDD N_A3_M7_g noxref_11 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M8 noxref_12 N_B1_M8_g VDD VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M9 N_Y_M9_d N_B2_M9_g noxref_12 VDD PMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.189
*
* 
* .include "OAI32xp33_ASAP7_75t_L.pex.sp.OAI32XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI32xp33_ASAP7_75t_L.pex.sp.OAI32XP33_ASAP7_75T_L.pxi"
* File: OAI32xp33_ASAP7_75t_L.pex.sp.OAI32XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:57:26 2017
* 
x_PM_OAI32XP33_ASAP7_75T_L%A1 N_A1_M0_g N_A1_c_2_p N_A1_M5_g N_A1_c_3_p
+ N_A1_c_4_p A1 VSS PM_OAI32XP33_ASAP7_75T_L%A1
x_PM_OAI32XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_16_n N_A2_M6_g N_A2_c_17_n
+ N_A2_c_18_n A2 VSS PM_OAI32XP33_ASAP7_75T_L%A2
x_PM_OAI32XP33_ASAP7_75T_L%A3 N_A3_M2_g N_A3_c_35_n N_A3_M7_g N_A3_c_47_p
+ N_A3_c_36_n N_A3_c_37_n A3 VSS PM_OAI32XP33_ASAP7_75T_L%A3
x_PM_OAI32XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_51_n N_B1_M8_g N_B1_c_52_n B1 VSS
+ PM_OAI32XP33_ASAP7_75T_L%B1
x_PM_OAI32XP33_ASAP7_75T_L%B2 N_B2_M4_g N_B2_c_62_n N_B2_M9_g B2 VSS
+ PM_OAI32XP33_ASAP7_75T_L%B2
x_PM_OAI32XP33_ASAP7_75T_L%Y N_Y_M4_s N_Y_M3_d N_Y_c_91_n N_Y_M5_s N_Y_c_72_n
+ N_Y_M9_d N_Y_c_85_n N_Y_c_74_n N_Y_c_75_n N_Y_c_78_n N_Y_c_99_p N_Y_c_80_n
+ N_Y_c_83_n N_Y_c_86_n N_Y_c_82_n N_Y_c_88_n N_Y_c_97_n N_Y_c_90_n Y VSS
+ PM_OAI32XP33_ASAP7_75T_L%Y
cc_1 N_A1_M0_g N_A2_M1_g 0.00354623f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A1_c_2_p N_A2_c_16_n 0.00104216f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p N_A2_c_17_n 0.00336701f $X=0.064 $Y=0.135 $X2=0.135 $Y2=0.189
cc_4 N_A1_c_4_p N_A2_c_18_n 7.95431e-19 $X=0.064 $Y=0.081 $X2=0.135 $Y2=0.135
cc_5 N_A1_c_3_p A2 0.00125891f $X=0.064 $Y=0.135 $X2=0.135 $Y2=0.1915
cc_6 N_A1_M0_g N_A3_M2_g 2.69148e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_7 VSS A1 8.09309e-19 $X=0.066 $Y=0.0355 $X2=0.135 $Y2=0.135
cc_8 VSS A1 0.00128996f $X=0.066 $Y=0.0355 $X2=0 $Y2=0
cc_9 N_A1_c_3_p N_Y_M5_s 2.00679e-19 $X=0.064 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_10 N_A1_c_2_p N_Y_c_72_n 4.59187e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 N_A1_c_3_p N_Y_c_72_n 0.00485527f $X=0.064 $Y=0.135 $X2=0 $Y2=0
cc_12 N_A1_c_3_p N_Y_c_74_n 0.00305998f $X=0.064 $Y=0.135 $X2=0 $Y2=0
cc_13 N_A1_M0_g N_Y_c_75_n 2.39633e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_14 N_A1_c_2_p N_Y_c_75_n 2.93604e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_15 N_A2_M1_g N_A3_M2_g 0.00323392f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_16 N_A2_c_16_n N_A3_c_35_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_17 N_A2_c_17_n N_A3_c_36_n 0.00216429f $X=0.135 $Y=0.189 $X2=0.064 $Y2=0.135
cc_18 A2 N_A3_c_37_n 0.00216429f $X=0.135 $Y=0.1915 $X2=0.064 $Y2=0.063
cc_19 N_A2_c_18_n A3 0.00216429f $X=0.135 $Y=0.135 $X2=0.066 $Y2=0.0355
cc_20 N_A2_M1_g N_B1_M3_g 2.34385e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_21 VSS N_A2_c_18_n 0.00211795f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 VSS N_A2_c_18_n 0.00412802f $X=0.135 $Y=0.135 $X2=0.066 $Y2=0.0355
cc_23 VSS N_A2_M1_g 2.34993e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_24 A2 N_Y_c_72_n 2.39233e-19 $X=0.135 $Y=0.1915 $X2=0.064 $Y2=0.045
cc_25 N_A2_M1_g N_Y_c_78_n 3.27325e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_26 A2 N_Y_c_78_n 0.00424732f $X=0.135 $Y=0.1915 $X2=0 $Y2=0
cc_27 VSS A2 2.99671e-19 $X=0.135 $Y=0.1915 $X2=0.081 $Y2=0.054
cc_28 N_A3_M2_g N_B1_M3_g 0.00323392f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_29 N_A3_c_35_n N_B1_c_51_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_30 N_A3_c_37_n N_B1_c_52_n 0.00383317f $X=0.189 $Y=0.1205 $X2=0 $Y2=0
cc_31 N_A3_M2_g N_B2_M4_g 2.69148e-19 $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_32 VSS A3 0.00222856f $X=0.187 $Y=0.0755 $X2=0 $Y2=0
cc_33 VSS N_A3_M2_g 2.34993e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_34 VSS A3 0.00413281f $X=0.187 $Y=0.0755 $X2=0 $Y2=0
cc_35 N_A3_M2_g N_Y_c_80_n 2.64276e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_36 N_A3_c_47_p N_Y_c_80_n 0.00125427f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_37 A3 N_Y_c_82_n 7.98429e-19 $X=0.187 $Y=0.0755 $X2=0 $Y2=0
cc_38 N_B1_M3_g N_B2_M4_g 0.0036697f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_39 N_B1_c_51_n N_B2_c_62_n 9.33263e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_40 N_B1_c_52_n B2 0.00487321f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.189
cc_41 VSS N_B1_M3_g 3.47199e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_42 VSS N_B1_c_52_n 5.30079e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_43 N_B1_M3_g N_Y_c_83_n 2.56935e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_44 N_B1_c_52_n N_Y_c_83_n 0.00123064f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_45 VSS N_B2_M4_g 2.38303e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_46 B2 N_Y_c_85_n 3.87865e-19 $X=0.298 $Y=0.1165 $X2=0.189 $Y2=0.1205
cc_47 N_B2_M4_g N_Y_c_86_n 2.64276e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_48 B2 N_Y_c_86_n 0.00124805f $X=0.298 $Y=0.1165 $X2=0 $Y2=0
cc_49 N_B2_M4_g N_Y_c_88_n 2.76185e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_50 B2 N_Y_c_88_n 0.0012322f $X=0.298 $Y=0.1165 $X2=0 $Y2=0
cc_51 B2 N_Y_c_90_n 0.00446403f $X=0.298 $Y=0.1165 $X2=0 $Y2=0
cc_52 VSS N_Y_c_91_n 0.00288888f $X=0.216 $Y=0.054 $X2=0.081 $Y2=0.135
cc_53 VSS N_Y_c_91_n 0.00302498f $X=0.322 $Y=0.054 $X2=0.081 $Y2=0.135
cc_54 VSS N_Y_c_91_n 0.00250965f $X=0.324 $Y=0.036 $X2=0.081 $Y2=0.135
cc_55 VSS N_Y_c_85_n 4.54531e-19 $X=0.322 $Y=0.054 $X2=0.064 $Y2=0.063
cc_56 VSS N_Y_c_82_n 2.56435e-19 $X=0.216 $Y=0.054 $X2=0 $Y2=0
cc_57 VSS N_Y_c_82_n 0.00705732f $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_58 VSS N_Y_c_97_n 0.00391824f $X=0.322 $Y=0.054 $X2=0 $Y2=0
cc_59 VSS N_Y_c_75_n 2.48104e-19 $X=0.099 $Y=0.234 $X2=0.081 $Y2=0.054
cc_60 VSS N_Y_c_99_p 4.8755e-19 $X=0.18 $Y=0.234 $X2=0.081 $Y2=0.054

* END of "./OAI32xp33_ASAP7_75t_L.pex.sp.OAI32XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI331xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:57:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI331xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI331xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI331xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:57:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI331XP33_ASAP7_75T_L%A3 2 5 7 10 14 VSS
c4 10 VSS 0.00613146f $X=0.081 $Y=0.135
c5 5 VSS 0.00238289f $X=0.081 $Y=0.135
c6 2 VSS 0.062704f $X=0.081 $Y=0.0675
r7 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.155
r8 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r9 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r10 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI331XP33_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c11 14 VSS 0.00132043f $X=0.135 $Y=0.155
c12 10 VSS 4.26629e-19 $X=0.135 $Y=0.135
c13 5 VSS 0.00123757f $X=0.135 $Y=0.135
c14 2 VSS 0.0598541f $X=0.135 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI331XP33_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c11 10 VSS 0.00101969f $X=0.189 $Y=0.135
c12 5 VSS 0.00121257f $X=0.189 $Y=0.135
c13 2 VSS 0.0608354f $X=0.189 $Y=0.0675
r14 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI331XP33_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.243 $Y=0.135
c14 5 VSS 0.00111336f $X=0.243 $Y=0.135
c15 2 VSS 0.0617786f $X=0.243 $Y=0.0675
r16 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.154
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI331XP33_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.297 $Y=0.135
c14 5 VSS 0.00112198f $X=0.297 $Y=0.135
c15 2 VSS 0.0616432f $X=0.297 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OAI331XP33_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c11 10 VSS 7.24259e-19 $X=0.351 $Y=0.135
c12 5 VSS 0.00113686f $X=0.351 $Y=0.135
c13 2 VSS 0.0618011f $X=0.351 $Y=0.0675
r14 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OAI331XP33_ASAP7_75T_L%C1 2 5 7 10 14 VSS
c8 10 VSS 0.00201948f $X=0.405 $Y=0.135
c9 5 VSS 0.00178636f $X=0.405 $Y=0.135
c10 2 VSS 0.0660367f $X=0.405 $Y=0.0675
r11 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.155
r12 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OAI331XP33_ASAP7_75T_L%Y 1 4 6 7 10 11 14 24 25 26 27 28 30 33 39 41
+ 49 VSS
c24 49 VSS 0.00190266f $X=0.45 $Y=0.072
c25 48 VSS 0.00163302f $X=0.459 $Y=0.072
c26 43 VSS 4.139e-19 $X=0.459 $Y=0.2125
c27 41 VSS 8.61055e-19 $X=0.459 $Y=0.1245
c28 40 VSS 0.00103118f $X=0.459 $Y=0.106
c29 39 VSS 0.00322429f $X=0.458 $Y=0.143
c30 37 VSS 3.97344e-19 $X=0.459 $Y=0.225
c31 35 VSS 6.94247e-19 $X=0.4245 $Y=0.234
c32 34 VSS 2.39163e-19 $X=0.417 $Y=0.234
c33 33 VSS 0.00146362f $X=0.414 $Y=0.234
c34 32 VSS 2.39163e-19 $X=0.396 $Y=0.234
c35 31 VSS 0.00617212f $X=0.393 $Y=0.234
c36 30 VSS 0.00142296f $X=0.36 $Y=0.234
c37 29 VSS 3.71649e-19 $X=0.342 $Y=0.234
c38 28 VSS 0.00311761f $X=0.339 $Y=0.234
c39 27 VSS 0.00146362f $X=0.306 $Y=0.234
c40 26 VSS 0.00340162f $X=0.288 $Y=0.234
c41 25 VSS 0.00146362f $X=0.252 $Y=0.234
c42 24 VSS 0.00417843f $X=0.234 $Y=0.234
c43 16 VSS 0.00591242f $X=0.45 $Y=0.234
c44 14 VSS 0.00701741f $X=0.43 $Y=0.2025
c45 10 VSS 0.00220422f $X=0.216 $Y=0.2025
c46 6 VSS 5.61153e-19 $X=0.233 $Y=0.2025
c47 4 VSS 0.0013176f $X=0.43 $Y=0.0675
r48 49 50 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.072 $X2=0.4545 $Y2=0.072
r49 48 50 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.072 $X2=0.4545 $Y2=0.072
r50 45 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.072 $X2=0.45 $Y2=0.072
r51 42 43 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.2 $X2=0.459 $Y2=0.2125
r52 40 41 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.106 $X2=0.459 $Y2=0.1245
r53 39 42 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.143 $X2=0.459 $Y2=0.2
r54 39 41 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.143 $X2=0.459 $Y2=0.1245
r55 37 43 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.2125
r56 36 48 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.072
r57 36 40 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.106
r58 34 35 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.417
+ $Y=0.234 $X2=0.4245 $Y2=0.234
r59 33 34 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.417 $Y2=0.234
r60 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r61 31 32 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.393
+ $Y=0.234 $X2=0.396 $Y2=0.234
r62 30 31 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.393 $Y2=0.234
r63 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r64 28 29 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.339
+ $Y=0.234 $X2=0.342 $Y2=0.234
r65 27 28 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.339 $Y2=0.234
r66 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r67 25 26 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.288 $Y2=0.234
r68 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r69 22 35 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.4245 $Y2=0.234
r70 18 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.234 $Y2=0.234
r71 16 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r72 16 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.432 $Y2=0.234
r73 14 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r74 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.43 $Y2=0.2025
r75 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r76 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r77 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r78 4 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.072 $X2=0.432
+ $Y2=0.072
r79 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.43 $Y2=0.0675
.ends


* END of "./OAI331xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI331xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C1 Y
* 
* Y	Y
* C1	C1
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 noxref_10 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_A2_M1_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_10 N_A1_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_11 N_B1_M3_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_10 N_B2_M4_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_11 N_B3_M5_g noxref_10 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 N_Y_M6_d N_C1_M6_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_13 N_A3_M7_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M8 noxref_14 N_A2_M8_g noxref_13 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M9 N_Y_M9_d N_A1_M9_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M10 noxref_15 N_B1_M10_g N_Y_M10_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M11 noxref_16 N_B2_M11_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M12 VDD N_B3_M12_g noxref_16 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M13 N_Y_M13_d N_C1_M13_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
*
* 
* .include "OAI331xp33_ASAP7_75t_L.pex.sp.OAI331XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI331xp33_ASAP7_75t_L.pex.sp.OAI331XP33_ASAP7_75T_L.pxi"
* File: OAI331xp33_ASAP7_75t_L.pex.sp.OAI331XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:57:48 2017
* 
x_PM_OAI331XP33_ASAP7_75T_L%A3 N_A3_M0_g N_A3_c_2_p N_A3_M7_g N_A3_c_3_p A3 VSS
+ PM_OAI331XP33_ASAP7_75T_L%A3
x_PM_OAI331XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_6_n N_A2_M8_g N_A2_c_7_n A2 VSS
+ PM_OAI331XP33_ASAP7_75T_L%A2
x_PM_OAI331XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_18_n N_A1_M9_g N_A1_c_19_n A1
+ VSS PM_OAI331XP33_ASAP7_75T_L%A1
x_PM_OAI331XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_29_n N_B1_M10_g N_B1_c_30_n B1
+ VSS PM_OAI331XP33_ASAP7_75T_L%B1
x_PM_OAI331XP33_ASAP7_75T_L%B2 N_B2_M4_g N_B2_c_42_n N_B2_M11_g N_B2_c_43_n B2
+ VSS PM_OAI331XP33_ASAP7_75T_L%B2
x_PM_OAI331XP33_ASAP7_75T_L%B3 N_B3_M5_g N_B3_c_55_n N_B3_M12_g N_B3_c_56_n B3
+ VSS PM_OAI331XP33_ASAP7_75T_L%B3
x_PM_OAI331XP33_ASAP7_75T_L%C1 N_C1_M6_g N_C1_c_66_n N_C1_M13_g N_C1_c_67_n C1
+ VSS PM_OAI331XP33_ASAP7_75T_L%C1
x_PM_OAI331XP33_ASAP7_75T_L%Y N_Y_M6_d N_Y_c_91_n N_Y_M10_s N_Y_M9_d N_Y_c_72_n
+ N_Y_M13_d N_Y_c_82_n N_Y_c_73_n N_Y_c_76_n N_Y_c_88_n N_Y_c_78_n N_Y_c_89_n
+ N_Y_c_80_n N_Y_c_83_n Y N_Y_c_85_n N_Y_c_90_n VSS PM_OAI331XP33_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_A2_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A3_c_2_p N_A2_c_6_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A3_c_3_p N_A2_c_7_n 0.00653171f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A3_M0_g N_A1_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 N_A2_M1_g N_A1_M2_g 0.00327995f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_6 N_A2_c_6_n N_A1_c_18_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_7 N_A2_c_7_n N_A1_c_19_n 0.00466039f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_8 N_A2_M1_g N_B1_M3_g 2.71887e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_9 VSS N_A2_M1_g 3.62029e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_10 VSS N_A2_c_7_n 0.0012376f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_11 A2 N_Y_c_72_n 5.87506e-19 $X=0.135 $Y=0.155 $X2=0.081 $Y2=0.135
cc_12 A2 N_Y_c_73_n 4.59602e-19 $X=0.135 $Y=0.155 $X2=0 $Y2=0
cc_13 N_A1_M2_g N_B1_M3_g 0.0036939f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_A1_c_18_n N_B1_c_29_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 N_A1_c_19_n N_B1_c_30_n 0.00406615f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_16 N_A1_M2_g N_B2_M4_g 3.06651e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 VSS N_A1_M2_g 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_18 VSS N_A1_c_19_n 0.0012322f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_19 N_A1_c_19_n N_Y_c_72_n 0.0013295f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_20 N_B1_M3_g N_B2_M4_g 0.00371573f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_21 N_B1_c_29_n N_B2_c_42_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_22 N_B1_c_30_n N_B2_c_43_n 0.00483372f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_23 N_B1_M3_g N_B3_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_24 VSS N_B1_M3_g 3.62029e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_25 VSS N_B1_c_30_n 0.0012322f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_26 N_B1_c_30_n N_Y_c_72_n 0.0013295f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_27 N_B1_M3_g N_Y_c_76_n 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_28 N_B1_c_30_n N_Y_c_76_n 0.00124805f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_29 N_B2_M4_g N_B3_M5_g 0.0036939f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_30 N_B2_c_42_n N_B3_c_55_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_31 N_B2_c_43_n N_B3_c_56_n 0.00483372f $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_32 N_B2_M4_g N_C1_M6_g 2.71887e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_33 VSS N_B2_M4_g 2.68514e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_34 VSS N_B2_c_43_n 0.00121543f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_35 VSS N_B2_M4_g 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B2_M4_g N_Y_c_78_n 3.48613e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_B2_c_43_n N_Y_c_78_n 0.00124805f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_38 N_B3_M5_g N_C1_M6_g 0.00333077f $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_39 N_B3_c_55_n N_C1_c_66_n 9.33263e-19 $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_40 N_B3_c_56_n N_C1_c_67_n 0.00406322f $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_41 VSS N_B3_M5_g 3.47199e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_42 VSS N_B3_c_56_n 5.30079e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_43 N_B3_M5_g N_Y_c_80_n 2.56935e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_B3_c_56_n N_Y_c_80_n 0.00123064f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_45 N_C1_c_67_n N_Y_c_82_n 0.00114532f $X=0.405 $Y=0.135 $X2=0.296 $Y2=0.155
cc_46 N_C1_M6_g N_Y_c_83_n 2.64276e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_C1_c_67_n N_Y_c_83_n 0.00124805f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_48 N_C1_c_67_n N_Y_c_85_n 0.00391301f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_49 VSS N_Y_c_72_n 0.00138157f $X=0.216 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_50 VSS N_Y_c_73_n 2.88662e-19 $X=0.2085 $Y=0.072 $X2=0 $Y2=0
cc_51 VSS N_Y_c_88_n 2.88662e-19 $X=0.254 $Y=0.072 $X2=0 $Y2=0
cc_52 VSS N_Y_c_89_n 2.88662e-19 $X=0.315 $Y=0.072 $X2=0 $Y2=0
cc_53 VSS N_Y_c_90_n 2.83845e-19 $X=0.324 $Y=0.072 $X2=0 $Y2=0
cc_54 VSS N_Y_c_91_n 3.11523e-19 $X=0.378 $Y=0.036 $X2=0.243 $Y2=0.135
cc_55 VSS N_Y_c_91_n 0.00333695f $X=0.378 $Y=0.036 $X2=0.243 $Y2=0.135
cc_56 VSS N_Y_c_90_n 4.47506e-19 $X=0.378 $Y=0.036 $X2=0 $Y2=0
cc_57 VSS N_Y_c_88_n 3.48201e-19 $X=0.288 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_58 VSS N_Y_c_89_n 3.30547e-19 $X=0.339 $Y=0.234 $X2=0.135 $Y2=0.0675

* END of "./OAI331xp33_ASAP7_75t_L.pex.sp.OAI331XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI332xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:58:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI332xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI332xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI332xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:58:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI332XP33_ASAP7_75T_L%A3 2 5 7 10 14 VSS
c4 10 VSS 0.00613146f $X=0.081 $Y=0.135
c5 5 VSS 0.00238289f $X=0.081 $Y=0.135
c6 2 VSS 0.062704f $X=0.081 $Y=0.0675
r7 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.155
r8 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r9 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r10 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI332XP33_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c11 14 VSS 0.00132043f $X=0.135 $Y=0.155
c12 10 VSS 4.26629e-19 $X=0.135 $Y=0.135
c13 5 VSS 0.00123757f $X=0.135 $Y=0.135
c14 2 VSS 0.0598541f $X=0.135 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI332XP33_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c11 10 VSS 0.00101969f $X=0.189 $Y=0.135
c12 5 VSS 0.00121257f $X=0.189 $Y=0.135
c13 2 VSS 0.0608354f $X=0.189 $Y=0.0675
r14 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI332XP33_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.243 $Y=0.135
c14 5 VSS 0.00111336f $X=0.243 $Y=0.135
c15 2 VSS 0.0617786f $X=0.243 $Y=0.0675
r16 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.154
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI332XP33_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.297 $Y=0.135
c14 5 VSS 0.00112198f $X=0.297 $Y=0.135
c15 2 VSS 0.0616432f $X=0.297 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OAI332XP33_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c12 10 VSS 7.27237e-19 $X=0.351 $Y=0.135
c13 5 VSS 0.00111185f $X=0.351 $Y=0.135
c14 2 VSS 0.0615515f $X=0.351 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OAI332XP33_ASAP7_75T_L%C2 2 5 7 10 14 VSS
c11 10 VSS 0.00167719f $X=0.405 $Y=0.135
c12 5 VSS 0.00113407f $X=0.405 $Y=0.135
c13 2 VSS 0.0618699f $X=0.405 $Y=0.0675
r14 10 14 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.156
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OAI332XP33_ASAP7_75T_L%C1 2 5 7 10 14 VSS
c11 10 VSS 4.90626e-19 $X=0.459 $Y=0.135
c12 5 VSS 0.00170346f $X=0.459 $Y=0.135
c13 2 VSS 0.0662985f $X=0.459 $Y=0.0675
r14 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OAI332XP33_ASAP7_75T_L%Y 1 2 5 6 7 10 11 14 24 25 26 27 28 30 32 34
+ 35 41 42 43 48 49 50 VSS
c36 52 VSS 5.10117e-19 $X=0.513 $Y=0.2125
c37 50 VSS 8.61055e-19 $X=0.513 $Y=0.1245
c38 49 VSS 0.00112176f $X=0.513 $Y=0.106
c39 48 VSS 0.00322429f $X=0.512 $Y=0.143
c40 46 VSS 6.07272e-19 $X=0.513 $Y=0.225
c41 44 VSS 4.93718e-20 $X=0.503 $Y=0.072
c42 43 VSS 4.1269e-19 $X=0.502 $Y=0.072
c43 42 VSS 8.46035e-21 $X=0.468 $Y=0.072
c44 41 VSS 4.70878e-19 $X=0.45 $Y=0.072
c45 36 VSS 0.0019286f $X=0.504 $Y=0.072
c46 35 VSS 0.00146362f $X=0.468 $Y=0.234
c47 34 VSS 0.00296425f $X=0.45 $Y=0.234
c48 33 VSS 3.35992e-19 $X=0.417 $Y=0.234
c49 32 VSS 0.00142296f $X=0.414 $Y=0.234
c50 31 VSS 0.00672869f $X=0.396 $Y=0.234
c51 30 VSS 0.00142296f $X=0.36 $Y=0.234
c52 29 VSS 3.35992e-19 $X=0.342 $Y=0.234
c53 28 VSS 0.00311761f $X=0.339 $Y=0.234
c54 27 VSS 0.00146362f $X=0.306 $Y=0.234
c55 26 VSS 0.00340162f $X=0.288 $Y=0.234
c56 25 VSS 0.00146362f $X=0.252 $Y=0.234
c57 24 VSS 0.00418453f $X=0.234 $Y=0.234
c58 16 VSS 0.00700674f $X=0.504 $Y=0.234
c59 14 VSS 0.0038436f $X=0.484 $Y=0.2025
c60 10 VSS 0.00220422f $X=0.216 $Y=0.2025
c61 6 VSS 5.61153e-19 $X=0.233 $Y=0.2025
c62 5 VSS 0.0023085f $X=0.432 $Y=0.0675
c63 1 VSS 5.70099e-19 $X=0.449 $Y=0.0675
r64 51 52 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.2 $X2=0.513 $Y2=0.2125
r65 49 50 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.106 $X2=0.513 $Y2=0.1245
r66 48 51 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.143 $X2=0.513 $Y2=0.2
r67 48 50 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.143 $X2=0.513 $Y2=0.1245
r68 46 52 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.2125
r69 45 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.081 $X2=0.513 $Y2=0.106
r70 43 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.502
+ $Y=0.072 $X2=0.503 $Y2=0.072
r71 42 43 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.072 $X2=0.502 $Y2=0.072
r72 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.072 $X2=0.468 $Y2=0.072
r73 38 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.072 $X2=0.45 $Y2=0.072
r74 36 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.072 $X2=0.513 $Y2=0.081
r75 36 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.072 $X2=0.503 $Y2=0.072
r76 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r77 33 34 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.417
+ $Y=0.234 $X2=0.45 $Y2=0.234
r78 32 33 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.417 $Y2=0.234
r79 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r80 30 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.396 $Y2=0.234
r81 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r82 28 29 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.339
+ $Y=0.234 $X2=0.342 $Y2=0.234
r83 27 28 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.339 $Y2=0.234
r84 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r85 25 26 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.288 $Y2=0.234
r86 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r87 22 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.468 $Y2=0.234
r88 18 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.234 $Y2=0.234
r89 16 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.234 $X2=0.513 $Y2=0.225
r90 16 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.486 $Y2=0.234
r91 14 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r92 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.484 $Y2=0.2025
r93 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r94 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r95 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r96 5 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.072 $X2=0.432
+ $Y2=0.072
r97 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.432 $Y2=0.0675
r98 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.449
+ $Y=0.0675 $X2=0.432 $Y2=0.0675
.ends


* END of "./OAI332xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI332xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 noxref_11 N_A3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_A2_M1_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_11 N_A1_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_12 N_B1_M3_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_11 N_B2_M4_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_12 N_B3_M5_g noxref_11 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 N_Y_M6_d N_C2_M6_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_12 N_C1_M7_g N_Y_M7_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 noxref_14 N_A3_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M9 noxref_15 N_A2_M9_g noxref_14 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M10 N_Y_M10_d N_A1_M10_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.179 $Y=0.162
M11 noxref_16 N_B1_M11_g N_Y_M11_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M12 noxref_17 N_B2_M12_g noxref_16 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M13 VDD N_B3_M13_g noxref_17 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M14 noxref_18 N_C2_M14_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M15 N_Y_M15_d N_C1_M15_g noxref_18 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
*
* 
* .include "OAI332xp33_ASAP7_75t_L.pex.sp.OAI332XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI332xp33_ASAP7_75t_L.pex.sp.OAI332XP33_ASAP7_75T_L.pxi"
* File: OAI332xp33_ASAP7_75t_L.pex.sp.OAI332XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:58:11 2017
* 
x_PM_OAI332XP33_ASAP7_75T_L%A3 N_A3_M0_g N_A3_c_2_p N_A3_M8_g N_A3_c_3_p A3 VSS
+ PM_OAI332XP33_ASAP7_75T_L%A3
x_PM_OAI332XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_6_n N_A2_M9_g N_A2_c_7_n A2 VSS
+ PM_OAI332XP33_ASAP7_75T_L%A2
x_PM_OAI332XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_18_n N_A1_M10_g N_A1_c_19_n A1
+ VSS PM_OAI332XP33_ASAP7_75T_L%A1
x_PM_OAI332XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_29_n N_B1_M11_g N_B1_c_30_n B1
+ VSS PM_OAI332XP33_ASAP7_75T_L%B1
x_PM_OAI332XP33_ASAP7_75T_L%B2 N_B2_M4_g N_B2_c_42_n N_B2_M12_g N_B2_c_43_n B2
+ VSS PM_OAI332XP33_ASAP7_75T_L%B2
x_PM_OAI332XP33_ASAP7_75T_L%B3 N_B3_M5_g N_B3_c_55_n N_B3_M13_g N_B3_c_56_n B3
+ VSS PM_OAI332XP33_ASAP7_75T_L%B3
x_PM_OAI332XP33_ASAP7_75T_L%C2 N_C2_M6_g N_C2_c_67_n N_C2_M14_g N_C2_c_68_n C2
+ VSS PM_OAI332XP33_ASAP7_75T_L%C2
x_PM_OAI332XP33_ASAP7_75T_L%C1 N_C1_M7_g N_C1_c_78_n N_C1_M15_g N_C1_c_79_n C1
+ VSS PM_OAI332XP33_ASAP7_75T_L%C1
x_PM_OAI332XP33_ASAP7_75T_L%Y N_Y_M7_s N_Y_M6_d N_Y_c_110_n N_Y_M11_s N_Y_M10_d
+ N_Y_c_87_n N_Y_M15_d N_Y_c_99_n N_Y_c_88_n N_Y_c_91_n N_Y_c_107_n N_Y_c_93_n
+ N_Y_c_108_n N_Y_c_95_n N_Y_c_97_n N_Y_c_122_p N_Y_c_100_n N_Y_c_109_n
+ N_Y_c_102_n N_Y_c_117_n Y N_Y_c_119_n N_Y_c_104_n VSS
+ PM_OAI332XP33_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_A2_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A3_c_2_p N_A2_c_6_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A3_c_3_p N_A2_c_7_n 0.00653171f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A3_M0_g N_A1_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 N_A2_M1_g N_A1_M2_g 0.00327995f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_6 N_A2_c_6_n N_A1_c_18_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_7 N_A2_c_7_n N_A1_c_19_n 0.00466039f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_8 N_A2_M1_g N_B1_M3_g 2.71887e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_9 VSS N_A2_M1_g 3.62029e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_10 VSS N_A2_c_7_n 0.0012376f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_11 A2 N_Y_c_87_n 5.87506e-19 $X=0.135 $Y=0.155 $X2=0.081 $Y2=0.135
cc_12 A2 N_Y_c_88_n 4.59821e-19 $X=0.135 $Y=0.155 $X2=0 $Y2=0
cc_13 N_A1_M2_g N_B1_M3_g 0.0036939f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_A1_c_18_n N_B1_c_29_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 N_A1_c_19_n N_B1_c_30_n 0.00406615f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_16 N_A1_M2_g N_B2_M4_g 3.06651e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 VSS N_A1_M2_g 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_18 VSS N_A1_c_19_n 0.0012322f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_19 N_A1_c_19_n N_Y_c_87_n 0.0013295f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_20 N_B1_M3_g N_B2_M4_g 0.00371573f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_21 N_B1_c_29_n N_B2_c_42_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_22 N_B1_c_30_n N_B2_c_43_n 0.00483372f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_23 N_B1_M3_g N_B3_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_24 VSS N_B1_M3_g 3.62029e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_25 VSS N_B1_c_30_n 0.0012322f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_26 N_B1_c_30_n N_Y_c_87_n 0.0013295f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_27 N_B1_M3_g N_Y_c_91_n 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_28 N_B1_c_30_n N_Y_c_91_n 0.00124805f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_29 N_B2_M4_g N_B3_M5_g 0.0036939f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_30 N_B2_c_42_n N_B3_c_55_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_31 N_B2_c_43_n N_B3_c_56_n 0.00483372f $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_32 N_B2_M4_g N_C2_M6_g 2.71887e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_33 VSS N_B2_M4_g 2.68514e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_34 VSS N_B2_c_43_n 0.00121543f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_35 VSS N_B2_M4_g 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B2_M4_g N_Y_c_93_n 3.48613e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_B2_c_43_n N_Y_c_93_n 0.00124805f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_38 N_B3_M5_g N_C2_M6_g 0.00333077f $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_39 N_B3_c_55_n N_C2_c_67_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_40 N_B3_c_56_n N_C2_c_68_n 0.00406615f $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_41 N_B3_M5_g N_C1_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_42 VSS N_B3_M5_g 3.47199e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_43 VSS N_B3_c_56_n 5.30079e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_44 N_B3_M5_g N_Y_c_95_n 2.56935e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_45 N_B3_c_56_n N_Y_c_95_n 0.00123064f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_46 N_C2_M6_g N_C1_M7_g 0.0036939f $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_47 N_C2_c_67_n N_C1_c_78_n 9.33263e-19 $X=0.405 $Y=0.135 $X2=0.297 $Y2=0.135
cc_48 N_C2_c_68_n N_C1_c_79_n 0.00477924f $X=0.405 $Y=0.135 $X2=0.297 $Y2=0.135
cc_49 VSS N_C2_M6_g 3.57119e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_50 VSS N_C2_c_68_n 5.37372e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_51 N_C2_M6_g N_Y_c_97_n 2.56935e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_52 N_C2_c_68_n N_Y_c_97_n 0.00123064f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_53 VSS N_C1_M7_g 2.15135e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_54 N_C1_c_79_n N_Y_c_99_n 0.0013399f $X=0.459 $Y=0.135 $X2=0.349 $Y2=0.155
cc_55 N_C1_M7_g N_Y_c_100_n 2.64276e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_56 N_C1_c_79_n N_Y_c_100_n 0.00124805f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_57 N_C1_M7_g N_Y_c_102_n 2.76185e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_C1_c_79_n N_Y_c_102_n 0.0012322f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_59 N_C1_c_79_n N_Y_c_104_n 0.00391301f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_60 VSS N_Y_c_87_n 0.00138157f $X=0.216 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_61 VSS N_Y_c_88_n 2.88662e-19 $X=0.2085 $Y=0.072 $X2=0 $Y2=0
cc_62 VSS N_Y_c_107_n 2.88662e-19 $X=0.254 $Y=0.072 $X2=0 $Y2=0
cc_63 VSS N_Y_c_108_n 2.88662e-19 $X=0.315 $Y=0.072 $X2=0 $Y2=0
cc_64 VSS N_Y_c_109_n 2.99055e-19 $X=0.324 $Y=0.072 $X2=0 $Y2=0
cc_65 VSS N_Y_c_110_n 0.00333582f $X=0.378 $Y=0.036 $X2=0.243 $Y2=0.135
cc_66 VSS N_Y_c_110_n 0.00371671f $X=0.486 $Y=0.036 $X2=0.243 $Y2=0.135
cc_67 VSS N_Y_c_110_n 0.00250965f $X=0.4515 $Y=0.036 $X2=0.243 $Y2=0.135
cc_68 VSS N_Y_c_99_n 0.00138157f $X=0.486 $Y=0.036 $X2=0.243 $Y2=0.154
cc_69 VSS N_Y_c_109_n 4.54465e-19 $X=0.378 $Y=0.036 $X2=0 $Y2=0
cc_70 VSS N_Y_c_109_n 0.00365373f $X=0.4515 $Y=0.036 $X2=0 $Y2=0
cc_71 VSS N_Y_c_102_n 0.00365373f $X=0.486 $Y=0.036 $X2=0 $Y2=0
cc_72 VSS N_Y_c_117_n 2.47657e-19 $X=0.484 $Y=0.0675 $X2=0 $Y2=0
cc_73 VSS N_Y_c_117_n 0.00260156f $X=0.486 $Y=0.036 $X2=0 $Y2=0
cc_74 VSS N_Y_c_119_n 3.97918e-19 $X=0.486 $Y=0.036 $X2=0 $Y2=0
cc_75 VSS N_Y_c_107_n 3.48201e-19 $X=0.288 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_76 VSS N_Y_c_108_n 3.30547e-19 $X=0.339 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_77 VSS N_Y_c_122_p 3.30547e-19 $X=0.45 $Y=0.234 $X2=0.135 $Y2=0.0675

* END of "./OAI332xp33_ASAP7_75t_L.pex.sp.OAI332XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI333xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:58:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI333xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI333xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI333xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:58:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI333XP33_ASAP7_75T_L%C3 2 5 7 10 14 VSS
c4 10 VSS 0.00613146f $X=0.081 $Y=0.135
c5 5 VSS 0.00238289f $X=0.081 $Y=0.135
c6 2 VSS 0.062704f $X=0.081 $Y=0.0675
r7 10 14 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.156
r8 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r9 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r10 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI333XP33_ASAP7_75T_L%C2 2 5 7 10 14 VSS
c11 14 VSS 0.00132043f $X=0.129 $Y=0.154
c12 10 VSS 4.26629e-19 $X=0.135 $Y=0.135
c13 5 VSS 0.00123757f $X=0.135 $Y=0.135
c14 2 VSS 0.0598541f $X=0.135 $Y=0.0675
r15 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.154
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI333XP33_ASAP7_75T_L%C1 2 5 7 10 14 VSS
c11 10 VSS 0.00101969f $X=0.189 $Y=0.135
c12 5 VSS 0.00121257f $X=0.189 $Y=0.135
c13 2 VSS 0.0608354f $X=0.189 $Y=0.0675
r14 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.155
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI333XP33_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.243 $Y=0.135
c14 5 VSS 0.00111336f $X=0.243 $Y=0.135
c15 2 VSS 0.0617786f $X=0.243 $Y=0.0675
r16 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.154
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI333XP33_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.297 $Y=0.135
c14 5 VSS 0.00112198f $X=0.297 $Y=0.135
c15 2 VSS 0.0616432f $X=0.297 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OAI333XP33_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c12 10 VSS 7.27237e-19 $X=0.351 $Y=0.135
c13 5 VSS 0.00111185f $X=0.351 $Y=0.135
c14 2 VSS 0.0615515f $X=0.351 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OAI333XP33_ASAP7_75T_L%A3 2 5 7 10 14 VSS
c12 10 VSS 7.27237e-19 $X=0.405 $Y=0.135
c13 5 VSS 0.00111774f $X=0.405 $Y=0.135
c14 2 VSS 0.0615416f $X=0.405 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OAI333XP33_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c12 10 VSS 4.78074e-19 $X=0.459 $Y=0.135
c13 5 VSS 0.00114557f $X=0.459 $Y=0.135
c14 2 VSS 0.0623815f $X=0.459 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OAI333XP33_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c9 10 VSS 4.90626e-19 $X=0.513 $Y=0.135
c10 5 VSS 0.00171614f $X=0.513 $Y=0.135
c11 2 VSS 0.0671256f $X=0.513 $Y=0.0675
r12 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.155
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OAI333XP33_ASAP7_75T_L%Y 1 2 5 6 9 11 12 15 16 19 29 30 31 32 33 35
+ 37 38 39 40 41 45 54 55 56 62 64 VSS
c38 66 VSS 5.10117e-19 $X=0.567 $Y=0.2125
c39 64 VSS 8.61055e-19 $X=0.567 $Y=0.1245
c40 63 VSS 0.00112176f $X=0.567 $Y=0.106
c41 62 VSS 0.00322429f $X=0.572 $Y=0.143
c42 60 VSS 6.07272e-19 $X=0.567 $Y=0.225
c43 58 VSS 4.0892e-19 $X=0.531 $Y=0.072
c44 57 VSS 3.28227e-19 $X=0.522 $Y=0.072
c45 56 VSS 1.7724e-19 $X=0.515 $Y=0.072
c46 55 VSS 4.2636e-19 $X=0.504 $Y=0.072
c47 54 VSS 8.46035e-21 $X=0.468 $Y=0.072
c48 53 VSS 3.93699e-19 $X=0.45 $Y=0.072
c49 45 VSS 3.25927e-19 $X=0.432 $Y=0.072
c50 43 VSS 0.00335467f $X=0.558 $Y=0.072
c51 42 VSS 8.36318e-19 $X=0.531 $Y=0.234
c52 41 VSS 0.00142296f $X=0.522 $Y=0.234
c53 40 VSS 0.00344621f $X=0.504 $Y=0.234
c54 39 VSS 0.00142296f $X=0.468 $Y=0.234
c55 38 VSS 0.00329285f $X=0.45 $Y=0.234
c56 37 VSS 0.00142296f $X=0.414 $Y=0.234
c57 36 VSS 0.00688205f $X=0.396 $Y=0.234
c58 35 VSS 0.00142296f $X=0.36 $Y=0.234
c59 34 VSS 2.83817e-19 $X=0.342 $Y=0.234
c60 33 VSS 0.00320869f $X=0.34 $Y=0.234
c61 32 VSS 0.00146362f $X=0.306 $Y=0.234
c62 31 VSS 0.00340162f $X=0.288 $Y=0.234
c63 30 VSS 0.00146362f $X=0.252 $Y=0.234
c64 29 VSS 0.0041898f $X=0.234 $Y=0.234
c65 21 VSS 0.00607902f $X=0.558 $Y=0.234
c66 19 VSS 0.00251001f $X=0.538 $Y=0.2025
c67 15 VSS 0.00220422f $X=0.216 $Y=0.2025
c68 11 VSS 5.61153e-19 $X=0.233 $Y=0.2025
c69 9 VSS 0.00113516f $X=0.538 $Y=0.0675
c70 5 VSS 0.0023085f $X=0.432 $Y=0.0675
c71 1 VSS 5.91014e-19 $X=0.449 $Y=0.0675
r72 65 66 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.2 $X2=0.567 $Y2=0.2125
r73 63 64 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.106 $X2=0.567 $Y2=0.1245
r74 62 65 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.143 $X2=0.567 $Y2=0.2
r75 62 64 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.143 $X2=0.567 $Y2=0.1245
r76 60 66 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.225 $X2=0.567 $Y2=0.2125
r77 59 63 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.567 $Y2=0.106
r78 57 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.072 $X2=0.531 $Y2=0.072
r79 56 57 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.515
+ $Y=0.072 $X2=0.522 $Y2=0.072
r80 55 56 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.072 $X2=0.515 $Y2=0.072
r81 54 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.072 $X2=0.504 $Y2=0.072
r82 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.072 $X2=0.468 $Y2=0.072
r83 51 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.072 $X2=0.531 $Y2=0.072
r84 45 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.072 $X2=0.45 $Y2=0.072
r85 43 59 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.072 $X2=0.567 $Y2=0.081
r86 43 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.072 $X2=0.54 $Y2=0.072
r87 41 42 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.234 $X2=0.531 $Y2=0.234
r88 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.522 $Y2=0.234
r89 39 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.504 $Y2=0.234
r90 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r91 37 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.45 $Y2=0.234
r92 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r93 35 36 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.396 $Y2=0.234
r94 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r95 33 34 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.34
+ $Y=0.234 $X2=0.342 $Y2=0.234
r96 32 33 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.34 $Y2=0.234
r97 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r98 30 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.288 $Y2=0.234
r99 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r100 27 42 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.531 $Y2=0.234
r101 23 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.234 $Y2=0.234
r102 21 60 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.234 $X2=0.567 $Y2=0.225
r103 21 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.54 $Y2=0.234
r104 19 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r105 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.538 $Y2=0.2025
r106 15 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r107 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r108 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r109 9 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.072 $X2=0.54
+ $Y2=0.072
r110 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.538 $Y2=0.0675
r111 5 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.072 $X2=0.432
+ $Y2=0.072
r112 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r113 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
.ends


* END of "./OAI333xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI333xp33_ASAP7_75t_L  VSS VDD C3 C2 C1 B1 B2 B3 A3 A2 A1 Y
* 
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* B3	B3
* B2	B2
* B1	B1
* C1	C1
* C2	C2
* C3	C3
M0 noxref_12 N_C3_M0_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_C2_M1_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_12 N_C1_M2_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_13 N_B1_M3_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_12 N_B2_M4_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_13 N_B3_M5_g noxref_12 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 N_Y_M6_d N_A3_M6_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_13 N_A2_M7_g N_Y_M7_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_Y_M8_d N_A1_M8_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 noxref_15 N_C3_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M10 noxref_16 N_C2_M10_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.125 $Y=0.162
M11 N_Y_M11_d N_C1_M11_g noxref_16 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.179 $Y=0.162
M12 noxref_17 N_B1_M12_g N_Y_M12_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M13 noxref_18 N_B2_M13_g noxref_17 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M14 VDD N_B3_M14_g noxref_18 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M15 noxref_19 N_A3_M15_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M16 noxref_20 N_A2_M16_g noxref_19 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M17 N_Y_M17_d N_A1_M17_g noxref_20 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
*
* 
* .include "OAI333xp33_ASAP7_75t_L.pex.sp.OAI333XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI333xp33_ASAP7_75t_L.pex.sp.OAI333XP33_ASAP7_75T_L.pxi"
* File: OAI333xp33_ASAP7_75t_L.pex.sp.OAI333XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:58:33 2017
* 
x_PM_OAI333XP33_ASAP7_75T_L%C3 N_C3_M0_g N_C3_c_2_p N_C3_M9_g N_C3_c_3_p C3 VSS
+ PM_OAI333XP33_ASAP7_75T_L%C3
x_PM_OAI333XP33_ASAP7_75T_L%C2 N_C2_M1_g N_C2_c_6_n N_C2_M10_g N_C2_c_7_n C2 VSS
+ PM_OAI333XP33_ASAP7_75T_L%C2
x_PM_OAI333XP33_ASAP7_75T_L%C1 N_C1_M2_g N_C1_c_18_n N_C1_M11_g N_C1_c_19_n C1
+ VSS PM_OAI333XP33_ASAP7_75T_L%C1
x_PM_OAI333XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_29_n N_B1_M12_g N_B1_c_30_n B1
+ VSS PM_OAI333XP33_ASAP7_75T_L%B1
x_PM_OAI333XP33_ASAP7_75T_L%B2 N_B2_M4_g N_B2_c_42_n N_B2_M13_g N_B2_c_43_n B2
+ VSS PM_OAI333XP33_ASAP7_75T_L%B2
x_PM_OAI333XP33_ASAP7_75T_L%B3 N_B3_M5_g N_B3_c_55_n N_B3_M14_g N_B3_c_56_n B3
+ VSS PM_OAI333XP33_ASAP7_75T_L%B3
x_PM_OAI333XP33_ASAP7_75T_L%A3 N_A3_M6_g N_A3_c_67_n N_A3_M15_g N_A3_c_68_n A3
+ VSS PM_OAI333XP33_ASAP7_75T_L%A3
x_PM_OAI333XP33_ASAP7_75T_L%A2 N_A2_M7_g N_A2_c_79_n N_A2_M16_g N_A2_c_80_n A2
+ VSS PM_OAI333XP33_ASAP7_75T_L%A2
x_PM_OAI333XP33_ASAP7_75T_L%A1 N_A1_M8_g N_A1_c_91_n N_A1_M17_g N_A1_c_92_n A1
+ VSS PM_OAI333XP33_ASAP7_75T_L%A1
x_PM_OAI333XP33_ASAP7_75T_L%Y N_Y_M7_s N_Y_M6_d N_Y_c_124_n N_Y_M8_d N_Y_c_127_n
+ N_Y_M12_s N_Y_M11_d N_Y_c_98_n N_Y_M17_d N_Y_c_114_n N_Y_c_99_n N_Y_c_102_n
+ N_Y_c_121_n N_Y_c_104_n N_Y_c_122_n N_Y_c_106_n N_Y_c_108_n N_Y_c_134_p
+ N_Y_c_110_n N_Y_c_135_p N_Y_c_115_n N_Y_c_123_n N_Y_c_112_n N_Y_c_131_n
+ N_Y_c_117_n Y N_Y_c_118_n VSS PM_OAI333XP33_ASAP7_75T_L%Y
cc_1 N_C3_M0_g N_C2_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_C3_c_2_p N_C2_c_6_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_C3_c_3_p N_C2_c_7_n 0.00653171f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_C3_M0_g N_C1_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 N_C2_M1_g N_C1_M2_g 0.00327995f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_6 N_C2_c_6_n N_C1_c_18_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_7 N_C2_c_7_n N_C1_c_19_n 0.00466039f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_8 N_C2_M1_g N_B1_M3_g 2.71887e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_9 VSS N_C2_M1_g 3.62029e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_10 VSS N_C2_c_7_n 0.0012376f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_11 C2 N_Y_c_98_n 5.87506e-19 $X=0.129 $Y=0.154 $X2=0 $Y2=0
cc_12 C2 N_Y_c_99_n 4.59979e-19 $X=0.129 $Y=0.154 $X2=0 $Y2=0
cc_13 N_C1_M2_g N_B1_M3_g 0.0036939f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_C1_c_18_n N_B1_c_29_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 N_C1_c_19_n N_B1_c_30_n 0.00406615f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_16 N_C1_M2_g N_B2_M4_g 3.06651e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 VSS N_C1_M2_g 3.62029e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_18 VSS N_C1_c_19_n 0.0012322f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_19 N_C1_c_19_n N_Y_c_98_n 0.0013295f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_20 N_B1_M3_g N_B2_M4_g 0.00371573f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_21 N_B1_c_29_n N_B2_c_42_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_22 N_B1_c_30_n N_B2_c_43_n 0.00483372f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_23 N_B1_M3_g N_B3_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_24 VSS N_B1_M3_g 3.62029e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_25 VSS N_B1_c_30_n 0.0012322f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_26 N_B1_c_30_n N_Y_c_98_n 0.0013295f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_27 N_B1_M3_g N_Y_c_102_n 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_28 N_B1_c_30_n N_Y_c_102_n 0.00124805f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_29 N_B2_M4_g N_B3_M5_g 0.0036939f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_30 N_B2_c_42_n N_B3_c_55_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_31 N_B2_c_43_n N_B3_c_56_n 0.00483372f $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_32 N_B2_M4_g N_A3_M6_g 2.71887e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_33 VSS N_B2_M4_g 2.68514e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_34 VSS N_B2_c_43_n 0.00121543f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_35 VSS N_B2_M4_g 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B2_M4_g N_Y_c_104_n 3.48613e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_B2_c_43_n N_Y_c_104_n 0.00124805f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_38 N_B3_M5_g N_A3_M6_g 0.00333077f $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_39 N_B3_c_55_n N_A3_c_67_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_40 N_B3_c_56_n N_A3_c_68_n 0.00406615f $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_41 N_B3_M5_g N_A2_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_42 VSS N_B3_M5_g 3.47199e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_43 VSS N_B3_c_56_n 5.30079e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_44 N_B3_M5_g N_Y_c_106_n 2.56935e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_45 N_B3_c_56_n N_Y_c_106_n 0.00123064f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_46 N_A3_M6_g N_A2_M7_g 0.0036939f $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_47 N_A3_c_67_n N_A2_c_79_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.297 $Y2=0.135
cc_48 N_A3_c_68_n N_A2_c_80_n 0.00483372f $X=0.405 $Y=0.135 $X2=0.297 $Y2=0.135
cc_49 N_A3_M6_g N_A1_M8_g 3.06651e-19 $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_50 VSS N_A3_M6_g 3.37279e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_51 VSS N_A3_c_68_n 5.22785e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_52 N_A3_M6_g N_Y_c_108_n 2.45924e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_53 N_A3_c_68_n N_Y_c_108_n 0.00123064f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_54 N_A2_M7_g N_A1_M8_g 0.00376655f $X=0.459 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_55 N_A2_c_79_n N_A1_c_91_n 9.33263e-19 $X=0.459 $Y=0.135 $X2=0.351 $Y2=0.135
cc_56 N_A2_c_80_n N_A1_c_92_n 0.0048308f $X=0.459 $Y=0.135 $X2=0.351 $Y2=0.135
cc_57 VSS N_A2_M7_g 2.38303e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_A2_M7_g N_Y_c_110_n 3.38929e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_59 N_A2_c_80_n N_Y_c_110_n 0.00123064f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_60 N_A2_M7_g N_Y_c_112_n 2.76185e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_61 N_A2_c_80_n N_Y_c_112_n 0.0012322f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_62 N_A1_c_92_n N_Y_c_114_n 0.0013295f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_63 N_A1_M8_g N_Y_c_115_n 2.56935e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_A1_c_92_n N_Y_c_115_n 0.00123064f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_65 N_A1_c_92_n N_Y_c_117_n 0.00121543f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_66 N_A1_c_92_n N_Y_c_118_n 0.00391301f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_67 VSS N_Y_c_98_n 0.00138157f $X=0.216 $Y=0.0675 $X2=0 $Y2=0
cc_68 VSS N_Y_c_99_n 2.9391e-19 $X=0.2085 $Y=0.072 $X2=0 $Y2=0
cc_69 VSS N_Y_c_121_n 2.9391e-19 $X=0.254 $Y=0.072 $X2=0 $Y2=0
cc_70 VSS N_Y_c_122_n 2.9391e-19 $X=0.315 $Y=0.072 $X2=0 $Y2=0
cc_71 VSS N_Y_c_123_n 3.22079e-19 $X=0.324 $Y=0.072 $X2=0 $Y2=0
cc_72 VSS N_Y_c_124_n 0.003332f $X=0.378 $Y=0.036 $X2=0.243 $Y2=0.135
cc_73 VSS N_Y_c_124_n 0.00250965f $X=0.486 $Y=0.036 $X2=0.243 $Y2=0.135
cc_74 VSS N_Y_c_124_n 0.00355403f $X=0.486 $Y=0.036 $X2=0.243 $Y2=0.135
cc_75 VSS N_Y_c_127_n 3.14809e-19 $X=0.486 $Y=0.036 $X2=0.243 $Y2=0.135
cc_76 VSS N_Y_c_127_n 0.00337424f $X=0.486 $Y=0.036 $X2=0.243 $Y2=0.135
cc_77 VSS N_Y_c_123_n 4.6373e-19 $X=0.378 $Y=0.036 $X2=0 $Y2=0
cc_78 VSS N_Y_c_123_n 0.00881219f $X=0.486 $Y=0.036 $X2=0 $Y2=0
cc_79 VSS N_Y_c_131_n 0.00233206f $X=0.486 $Y=0.036 $X2=0 $Y2=0
cc_80 VSS N_Y_c_121_n 3.48201e-19 $X=0.288 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_81 VSS N_Y_c_122_n 3.4467e-19 $X=0.34 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_82 VSS N_Y_c_134_p 3.48201e-19 $X=0.45 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_83 VSS N_Y_c_135_p 3.48201e-19 $X=0.504 $Y=0.234 $X2=0.135 $Y2=0.0675

* END of "./OAI333xp33_ASAP7_75t_L.pex.sp.OAI333XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: OAI33xp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:58:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OAI33xp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./OAI33xp33_ASAP7_75t_L.pex.sp.pex"
* File: OAI33xp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:58:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OAI33XP33_ASAP7_75T_L%A3 2 5 7 11 15 VSS
c10 15 VSS 0.00163529f $X=0.081 $Y=0.155
c11 11 VSS 8.01854e-19 $X=0.081 $Y=0.135
c12 5 VSS 0.00168113f $X=0.081 $Y=0.135
c13 2 VSS 0.0658433f $X=0.081 $Y=0.0675
r14 11 15 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.155
r15 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OAI33XP33_ASAP7_75T_L%A2 2 5 7 10 14 VSS
c12 10 VSS 4.78074e-19 $X=0.135 $Y=0.135
c13 5 VSS 0.00114323f $X=0.135 $Y=0.135
c14 2 VSS 0.0623258f $X=0.135 $Y=0.0675
r15 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.155
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OAI33XP33_ASAP7_75T_L%A1 2 5 7 10 14 VSS
c14 10 VSS 4.81053e-19 $X=0.189 $Y=0.135
c15 5 VSS 0.00112856f $X=0.189 $Y=0.135
c16 2 VSS 0.0624435f $X=0.189 $Y=0.0675
r17 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.155
r18 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r19 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r20 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OAI33XP33_ASAP7_75T_L%B1 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.243 $Y=0.135
c14 5 VSS 0.00112856f $X=0.243 $Y=0.135
c15 2 VSS 0.0627054f $X=0.243 $Y=0.0675
r16 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.154
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OAI33XP33_ASAP7_75T_L%B2 2 5 7 10 14 VSS
c13 10 VSS 4.81053e-19 $X=0.297 $Y=0.135
c14 5 VSS 0.00112198f $X=0.297 $Y=0.135
c15 2 VSS 0.0616432f $X=0.297 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OAI33XP33_ASAP7_75T_L%B3 2 5 7 10 14 VSS
c13 10 VSS 7.13761e-19 $X=0.351 $Y=0.135
c14 5 VSS 0.00111707f $X=0.351 $Y=0.135
c15 2 VSS 0.0611572f $X=0.351 $Y=0.0675
r16 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.155
r17 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OAI33XP33_ASAP7_75T_L%C3 2 5 7 10 16 VSS
c14 10 VSS 0.00175162f $X=0.405 $Y=0.135
c15 5 VSS 0.00110628f $X=0.405 $Y=0.135
c16 2 VSS 0.059756f $X=0.405 $Y=0.0675
r17 10 16 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.156
r18 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r19 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r20 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_OAI33XP33_ASAP7_75T_L%C2 2 5 7 10 14 VSS
c12 10 VSS 0.00154575f $X=0.459 $Y=0.135
c13 5 VSS 0.00113128f $X=0.459 $Y=0.135
c14 2 VSS 0.0597446f $X=0.459 $Y=0.0675
r15 10 14 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.154
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_OAI33XP33_ASAP7_75T_L%C1 2 5 7 10 14 VSS
c10 10 VSS 0.00299346f $X=0.513 $Y=0.135
c11 5 VSS 0.00222969f $X=0.513 $Y=0.135
c12 2 VSS 0.0636632f $X=0.513 $Y=0.0675
r13 10 14 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.155
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_OAI33XP33_ASAP7_75T_L%Y 1 6 7 11 12 15 16 19 24 26 28 30 34 38 39 48
+ 49 50 51 52 56 57 58 59 60 61 62 63 64 65 66 67 VSS
c50 67 VSS 0.00146362f $X=0.522 $Y=0.234
c51 66 VSS 0.00347187f $X=0.504 $Y=0.234
c52 65 VSS 0.00146362f $X=0.468 $Y=0.234
c53 64 VSS 0.00356553f $X=0.45 $Y=0.234
c54 63 VSS 0.00146362f $X=0.414 $Y=0.234
c55 62 VSS 0.0067709f $X=0.396 $Y=0.234
c56 61 VSS 0.00146362f $X=0.36 $Y=0.234
c57 60 VSS 0.00340842f $X=0.342 $Y=0.234
c58 59 VSS 0.00146362f $X=0.306 $Y=0.234
c59 58 VSS 0.00340842f $X=0.288 $Y=0.234
c60 57 VSS 0.00146362f $X=0.252 $Y=0.234
c61 56 VSS 0.00347104f $X=0.234 $Y=0.234
c62 54 VSS 0.00690733f $X=0.54 $Y=0.234
c63 52 VSS 0.00146362f $X=0.198 $Y=0.234
c64 51 VSS 0.00325506f $X=0.18 $Y=0.234
c65 50 VSS 0.00146362f $X=0.144 $Y=0.234
c66 49 VSS 0.00340842f $X=0.126 $Y=0.234
c67 48 VSS 0.00470799f $X=0.09 $Y=0.234
c68 47 VSS 0.00451896f $X=0.053 $Y=0.234
c69 43 VSS 0.00328056f $X=0.027 $Y=0.234
c70 41 VSS 6.55192e-19 $X=0.077 $Y=0.036
c71 40 VSS 0.00192646f $X=0.072 $Y=0.036
c72 39 VSS 0.00238885f $X=0.162 $Y=0.036
c73 38 VSS 0.00914531f $X=0.162 $Y=0.036
c74 35 VSS 0.00303439f $X=0.053 $Y=0.036
c75 34 VSS 0.00345727f $X=0.054 $Y=0.036
c76 31 VSS 0.00322101f $X=0.027 $Y=0.036
c77 30 VSS 7.47379e-19 $X=0.018 $Y=0.207
c78 28 VSS 9.68e-19 $X=0.018 $Y=0.1245
c79 27 VSS 9.60196e-19 $X=0.018 $Y=0.106
c80 26 VSS 7.3752e-19 $X=0.018 $Y=0.081
c81 25 VSS 8.29409e-19 $X=0.018 $Y=0.063
c82 24 VSS 0.00294659f $X=0.018 $Y=0.143
c83 22 VSS 8.29409e-19 $X=0.018 $Y=0.225
c84 19 VSS 0.00358415f $X=0.538 $Y=0.2025
c85 15 VSS 0.00233324f $X=0.216 $Y=0.2025
c86 11 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c87 6 VSS 6.29123e-19 $X=0.179 $Y=0.0675
c88 1 VSS 2.69461e-19 $X=0.071 $Y=0.0675
r89 66 67 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.522 $Y2=0.234
r90 65 66 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.504 $Y2=0.234
r91 64 65 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r92 63 64 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.45 $Y2=0.234
r93 62 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r94 61 62 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.234 $X2=0.396 $Y2=0.234
r95 60 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.36 $Y2=0.234
r96 59 60 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.342 $Y2=0.234
r97 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r98 57 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.288 $Y2=0.234
r99 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r100 54 67 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.522 $Y2=0.234
r101 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r102 50 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.18 $Y2=0.234
r103 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r104 48 49 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.126 $Y2=0.234
r105 47 48 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.053
+ $Y=0.234 $X2=0.09 $Y2=0.234
r106 45 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.234 $Y2=0.234
r107 45 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.198 $Y2=0.234
r108 43 47 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.053 $Y2=0.234
r109 40 41 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.077 $Y2=0.036
r110 38 41 5.77161 $w=1.8e-08 $l=8.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.077 $Y2=0.036
r111 38 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r112 35 36 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.053
+ $Y=0.036 $X2=0.0535 $Y2=0.036
r113 33 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.072 $Y2=0.036
r114 33 36 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0535 $Y2=0.036
r115 33 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r116 31 35 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.053 $Y2=0.036
r117 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.207
r118 27 28 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.106 $X2=0.018 $Y2=0.1245
r119 26 27 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.106
r120 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.081
r121 24 29 3.12346 $w=1.8e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.143 $X2=0.018 $Y2=0.189
r122 24 28 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.143 $X2=0.018 $Y2=0.1245
r123 22 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r124 22 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.207
r125 21 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r126 21 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r127 19 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r128 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.538 $Y2=0.2025
r129 15 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r130 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r131 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r132 10 39 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.162 $Y=0.0675 $X2=0.162 $Y2=0.036
r133 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r134 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r135 4 34 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r136 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./OAI33xp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt OAI33xp33_ASAP7_75t_L  VSS VDD A3 A2 A1 B1 B2 B3 C3 C2 C1 Y
* 
* Y	Y
* C1	C1
* C2	C2
* C3	C3
* B3	B3
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
M0 noxref_13 N_A3_M0_g N_Y_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_Y_M1_d N_A2_M1_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 noxref_13 N_A1_M2_g N_Y_M2_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 noxref_14 N_B1_M3_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 noxref_13 N_B2_M4_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 noxref_14 N_B3_M5_g noxref_13 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 VSS N_C3_M6_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 noxref_14 N_C2_M7_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 VSS N_C1_M8_g noxref_14 VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 noxref_15 N_A3_M9_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M10 noxref_16 N_A2_M10_g noxref_15 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.125 $Y=0.162
M11 N_Y_M11_d N_A1_M11_g noxref_16 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.179 $Y=0.162
M12 noxref_17 N_B1_M12_g N_Y_M12_s VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M13 noxref_18 N_B2_M13_g noxref_17 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M14 VDD N_B3_M14_g noxref_18 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M15 noxref_19 N_C3_M15_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M16 noxref_20 N_C2_M16_g noxref_19 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M17 N_Y_M17_d N_C1_M17_g noxref_20 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
*
* 
* .include "OAI33xp33_ASAP7_75t_L.pex.sp.OAI33XP33_ASAP7_75T_L.pxi"
* BEGIN of "./OAI33xp33_ASAP7_75t_L.pex.sp.OAI33XP33_ASAP7_75T_L.pxi"
* File: OAI33xp33_ASAP7_75t_L.pex.sp.OAI33XP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:58:56 2017
* 
x_PM_OAI33XP33_ASAP7_75T_L%A3 N_A3_M0_g N_A3_c_2_p N_A3_M9_g N_A3_c_3_p A3 VSS
+ PM_OAI33XP33_ASAP7_75T_L%A3
x_PM_OAI33XP33_ASAP7_75T_L%A2 N_A2_M1_g N_A2_c_12_n N_A2_M10_g N_A2_c_13_n A2
+ VSS PM_OAI33XP33_ASAP7_75T_L%A2
x_PM_OAI33XP33_ASAP7_75T_L%A1 N_A1_M2_g N_A1_c_25_n N_A1_M11_g N_A1_c_26_n A1
+ VSS PM_OAI33XP33_ASAP7_75T_L%A1
x_PM_OAI33XP33_ASAP7_75T_L%B1 N_B1_M3_g N_B1_c_39_n N_B1_M12_g N_B1_c_40_n B1
+ VSS PM_OAI33XP33_ASAP7_75T_L%B1
x_PM_OAI33XP33_ASAP7_75T_L%B2 N_B2_M4_g N_B2_c_52_n N_B2_M13_g N_B2_c_53_n B2
+ VSS PM_OAI33XP33_ASAP7_75T_L%B2
x_PM_OAI33XP33_ASAP7_75T_L%B3 N_B3_M5_g N_B3_c_65_n N_B3_M14_g N_B3_c_66_n B3
+ VSS PM_OAI33XP33_ASAP7_75T_L%B3
x_PM_OAI33XP33_ASAP7_75T_L%C3 N_C3_M6_g N_C3_c_78_n N_C3_M15_g N_C3_c_79_n C3
+ VSS PM_OAI33XP33_ASAP7_75T_L%C3
x_PM_OAI33XP33_ASAP7_75T_L%C2 N_C2_M7_g N_C2_c_92_n N_C2_M16_g N_C2_c_93_n C2
+ VSS PM_OAI33XP33_ASAP7_75T_L%C2
x_PM_OAI33XP33_ASAP7_75T_L%C1 N_C1_M8_g N_C1_c_104_n N_C1_M17_g N_C1_c_105_n C1
+ VSS PM_OAI33XP33_ASAP7_75T_L%C1
x_PM_OAI33XP33_ASAP7_75T_L%Y N_Y_M0_s N_Y_M2_s N_Y_M1_d N_Y_M12_s N_Y_M11_d
+ N_Y_c_119_n N_Y_M17_d N_Y_c_134_n Y N_Y_c_143_p N_Y_c_112_n N_Y_c_113_n
+ N_Y_c_137_p N_Y_c_116_n N_Y_c_139_p N_Y_c_114_n N_Y_c_146_p N_Y_c_117_n
+ N_Y_c_147_p N_Y_c_121_n N_Y_c_149_p N_Y_c_124_n N_Y_c_150_p N_Y_c_126_n
+ N_Y_c_151_p N_Y_c_128_n N_Y_c_154_p N_Y_c_130_n N_Y_c_155_p N_Y_c_132_n
+ N_Y_c_153_p N_Y_c_135_n VSS PM_OAI33XP33_ASAP7_75T_L%Y
cc_1 N_A3_M0_g N_A2_M1_g 0.0036939f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A3_c_2_p N_A2_c_12_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A3_c_3_p N_A2_c_13_n 0.00473719f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A3_M0_g N_A1_M2_g 3.06651e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 N_A3_c_3_p N_Y_c_112_n 0.0026314f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_6 A3 N_Y_c_113_n 9.68179e-19 $X=0.081 $Y=0.155 $X2=0 $Y2=0
cc_7 N_A3_M0_g N_Y_c_114_n 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_8 A3 N_Y_c_114_n 0.00380759f $X=0.081 $Y=0.155 $X2=0 $Y2=0
cc_9 VSS N_A3_M0_g 3.32429e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_10 VSS N_A3_c_3_p 0.00112429f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 N_A2_M1_g N_A1_M2_g 0.00376655f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_12 N_A2_c_12_n N_A1_c_25_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_13 N_A2_c_13_n N_A1_c_26_n 0.00483372f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 N_A2_M1_g N_B1_M3_g 3.12393e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_15 N_A2_M1_g N_Y_c_116_n 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_16 N_A2_M1_g N_Y_c_117_n 3.48613e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_17 N_A2_c_13_n N_Y_c_117_n 0.00124805f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_18 VSS N_A2_M1_g 2.76185e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 VSS N_A2_c_13_n 0.0012322f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_20 N_A1_M2_g N_B1_M3_g 0.00381737f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_21 N_A1_c_25_n N_B1_c_39_n 8.86777e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 N_A1_c_26_n N_B1_c_40_n 0.00406615f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 N_A1_M2_g N_B2_M4_g 3.12393e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_24 N_A1_c_26_n N_Y_c_119_n 0.0013295f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.155
cc_25 N_A1_M2_g N_Y_c_116_n 2.04849e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_A1_M2_g N_Y_c_121_n 2.56935e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_A1_c_26_n N_Y_c_121_n 0.00124805f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_28 VSS N_A1_c_26_n 0.00120704f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_29 VSS N_A1_M2_g 2.86606e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_B1_M3_g N_B2_M4_g 0.00376655f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_31 N_B1_c_39_n N_B2_c_52_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_32 N_B1_c_40_n N_B2_c_53_n 0.00483372f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_33 N_B1_M3_g N_B3_M5_g 3.06651e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_34 N_B1_c_40_n N_Y_c_119_n 0.0013295f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_35 N_B1_M3_g N_Y_c_124_n 2.64276e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B1_c_40_n N_Y_c_124_n 0.00124805f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_37 VSS N_B1_c_40_n 0.00121543f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_38 VSS N_B1_M3_g 2.81289e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_B2_M4_g N_B3_M5_g 0.00364308f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_40 N_B2_c_52_n N_B3_c_65_n 8.86777e-19 $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_41 N_B2_c_53_n N_B3_c_66_n 0.00483372f $X=0.297 $Y=0.135 $X2=0.189 $Y2=0.135
cc_42 N_B2_M4_g N_C3_M6_g 2.66145e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_43 N_B2_M4_g N_Y_c_126_n 3.48613e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_B2_c_53_n N_Y_c_126_n 0.00124805f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_45 VSS N_B2_M4_g 2.68514e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_46 VSS N_B2_c_53_n 0.00121543f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_47 VSS N_B2_M4_g 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_48 N_B3_M5_g N_C3_M6_g 0.0032073f $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_49 N_B3_c_65_n N_C3_c_78_n 8.86777e-19 $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_50 N_B3_c_66_n N_C3_c_79_n 0.00389755f $X=0.351 $Y=0.135 $X2=0.243 $Y2=0.135
cc_51 N_B3_M5_g N_C2_M7_g 2.31381e-19 $X=0.351 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_52 N_B3_M5_g N_Y_c_128_n 2.64276e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_53 N_B3_c_66_n N_Y_c_128_n 0.00124805f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_54 VSS N_B3_M5_g 2.34106e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_55 VSS N_B3_c_66_n 7.19406e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_56 VSS N_B3_c_66_n 2.9854e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_57 N_C3_M6_g N_C2_M7_g 0.0032073f $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_58 N_C3_c_78_n N_C2_c_92_n 8.86777e-19 $X=0.405 $Y=0.135 $X2=0.297 $Y2=0.135
cc_59 N_C3_c_79_n N_C2_c_93_n 0.00581998f $X=0.405 $Y=0.135 $X2=0.297 $Y2=0.135
cc_60 N_C3_M6_g N_C1_M8_g 2.66145e-19 $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_61 N_C3_M6_g N_Y_c_130_n 2.64276e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_62 N_C3_c_79_n N_Y_c_130_n 0.00125352f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_63 VSS N_C3_c_79_n 3.41423e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_64 VSS N_C3_c_79_n 8.59553e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_65 VSS N_C3_M6_g 2.64276e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_66 VSS N_C3_c_79_n 0.00125352f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_67 N_C2_M7_g N_C1_M8_g 0.0035196f $X=0.459 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_68 N_C2_c_92_n N_C1_c_104_n 9.33263e-19 $X=0.459 $Y=0.135 $X2=0.351 $Y2=0.135
cc_69 N_C2_c_93_n N_C1_c_105_n 0.00582751f $X=0.459 $Y=0.135 $X2=0.351 $Y2=0.135
cc_70 N_C2_M7_g N_Y_c_132_n 3.48613e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_71 N_C2_c_93_n N_Y_c_132_n 0.00125352f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_72 VSS N_C2_c_93_n 0.00114532f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_73 VSS N_C2_M7_g 2.64276e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_74 VSS N_C2_c_93_n 0.00125352f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_75 N_C1_c_105_n N_Y_c_134_n 0.00165292f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_76 N_C1_M8_g N_Y_c_135_n 2.64276e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_77 N_C1_c_105_n N_Y_c_135_n 0.00125352f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_78 VSS N_C1_M8_g 2.1563e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_79 VSS N_C1_c_105_n 0.00101217f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_80 VSS N_C1_c_105_n 0.00114532f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_81 VSS N_Y_c_137_p 0.00336248f $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.135
cc_82 VSS N_Y_c_116_n 0.00250965f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_83 VSS N_Y_c_139_p 0.00355401f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_84 VSS N_Y_c_119_n 0.00138157f $X=0.216 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_85 VSS N_Y_c_116_n 4.51937e-19 $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_86 VSS N_Y_c_139_p 0.00322522f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_87 VSS N_Y_c_143_p 3.9223e-19 $X=0.018 $Y=0.081 $X2=0 $Y2=0
cc_88 VSS N_Y_c_137_p 5.38872e-19 $X=0.054 $Y=0.036 $X2=0 $Y2=0
cc_89 VSS N_Y_c_116_n 0.00906393f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_90 VSS N_Y_c_146_p 3.20199e-19 $X=0.126 $Y=0.234 $X2=0 $Y2=0
cc_91 VSS N_Y_c_147_p 3.20199e-19 $X=0.18 $Y=0.234 $X2=0 $Y2=0
cc_92 VSS N_Y_c_139_p 0.00233206f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_93 VSS N_Y_c_149_p 3.20199e-19 $X=0.234 $Y=0.234 $X2=0 $Y2=0
cc_94 VSS N_Y_c_150_p 3.20199e-19 $X=0.288 $Y=0.234 $X2=0 $Y2=0
cc_95 VSS N_Y_c_151_p 3.20199e-19 $X=0.342 $Y=0.234 $X2=0 $Y2=0
cc_96 VSS N_Y_c_116_n 3.9033e-19 $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_97 VSS N_Y_c_153_p 2.18766e-19 $X=0.504 $Y=0.234 $X2=0 $Y2=0
cc_98 VSS N_Y_c_154_p 2.18766e-19 $X=0.396 $Y=0.234 $X2=0 $Y2=0
cc_99 VSS N_Y_c_155_p 2.18766e-19 $X=0.45 $Y=0.234 $X2=0 $Y2=0
cc_100 VSS N_Y_c_146_p 3.62324e-19 $X=0.126 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_101 VSS N_Y_c_147_p 3.62324e-19 $X=0.18 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_102 VSS N_Y_c_150_p 3.62324e-19 $X=0.288 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_103 VSS N_Y_c_151_p 3.62324e-19 $X=0.342 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_104 VSS N_Y_c_155_p 3.71563e-19 $X=0.45 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_105 VSS N_Y_c_153_p 3.71563e-19 $X=0.504 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./OAI33xp33_ASAP7_75t_L.pex.sp.OAI33XP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: O2A1O1Ixp33_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:46:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "O2A1O1Ixp33_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./O2A1O1Ixp33_ASAP7_75t_L.pex.sp.pex"
* File: O2A1O1Ixp33_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:46:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_O2A1O1IXP33_ASAP7_75T_L%A2 2 5 7 13 VSS
c9 13 VSS 0.0010791f $X=0.082 $Y=0.138
c10 5 VSS 0.00220625f $X=0.081 $Y=0.135
c11 2 VSS 0.0633348f $X=0.081 $Y=0.0675
r12 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_O2A1O1IXP33_ASAP7_75T_L%A1 2 5 7 13 VSS
c12 13 VSS 0.00164686f $X=0.136 $Y=0.138
c13 5 VSS 0.00114698f $X=0.135 $Y=0.135
c14 2 VSS 0.0587206f $X=0.135 $Y=0.0675
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_O2A1O1IXP33_ASAP7_75T_L%B 2 5 7 13 VSS
c12 13 VSS 0.00167842f $X=0.191 $Y=0.136
c13 5 VSS 0.00113686f $X=0.189 $Y=0.135
c14 2 VSS 0.0582057f $X=0.189 $Y=0.0675
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_O2A1O1IXP33_ASAP7_75T_L%C 2 5 7 15 VSS
c11 15 VSS 0.00221489f $X=0.242 $Y=0.136
c12 5 VSS 0.00178699f $X=0.243 $Y=0.135
c13 2 VSS 0.0626166f $X=0.243 $Y=0.054
r14 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r16 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_O2A1O1IXP33_ASAP7_75T_L%7 1 4 6 7 10 16 18 19 20 21 22 23 VSS
c15 23 VSS 1.34897e-19 $X=0.153 $Y=0.072
c16 22 VSS 8.46035e-21 $X=0.144 $Y=0.072
c17 21 VSS 3.38991e-19 $X=0.126 $Y=0.072
c18 20 VSS 2.03419e-19 $X=0.094 $Y=0.072
c19 19 VSS 5.31938e-19 $X=0.09 $Y=0.072
c20 18 VSS 0.002538f $X=0.072 $Y=0.072
c21 16 VSS 0.00100696f $X=0.162 $Y=0.072
c22 10 VSS 0.00757825f $X=0.162 $Y=0.0675
c23 6 VSS 5.76042e-19 $X=0.179 $Y=0.0675
c24 4 VSS 8.25856e-19 $X=0.056 $Y=0.0675
c25 1 VSS 3.34937e-19 $X=0.071 $Y=0.0675
r26 22 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.153 $Y2=0.072
r27 21 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.144 $Y2=0.072
r28 20 21 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.072 $X2=0.126 $Y2=0.072
r29 19 20 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.094 $Y2=0.072
r30 18 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.072 $X2=0.09 $Y2=0.072
r31 16 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.072 $X2=0.153 $Y2=0.072
r32 12 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.072 $X2=0.072 $Y2=0.072
r33 10 16 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.072 $X2=0.162
+ $Y2=0.072
r34 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r35 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r36 4 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.072 $X2=0.054
+ $Y2=0.072
r37 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends

.subckt PM_O2A1O1IXP33_ASAP7_75T_L%Y 1 2 6 9 11 14 19 24 26 29 35 45 VSS
c16 45 VSS 0.00328191f $X=0.288 $Y=0.234
c17 44 VSS 0.00277971f $X=0.297 $Y=0.234
c18 39 VSS 3.14564e-19 $X=0.297 $Y=0.2155
c19 37 VSS 2.86471e-19 $X=0.297 $Y=0.07
c20 36 VSS 5.7946e-19 $X=0.297 $Y=0.063
c21 35 VSS 0.0059242f $X=0.298 $Y=0.136
c22 33 VSS 7.46764e-19 $X=0.297 $Y=0.225
c23 31 VSS 4.50206e-19 $X=0.2655 $Y=0.036
c24 30 VSS 8.40992e-19 $X=0.261 $Y=0.036
c25 29 VSS 0.00146362f $X=0.252 $Y=0.036
c26 28 VSS 0.00140647f $X=0.234 $Y=0.036
c27 27 VSS 0.00457115f $X=0.225 $Y=0.036
c28 26 VSS 0.00142296f $X=0.198 $Y=0.036
c29 25 VSS 4.81555e-19 $X=0.18 $Y=0.036
c30 24 VSS 0.00691396f $X=0.176 $Y=0.036
c31 19 VSS 0.00272524f $X=0.108 $Y=0.036
c32 16 VSS 0.00565494f $X=0.288 $Y=0.036
c33 14 VSS 0.0032709f $X=0.268 $Y=0.2025
c34 9 VSS 0.00592134f $X=0.268 $Y=0.054
c35 1 VSS 6.469e-19 $X=0.125 $Y=0.0675
r36 45 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.2925 $Y2=0.234
r37 44 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.234 $X2=0.2925 $Y2=0.234
r38 41 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.288 $Y2=0.234
r39 38 39 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.206 $X2=0.297 $Y2=0.2155
r40 36 37 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.063 $X2=0.297 $Y2=0.07
r41 35 38 4.75309 $w=1.8e-08 $l=7e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.136 $X2=0.297 $Y2=0.206
r42 35 37 4.48148 $w=1.8e-08 $l=6.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.136 $X2=0.297 $Y2=0.07
r43 33 44 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.234
r44 33 39 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.2155
r45 32 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.063
r46 30 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.036 $X2=0.2655 $Y2=0.036
r47 29 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.261 $Y2=0.036
r48 28 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r49 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.036 $X2=0.234 $Y2=0.036
r50 26 27 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.225 $Y2=0.036
r51 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r52 24 25 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.036 $X2=0.18 $Y2=0.036
r53 22 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.2655 $Y2=0.036
r54 18 24 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.176 $Y2=0.036
r55 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r56 16 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r57 16 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.27 $Y2=0.036
r58 14 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r59 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.268 $Y2=0.2025
r60 9 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r61 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.054 $X2=0.268 $Y2=0.054
r62 5 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r63 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r64 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./O2A1O1Ixp33_ASAP7_75t_L.pex.sp.pex"
* 
.subckt O2A1O1Ixp33_ASAP7_75t_L  VSS VDD A2 A1 B C Y
* 
* Y	Y
* C	C
* B	B
* A1	A1
* A2	A2
M0 N_Y_M0_d N_A2_M0_g N_7_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_7_M1_d N_A1_M1_g N_Y_M1_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_B_M2_g N_7_M2_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_C_M3_g VSS VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 noxref_10 N_A2_M4_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 VDD N_A1_M5_g noxref_10 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 noxref_8 N_B_M6_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M7 N_Y_M7_d N_C_M7_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
*
* 
* .include "O2A1O1Ixp33_ASAP7_75t_L.pex.sp.O2A1O1IXP33_ASAP7_75T_L.pxi"
* BEGIN of "./O2A1O1Ixp33_ASAP7_75t_L.pex.sp.O2A1O1IXP33_ASAP7_75T_L.pxi"
* File: O2A1O1Ixp33_ASAP7_75t_L.pex.sp.O2A1O1IXP33_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:46:34 2017
* 
x_PM_O2A1O1IXP33_ASAP7_75T_L%A2 N_A2_M0_g N_A2_c_2_p N_A2_M4_g A2 VSS
+ PM_O2A1O1IXP33_ASAP7_75T_L%A2
x_PM_O2A1O1IXP33_ASAP7_75T_L%A1 N_A1_M1_g N_A1_c_11_n N_A1_M5_g A1 VSS
+ PM_O2A1O1IXP33_ASAP7_75T_L%A1
x_PM_O2A1O1IXP33_ASAP7_75T_L%B N_B_M2_g N_B_c_24_n N_B_M6_g B VSS
+ PM_O2A1O1IXP33_ASAP7_75T_L%B
x_PM_O2A1O1IXP33_ASAP7_75T_L%C N_C_M3_g N_C_c_36_n N_C_M7_g C VSS
+ PM_O2A1O1IXP33_ASAP7_75T_L%C
x_PM_O2A1O1IXP33_ASAP7_75T_L%7 N_7_M0_s N_7_c_50_p N_7_M2_s N_7_M1_d N_7_c_55_p
+ N_7_c_49_n N_7_c_51_p N_7_c_45_n N_7_c_52_p N_7_c_56_p N_7_c_47_n N_7_c_53_p
+ VSS PM_O2A1O1IXP33_ASAP7_75T_L%7
x_PM_O2A1O1IXP33_ASAP7_75T_L%Y N_Y_M1_s N_Y_M0_d N_Y_M3_d N_Y_c_63_n N_Y_M7_d
+ N_Y_c_64_n N_Y_c_68_n N_Y_c_60_n N_Y_c_61_n N_Y_c_65_n Y N_Y_c_75_n VSS
+ PM_O2A1O1IXP33_ASAP7_75T_L%Y
cc_1 N_A2_M0_g N_A1_M1_g 0.00348334f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A2_c_2_p N_A1_c_11_n 9.33263e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A2 A1 0.00477924f $X=0.082 $Y=0.138 $X2=0.136 $Y2=0.138
cc_4 N_A2_M0_g N_B_M2_g 2.48122e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 N_A2_M0_g N_7_c_45_n 3.62029e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_6 A2 N_7_c_45_n 0.0012322f $X=0.082 $Y=0.138 $X2=0 $Y2=0
cc_7 VSS A2 8.92951e-19 $X=0.082 $Y=0.138 $X2=0.135 $Y2=0.135
cc_8 VSS N_A2_M0_g 2.64276e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_9 VSS A2 0.00124805f $X=0.082 $Y=0.138 $X2=0 $Y2=0
cc_10 N_A1_M1_g N_B_M2_g 0.00304756f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_11 N_A1_c_11_n N_B_c_24_n 8.86777e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_12 A1 B 0.00406615f $X=0.136 $Y=0.138 $X2=0.082 $Y2=0.138
cc_13 N_A1_M1_g N_C_M3_g 2.13359e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_A1_M1_g N_7_c_47_n 2.68514e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 A1 N_7_c_47_n 0.00121543f $X=0.136 $Y=0.138 $X2=0 $Y2=0
cc_16 VSS N_A1_M1_g 2.64276e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_17 VSS A1 0.00124805f $X=0.136 $Y=0.138 $X2=0 $Y2=0
cc_18 N_A1_M1_g N_Y_c_60_n 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 N_B_M2_g N_C_M3_g 0.00304756f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_20 N_B_c_24_n N_C_c_36_n 9.33263e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 B C 0.00382941f $X=0.191 $Y=0.136 $X2=0 $Y2=0
cc_22 VSS B 0.00114532f $X=0.191 $Y=0.136 $X2=0.081 $Y2=0.135
cc_23 VSS N_B_M2_g 2.56935e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 VSS B 0.00123064f $X=0.191 $Y=0.136 $X2=0 $Y2=0
cc_25 N_B_M2_g N_Y_c_61_n 3.47199e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 B N_Y_c_61_n 5.30079e-19 $X=0.191 $Y=0.136 $X2=0 $Y2=0
cc_27 C N_7_c_49_n 2.63981e-19 $X=0.242 $Y=0.136 $X2=0 $Y2=0
cc_28 VSS C 0.00124888f $X=0.242 $Y=0.136 $X2=0.135 $Y2=0.135
cc_29 C N_Y_c_63_n 3.24828e-19 $X=0.242 $Y=0.136 $X2=0 $Y2=0
cc_30 C N_Y_c_64_n 0.00131945f $X=0.242 $Y=0.136 $X2=0 $Y2=0
cc_31 N_C_M3_g N_Y_c_65_n 2.64276e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_32 C N_Y_c_65_n 0.00125417f $X=0.242 $Y=0.136 $X2=0 $Y2=0
cc_33 C Y 0.00559493f $X=0.242 $Y=0.136 $X2=0 $Y2=0
cc_34 VSS N_7_c_50_p 0.00138157f $X=0.056 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_35 VSS N_7_c_51_p 2.62991e-19 $X=0.072 $Y=0.072 $X2=0 $Y2=0
cc_36 VSS N_7_c_52_p 2.62991e-19 $X=0.094 $Y=0.072 $X2=0 $Y2=0
cc_37 VSS N_7_c_53_p 2.62991e-19 $X=0.153 $Y=0.072 $X2=0 $Y2=0
cc_38 N_7_c_50_p N_Y_c_68_n 0.00328221f $X=0.056 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_7_c_55_p N_Y_c_68_n 0.00355395f $X=0.162 $Y=0.0675 $X2=0 $Y2=0
cc_40 N_7_c_56_p N_Y_c_68_n 0.00233206f $X=0.126 $Y=0.072 $X2=0 $Y2=0
cc_41 N_7_c_50_p N_Y_c_60_n 3.09693e-19 $X=0.056 $Y=0.0675 $X2=0 $Y2=0
cc_42 N_7_c_55_p N_Y_c_60_n 0.00250962f $X=0.162 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_7_c_56_p N_Y_c_60_n 0.00675381f $X=0.126 $Y=0.072 $X2=0 $Y2=0
cc_44 VSS N_Y_c_64_n 0.00389029f $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_45 VSS N_Y_c_75_n 6.56506e-19 $X=0.216 $Y=0.234 $X2=0 $Y2=0

* END of "./O2A1O1Ixp33_ASAP7_75t_L.pex.sp.O2A1O1IXP33_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

* File: O2A1O1Ixp5_ASAP7_75t_L.pex.sp
* Created: Tue Sep  5 12:46:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "O2A1O1Ixp5_ASAP7_75t_L.pex.sp.pex"
* BEGIN of "./O2A1O1Ixp5_ASAP7_75t_L.pex.sp.pex"
* File: O2A1O1Ixp5_ASAP7_75t_L.pex.sp.pex
* Created: Tue Sep  5 12:46:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_O2A1O1IXP5_ASAP7_75T_L%A1 2 5 8 11 13 25 28 31 32 33 34 37 43 46 49
+ VSS
c29 49 VSS 0.00793702f $X=0.018 $Y=0.135
c30 46 VSS 3.38114e-19 $X=0.243 $Y=0.106
c31 45 VSS 9.46734e-19 $X=0.243 $Y=0.099
c32 43 VSS 5.5624e-19 $X=0.243 $Y=0.135
c33 37 VSS 0.00350999f $X=0.081 $Y=0.135
c34 34 VSS 1.97726e-19 $X=0.1985 $Y=0.072
c35 33 VSS 7.004e-20 $X=0.163 $Y=0.072
c36 32 VSS 1.60995e-19 $X=0.148 $Y=0.072
c37 31 VSS 5.17397e-19 $X=0.144 $Y=0.072
c38 30 VSS 0.00202608f $X=0.126 $Y=0.072
c39 29 VSS 0.00302348f $X=0.095 $Y=0.072
c40 26 VSS 0.00205016f $X=0.027 $Y=0.072
c41 25 VSS 0.00199463f $X=0.234 $Y=0.072
c42 18 VSS 5.05955e-19 $X=0.018 $Y=0.116
c43 17 VSS 0.00120676f $X=0.018 $Y=0.106
c44 16 VSS 4.10062e-19 $X=0.018 $Y=0.126
c45 11 VSS 0.00105091f $X=0.243 $Y=0.135
c46 8 VSS 0.0607085f $X=0.243 $Y=0.0675
c47 2 VSS 0.0693372f $X=0.081 $Y=0.135
r48 45 46 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.099 $X2=0.243 $Y2=0.106
r49 43 46 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.106
r50 41 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.243 $Y2=0.099
r51 35 49 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r52 35 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.081 $Y2=0.135
r53 33 34 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.163
+ $Y=0.072 $X2=0.1985 $Y2=0.072
r54 32 33 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.072 $X2=0.163 $Y2=0.072
r55 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.148 $Y2=0.072
r56 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.144 $Y2=0.072
r57 29 30 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.072 $X2=0.126 $Y2=0.072
r58 28 29 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.067
+ $Y=0.072 $X2=0.095 $Y2=0.072
r59 26 28 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.072 $X2=0.067 $Y2=0.072
r60 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.072 $X2=0.243 $Y2=0.081
r61 25 34 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.1985 $Y2=0.072
r62 17 18 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.106 $X2=0.018 $Y2=0.116
r63 16 49 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.135
r64 16 18 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.116
r65 15 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.081 $X2=0.027 $Y2=0.072
r66 15 17 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.106
r67 11 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r68 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r69 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r70 2 37 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r71 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
.ends

.subckt PM_O2A1O1IXP5_ASAP7_75T_L%A2 2 5 8 11 13 17 23 25 VSS
c28 25 VSS 2.14622e-20 $X=0.135 $Y=0.147
c29 23 VSS 6.08933e-19 $X=0.139 $Y=0.15
c30 17 VSS 5.74468e-19 $X=0.135 $Y=0.135
c31 11 VSS 0.00313854f $X=0.189 $Y=0.135
c32 8 VSS 0.0626362f $X=0.189 $Y=0.0675
c33 2 VSS 0.0638717f $X=0.135 $Y=0.135
r34 24 25 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.147
r35 23 25 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.15 $X2=0.135 $Y2=0.147
r36 17 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r37 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r38 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r39 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r40 2 17 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r41 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
.ends

.subckt PM_O2A1O1IXP5_ASAP7_75T_L%B 2 5 7 10 VSS
c11 10 VSS 7.73504e-19 $X=0.296 $Y=0.128
c12 5 VSS 0.00125105f $X=0.297 $Y=0.135
c13 2 VSS 0.0610856f $X=0.297 $Y=0.0675
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_O2A1O1IXP5_ASAP7_75T_L%C 2 7 11 16 VSS
c12 16 VSS 0.0039869f $X=0.368 $Y=0.135
c13 11 VSS 0.00299117f $X=0.371 $Y=0.116
c14 2 VSS 0.0659251f $X=0.351 $Y=0.054
r15 15 16 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.368 $Y=0.135 $X2=0.368
+ $Y2=0.135
r16 11 15 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.368
+ $Y=0.116 $X2=0.368 $Y2=0.135
r17 5 16 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.368 $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r19 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.054 $X2=0.351 $Y2=0.135
.ends

.subckt PM_O2A1O1IXP5_ASAP7_75T_L%9 1 6 7 13 16 17 18 VSS
c12 19 VSS 9.71907e-19 $X=0.261 $Y=0.036
c13 18 VSS 0.0118667f $X=0.252 $Y=0.036
c14 17 VSS 0.00756655f $X=0.27 $Y=0.036
c15 16 VSS 0.00247812f $X=0.27 $Y=0.036
c16 13 VSS 0.00669097f $X=0.162 $Y=0.036
c17 6 VSS 5.945e-19 $X=0.287 $Y=0.0675
c18 1 VSS 5.05892e-19 $X=0.179 $Y=0.0675
r19 18 19 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.261 $Y2=0.036
r20 16 19 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.261 $Y2=0.036
r21 16 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r22 12 18 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.252 $Y2=0.036
r23 12 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r24 10 17 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r25 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r26 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r27 4 13 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r28 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.164 $Y2=0.0675
.ends

.subckt PM_O2A1O1IXP5_ASAP7_75T_L%Y 2 3 10 13 18 20 21 25 27 30 33 VSS
c15 39 VSS 0.00191594f $X=0.396 $Y=0.234
c16 38 VSS 0.00278493f $X=0.405 $Y=0.234
c17 33 VSS 0.00161166f $X=0.378 $Y=0.234
c18 31 VSS 2.98008e-19 $X=0.405 $Y=0.216
c19 30 VSS 6.54272e-19 $X=0.405 $Y=0.207
c20 29 VSS 6.80352e-19 $X=0.405 $Y=0.189
c21 28 VSS 2.45683e-19 $X=0.405 $Y=0.171
c22 27 VSS 0.00397351f $X=0.405 $Y=0.164
c23 26 VSS 0.00108941f $X=0.405 $Y=0.063
c24 25 VSS 0.00332962f $X=0.405 $Y=0.045
c25 23 VSS 7.30208e-19 $X=0.405 $Y=0.225
c26 21 VSS 0.00452798f $X=0.377 $Y=0.036
c27 20 VSS 0.00260728f $X=0.335 $Y=0.036
c28 18 VSS 0.00538096f $X=0.324 $Y=0.036
c29 15 VSS 0.00280886f $X=0.396 $Y=0.036
c30 13 VSS 0.00458137f $X=0.376 $Y=0.2025
c31 9 VSS 2.53915e-20 $X=0.324 $Y=0.0675
c32 4 VSS 6.14564e-19 $X=0.324 $Y=0.0455
r33 39 40 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.4005 $Y2=0.234
r34 38 40 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.234 $X2=0.4005 $Y2=0.234
r35 33 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r36 30 31 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.207 $X2=0.405 $Y2=0.216
r37 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.207
r38 28 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.171 $X2=0.405 $Y2=0.189
r39 27 28 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.164 $X2=0.405 $Y2=0.171
r40 26 27 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.063 $X2=0.405 $Y2=0.164
r41 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.063
r42 23 38 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.234
r43 23 31 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.216
r44 20 21 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.335
+ $Y=0.036 $X2=0.377 $Y2=0.036
r45 17 20 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.335 $Y2=0.036
r46 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r47 15 25 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.405 $Y2=0.036
r48 15 21 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.377 $Y2=0.036
r49 13 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r50 10 13 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.376 $Y2=0.2025
r51 9 18 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r52 3 4 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0455 $X2=0.324 $Y2=0.0455
r53 2 4 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.0455 $X2=0.324 $Y2=0.0455
r54 1 9 3.12934 $w=6.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.324
+ $Y=0.064 $X2=0.307 $Y2=0.064
r55 1 4 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.324 $Y=0.064 $X2=0.324 $Y2=0.0455
.ends


* END of "./O2A1O1Ixp5_ASAP7_75t_L.pex.sp.pex"
* 
.subckt O2A1O1Ixp5_ASAP7_75t_L  VSS VDD A1 A2 B C Y
* 
* Y	Y
* C	C
* B	B
* A2	A2
* A1	A1
M0 VSS N_A2_M0_g N_9_M0_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M1 N_9_M1_d N_A1_M1_g VSS VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M2 N_Y_M2_d N_B_M2_g N_9_M2_s VSS NMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 VSS N_C_M3_g N_Y_M3_s VSS NMOS_LVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341 $Y=0.027
M4 noxref_7 N_A1_M4_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 noxref_8 N_A2_M5_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 noxref_8 N_A2_M6_g noxref_7 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M7 noxref_7 N_A1_M7_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M8 noxref_8 N_B_M8_g VDD VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
M9 N_Y_M9_d N_C_M9_g noxref_8 VDD PMOS_LVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "O2A1O1Ixp5_ASAP7_75t_L.pex.sp.O2A1O1IXP5_ASAP7_75T_L.pxi"
* BEGIN of "./O2A1O1Ixp5_ASAP7_75t_L.pex.sp.O2A1O1IXP5_ASAP7_75T_L.pxi"
* File: O2A1O1Ixp5_ASAP7_75t_L.pex.sp.O2A1O1IXP5_ASAP7_75T_L.pxi
* Created: Tue Sep  5 12:46:56 2017
* 
x_PM_O2A1O1IXP5_ASAP7_75T_L%A1 N_A1_c_1_p N_A1_M4_g N_A1_M1_g N_A1_c_8_p
+ N_A1_M7_g N_A1_c_20_p A1 N_A1_c_3_p N_A1_c_9_p N_A1_c_24_p N_A1_c_6_p
+ N_A1_c_11_p N_A1_c_12_p N_A1_c_18_p N_A1_c_15_p VSS
+ PM_O2A1O1IXP5_ASAP7_75T_L%A1
x_PM_O2A1O1IXP5_ASAP7_75T_L%A2 N_A2_c_30_n N_A2_M5_g N_A2_M0_g N_A2_c_36_n
+ N_A2_M6_g N_A2_c_39_n A2 N_A2_c_44_n VSS PM_O2A1O1IXP5_ASAP7_75T_L%A2
x_PM_O2A1O1IXP5_ASAP7_75T_L%B N_B_M2_g N_B_c_59_n N_B_M8_g B VSS
+ PM_O2A1O1IXP5_ASAP7_75T_L%B
x_PM_O2A1O1IXP5_ASAP7_75T_L%C N_C_M3_g N_C_M9_g C N_C_c_73_n VSS
+ PM_O2A1O1IXP5_ASAP7_75T_L%C
x_PM_O2A1O1IXP5_ASAP7_75T_L%9 N_9_M0_s N_9_M2_s N_9_M1_d N_9_c_82_n N_9_c_92_p
+ N_9_c_84_n N_9_c_85_n VSS PM_O2A1O1IXP5_ASAP7_75T_L%9
x_PM_O2A1O1IXP5_ASAP7_75T_L%Y N_Y_M3_s N_Y_M2_d N_Y_M9_d N_Y_c_94_n N_Y_c_93_n
+ N_Y_c_107_n N_Y_c_97_n Y N_Y_c_99_n N_Y_c_104_n N_Y_c_100_n VSS
+ PM_O2A1O1IXP5_ASAP7_75T_L%Y
cc_1 N_A1_c_1_p N_A2_c_30_n 0.0036697f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_2 N_A1_M1_g N_A2_c_30_n 2.69148e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_3 N_A1_c_3_p N_A2_c_30_n 3.51973e-19 $X=0.144 $Y=0.072 $X2=0.135 $Y2=0.135
cc_4 N_A1_c_1_p N_A2_M0_g 3.03912e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_5 N_A1_M1_g N_A2_M0_g 0.00323392f $X=0.243 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_6 N_A1_c_6_p N_A2_M0_g 3.8965e-19 $X=0.1985 $Y=0.072 $X2=0.189 $Y2=0.0675
cc_7 N_A1_c_1_p N_A2_c_36_n 0.00122296f $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_8 N_A1_c_8_p N_A2_c_36_n 0.00121817f $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.135
cc_9 N_A1_c_9_p N_A2_c_36_n 7.17367e-19 $X=0.148 $Y=0.072 $X2=0.189 $Y2=0.135
cc_10 N_A1_c_3_p N_A2_c_39_n 0.00120736f $X=0.144 $Y=0.072 $X2=0.135 $Y2=0.135
cc_11 N_A1_c_11_p N_A2_c_39_n 8.78098e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_12 N_A1_c_12_p N_A2_c_39_n 6.84703e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_13 N_A1_c_9_p A2 3.82448e-19 $X=0.148 $Y=0.072 $X2=0.139 $Y2=0.15
cc_14 N_A1_c_12_p A2 2.76524e-19 $X=0.243 $Y=0.135 $X2=0.139 $Y2=0.15
cc_15 N_A1_c_15_p N_A2_c_44_n 3.90421e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.147
cc_16 N_A1_M1_g N_B_M2_g 0.0031831f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_17 N_A1_c_8_p N_B_c_59_n 8.86777e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_18 N_A1_c_18_p B 0.00306489f $X=0.243 $Y=0.106 $X2=0.189 $Y2=0.135
cc_19 N_A1_M1_g N_C_M3_g 2.63406e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_20 N_A1_c_20_p C 2.17364e-19 $X=0.234 $Y=0.072 $X2=0.189 $Y2=0.135
cc_21 VSS N_A1_c_9_p 4.65344e-19 $X=0.148 $Y=0.072 $X2=0 $Y2=0
cc_22 VSS N_A1_M1_g 3.62029e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_23 VSS N_A1_c_12_p 0.00123353f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_24 N_A1_c_24_p N_9_M0_s 2.87556e-19 $X=0.163 $Y=0.072 $X2=0.135 $Y2=0.135
cc_25 N_A1_c_24_p N_9_c_82_n 0.00156633f $X=0.163 $Y=0.072 $X2=0.189 $Y2=0.2025
cc_26 N_A1_c_6_p N_9_c_82_n 0.00109303f $X=0.1985 $Y=0.072 $X2=0.189 $Y2=0.2025
cc_27 N_A1_c_20_p N_9_c_84_n 0.00153136f $X=0.234 $Y=0.072 $X2=0.135 $Y2=0.135
cc_28 N_A1_M1_g N_9_c_85_n 2.34993e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_29 N_A1_c_24_p N_9_c_85_n 0.00931117f $X=0.163 $Y=0.072 $X2=0.135 $Y2=0.135
cc_30 N_A2_M0_g N_B_M2_g 2.34385e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_31 VSS A2 3.11986e-19 $X=0.139 $Y=0.15 $X2=0.081 $Y2=0.2025
cc_32 VSS N_A2_M0_g 2.64781e-19 $X=0.189 $Y=0.0675 $X2=0.018 $Y2=0.116
cc_33 VSS N_A2_c_30_n 2.38303e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_34 VSS N_A2_c_36_n 3.78279e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_35 VSS N_A2_c_36_n 8.00372e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_36 VSS A2 8.38539e-19 $X=0.139 $Y=0.15 $X2=0.081 $Y2=0.2025
cc_37 VSS N_A2_c_30_n 2.92813e-19 $X=0.135 $Y=0.135 $X2=0.018 $Y2=0.116
cc_38 VSS A2 0.0040524f $X=0.139 $Y=0.15 $X2=0.018 $Y2=0.116
cc_39 VSS N_A2_M0_g 3.99641e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_40 VSS N_A2_c_36_n 5.14484e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_41 N_A2_c_36_n N_9_c_82_n 8.00061e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.2025
cc_42 N_A2_M0_g N_9_c_85_n 2.64781e-19 $X=0.189 $Y=0.0675 $X2=0.018 $Y2=0.116
cc_43 N_B_M2_g N_C_M3_g 0.00354623f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_44 B C 0.00195119f $X=0.296 $Y=0.128 $X2=0.243 $Y2=0.135
cc_45 N_B_c_59_n N_C_c_73_n 0.00104216f $X=0.297 $Y=0.135 $X2=0.018 $Y2=0.126
cc_46 VSS N_B_M2_g 3.51973e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_47 VSS B 0.00120736f $X=0.296 $Y=0.128 $X2=0 $Y2=0
cc_48 B N_9_c_84_n 2.71261e-19 $X=0.296 $Y=0.128 $X2=0.018 $Y2=0.106
cc_49 B N_Y_c_93_n 2.97606e-19 $X=0.296 $Y=0.128 $X2=0.018 $Y2=0.116
cc_50 C N_Y_c_94_n 8.37647e-19 $X=0.371 $Y=0.116 $X2=0.243 $Y2=0.2025
cc_51 N_C_c_73_n N_Y_c_94_n 4.59187e-19 $X=0.368 $Y=0.135 $X2=0.243 $Y2=0.2025
cc_52 C N_Y_c_93_n 0.0015775f $X=0.371 $Y=0.116 $X2=0.018 $Y2=0.116
cc_53 N_C_M3_g N_Y_c_97_n 2.64781e-19 $X=0.351 $Y=0.054 $X2=0 $Y2=0
cc_54 C N_Y_c_97_n 0.00424763f $X=0.371 $Y=0.116 $X2=0 $Y2=0
cc_55 C N_Y_c_99_n 0.00861419f $X=0.371 $Y=0.116 $X2=0.067 $Y2=0.072
cc_56 C N_Y_c_100_n 2.86085e-19 $X=0.371 $Y=0.116 $X2=0.163 $Y2=0.072
cc_57 VSS N_9_c_82_n 0.00149637f $X=0.162 $Y=0.2025 $X2=0.243 $Y2=0.2025
cc_58 VSS N_Y_c_94_n 0.00363024f $X=0.324 $Y=0.2025 $X2=0.243 $Y2=0.2025
cc_59 VSS N_Y_c_94_n 3.95522e-19 $X=0.324 $Y=0.198 $X2=0.243 $Y2=0.2025
cc_60 VSS N_Y_c_93_n 0.00138157f $X=0.324 $Y=0.2025 $X2=0.018 $Y2=0.116
cc_61 VSS N_Y_c_104_n 3.44171e-19 $X=0.324 $Y=0.198 $X2=0.126 $Y2=0.072
cc_62 VSS N_Y_c_100_n 5.01727e-19 $X=0.324 $Y=0.2025 $X2=0.163 $Y2=0.072
cc_63 N_9_c_84_n N_Y_c_93_n 0.00342796f $X=0.27 $Y=0.036 $X2=0.018 $Y2=0.116
cc_64 N_9_c_92_p N_Y_c_107_n 6.82184e-19 $X=0.27 $Y=0.036 $X2=0 $Y2=0

* END of "./O2A1O1Ixp5_ASAP7_75t_L.pex.sp.O2A1O1IXP5_ASAP7_75T_L.pxi"
* 
*
.ends
*
*

