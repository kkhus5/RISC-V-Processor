* File: DFFHQNx1_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:24:08 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DFFHQNx1_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DFFHQNx1_ASAP7_75t_SRAM.pex.sp.pex"
* File: DFFHQNx1_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:24:08 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%CLK 2 5 7 12 14 VSS
c20 14 VSS 0.00674559f $X=0.081 $Y=0.135
c21 12 VSS 0.00682604f $X=0.082 $Y=0.119
c22 5 VSS 0.00206449f $X=0.081 $Y=0.135
c23 2 VSS 0.0629f $X=0.081 $Y=0.054
r24 12 14 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.135
r25 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r26 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r27 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%4 2 7 10 13 15 18 21 23 25 28 30 36 37 38 41 42
+ 45 52 59 67 68 70 72 73 78 79 83 88 VSS
c77 114 VSS 1.06551e-19 $X=0.03 $Y=0.153
c78 113 VSS 6.89947e-19 $X=0.027 $Y=0.153
c79 88 VSS 0.00102973f $X=0.675 $Y=0.135
c80 83 VSS 8.66895e-19 $X=0.405 $Y=0.135
c81 79 VSS 0.00121012f $X=0.151 $Y=0.135
c82 78 VSS 0.00390107f $X=0.151 $Y=0.135
c83 73 VSS 0.00263053f $X=0.601 $Y=0.153
c84 72 VSS 0.00556612f $X=0.527 $Y=0.153
c85 70 VSS 0.00405122f $X=0.675 $Y=0.153
c86 68 VSS 0.00330975f $X=0.29 $Y=0.153
c87 67 VSS 0.00602706f $X=0.175 $Y=0.153
c88 59 VSS 6.74716e-19 $X=0.033 $Y=0.153
c89 55 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c90 54 VSS 0.00180216f $X=0.047 $Y=0.234
c91 52 VSS 0.00250119f $X=0.054 $Y=0.234
c92 50 VSS 0.00305101f $X=0.027 $Y=0.234
c93 48 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c94 47 VSS 0.00199699f $X=0.047 $Y=0.036
c95 45 VSS 0.00250119f $X=0.054 $Y=0.036
c96 43 VSS 0.00305101f $X=0.027 $Y=0.036
c97 42 VSS 4.88707e-19 $X=0.018 $Y=0.2125
c98 41 VSS 0.00180713f $X=0.018 $Y=0.2
c99 40 VSS 4.69158e-19 $X=0.018 $Y=0.225
c100 38 VSS 0.00173342f $X=0.018 $Y=0.107
c101 37 VSS 9.57865e-19 $X=0.018 $Y=0.07
c102 36 VSS 0.00172854f $X=0.018 $Y=0.144
c103 33 VSS 0.00509483f $X=0.056 $Y=0.216
c104 30 VSS 2.98509e-19 $X=0.071 $Y=0.216
c105 28 VSS 0.00497933f $X=0.056 $Y=0.054
c106 25 VSS 2.98509e-19 $X=0.071 $Y=0.054
c107 21 VSS 0.00214819f $X=0.675 $Y=0.135
c108 18 VSS 0.0585656f $X=0.675 $Y=0.0405
c109 13 VSS 0.00214124f $X=0.405 $Y=0.135
c110 10 VSS 0.058827f $X=0.405 $Y=0.0675
c111 2 VSS 0.0628024f $X=0.135 $Y=0.054
r112 113 114 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r113 110 113 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r114 78 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.151 $Y=0.135 $X2=0.151
+ $Y2=0.135
r115 72 73 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.601 $Y2=0.153
r116 70 73 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.675
+ $Y=0.153 $X2=0.601 $Y2=0.153
r117 70 88 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.675 $Y=0.153 $X2=0.675
+ $Y2=0.153
r118 67 68 7.80864 $w=1.8e-08 $l=1.15e-07 $layer=M2 $thickness=3.6e-08 $X=0.175
+ $Y=0.153 $X2=0.29 $Y2=0.153
r119 65 72 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.527 $Y2=0.153
r120 65 68 7.80864 $w=1.8e-08 $l=1.15e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.29 $Y2=0.153
r121 65 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r122 62 67 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.151
+ $Y=0.153 $X2=0.175 $Y2=0.153
r123 62 79 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.151 $Y=0.153 $X2=0.151
+ $Y2=0.153
r124 59 114 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r125 58 62 8.01235 $w=1.8e-08 $l=1.18e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.151 $Y2=0.153
r126 58 59 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r127 54 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r128 52 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r129 50 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r130 47 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r131 45 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r132 43 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r133 41 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r134 40 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r135 40 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r136 39 110 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r137 39 41 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.2
r138 37 38 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.107
r139 36 110 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r140 36 38 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.107
r141 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r142 35 37 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r143 33 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r144 30 33 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r145 28 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r146 25 28 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r147 21 88 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.135 $X2=0.675
+ $Y2=0.135
r148 21 23 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2295
r149 18 21 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.135
r150 13 83 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r151 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2295
r152 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r153 5 78 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.151 $Y2=0.135
r154 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r155 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%D 2 5 7 10 12 14 21 23 28 VSS
c18 28 VSS 0.00931225f $X=0.243 $Y=0.135
c19 24 VSS 2.45662e-20 $X=0.276 $Y=0.135
c20 23 VSS 0.00111822f $X=0.271 $Y=0.135
c21 21 VSS 2.56376e-19 $X=0.281 $Y=0.135
c22 14 VSS 2.7811e-19 $X=0.243 $Y=0.116
c23 12 VSS 0.00925957f $X=0.244 $Y=0.082
c24 10 VSS 2.38113e-19 $X=0.243 $Y=0.126
c25 5 VSS 0.00522238f $X=0.297 $Y=0.135
c26 2 VSS 0.0630392f $X=0.297 $Y=0.0675
r27 23 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.271
+ $Y=0.135 $X2=0.276 $Y2=0.135
r28 21 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.281
+ $Y=0.135 $X2=0.276 $Y2=0.135
r29 21 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.281 $Y=0.135 $X2=0.281
+ $Y2=0.135
r30 19 28 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.243 $Y2=0.135
r31 19 23 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.271 $Y2=0.135
r32 13 14 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.106 $X2=0.243 $Y2=0.116
r33 12 13 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.082 $X2=0.243 $Y2=0.106
r34 10 28 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.135
r35 10 14 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.116
r36 5 22 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.281 $Y2=0.135
r37 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r38 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%6 2 5 8 14 17 20 23 28 35 39 44 50 55 57 61 66
+ 67 68 75 77 78 87 89 105 110 111 113 114 VSS
c102 114 VSS 2.23151e-19 $X=0.324 $Y=0.178
c103 113 VSS 4.08645e-19 $X=0.324 $Y=0.167
c104 111 VSS 7.77947e-19 $X=0.189 $Y=0.167
c105 110 VSS 9.60988e-19 $X=0.189 $Y=0.106
c106 105 VSS 6.81413e-19 $X=0.513 $Y=0.18
c107 89 VSS 0.0113851f $X=0.513 $Y=0.189
c108 87 VSS 0.00141172f $X=0.324 $Y=0.189
c109 78 VSS 4.01771e-19 $X=0.342 $Y=0.135
c110 77 VSS 5.28662e-19 $X=0.333 $Y=0.135
c111 75 VSS 7.4105e-19 $X=0.351 $Y=0.135
c112 68 VSS 0.00169555f $X=0.18 $Y=0.234
c113 67 VSS 9.43175e-19 $X=0.189 $Y=0.225
c114 66 VSS 0.00196236f $X=0.189 $Y=0.234
c115 61 VSS 0.00196921f $X=0.162 $Y=0.234
c116 57 VSS 0.00170883f $X=0.18 $Y=0.036
c117 55 VSS 0.00196236f $X=0.189 $Y=0.036
c118 50 VSS 0.00193426f $X=0.162 $Y=0.036
c119 47 VSS 0.00715944f $X=0.16 $Y=0.216
c120 42 VSS 0.00719538f $X=0.16 $Y=0.054
c121 35 VSS 0.0611368f $X=0.725 $Y=0.178
c122 28 VSS 0.00126548f $X=0.464 $Y=0.178
c123 20 VSS 0.0618767f $X=0.729 $Y=0.178
c124 17 VSS 1.08457e-19 $X=0.621 $Y=0.178
c125 14 VSS 0.0600454f $X=0.621 $Y=0.0405
c126 8 VSS 0.0602427f $X=0.459 $Y=0.0405
c127 2 VSS 0.0623279f $X=0.351 $Y=0.135
r128 113 114 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.324 $Y=0.167 $X2=0.324 $Y2=0.178
r129 110 111 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.106 $X2=0.189 $Y2=0.167
r130 104 105 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r131 89 105 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r132 87 114 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.189 $X2=0.324 $Y2=0.178
r133 86 89 12.8333 $w=1.8e-08 $l=1.89e-07 $layer=M2 $thickness=3.6e-08 $X=0.324
+ $Y=0.189 $X2=0.513 $Y2=0.189
r134 86 87 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.324 $Y=0.189 $X2=0.324
+ $Y2=0.189
r135 83 111 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.167
r136 82 86 9.16667 $w=1.8e-08 $l=1.35e-07 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.324 $Y2=0.189
r137 82 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.189 $X2=0.189
+ $Y2=0.189
r138 77 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.135 $X2=0.342 $Y2=0.135
r139 75 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.342 $Y2=0.135
r140 72 113 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.144 $X2=0.324 $Y2=0.167
r141 71 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.135 $X2=0.333 $Y2=0.135
r142 71 72 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.135 $X2=0.324 $Y2=0.144
r143 68 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r144 67 83 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.189
r145 66 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r146 66 67 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.189 $Y2=0.225
r147 61 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r148 57 58 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r149 56 110 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.106
r150 55 58 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r151 55 56 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r152 50 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r153 47 61 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r154 44 47 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r155 42 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r156 39 42 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r157 28 104 39.0385 $w=2.6e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.178 $X2=0.513 $Y2=0.178
r158 20 35 3.07692 $w=2.6e-08 $l=4e-09 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.178 $X2=0.725 $Y2=0.178
r159 20 23 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.178 $X2=0.729 $Y2=0.2295
r160 17 35 82.8571 $w=2.6e-08 $l=1.04e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.725 $Y2=0.178
r161 17 104 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.513 $Y2=0.178
r162 14 17 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0405 $X2=0.621 $Y2=0.178
r163 11 28 3.84615 $w=2.6e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.178 $X2=0.464 $Y2=0.178
r164 8 11 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.178
r165 2 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r166 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%7 2 5 7 9 10 13 14 17 19 22 29 30 31 38 43 44 45
+ 46 47 48 52 53 VSS
c43 54 VSS 3.52511e-19 $X=0.612 $Y=0.09
c44 53 VSS 1.80704e-19 $X=0.603 $Y=0.09
c45 52 VSS 5.96246e-19 $X=0.621 $Y=0.09
c46 49 VSS 6.86664e-19 $X=0.621 $Y=0.224
c47 48 VSS 4.95788e-19 $X=0.621 $Y=0.203
c48 47 VSS 1.19762e-19 $X=0.621 $Y=0.167
c49 46 VSS 3.19764e-19 $X=0.621 $Y=0.165
c50 45 VSS 3.13056e-19 $X=0.621 $Y=0.14
c51 44 VSS 3.62783e-19 $X=0.621 $Y=0.122
c52 43 VSS 1.48552e-19 $X=0.621 $Y=0.101
c53 38 VSS 0.00113884f $X=0.594 $Y=0.054
c54 31 VSS 0.00668633f $X=0.612 $Y=0.234
c55 30 VSS 3.5821e-19 $X=0.5805 $Y=0.09
c56 29 VSS 0.00257846f $X=0.576 $Y=0.09
c57 24 VSS 1.48201e-19 $X=0.585 $Y=0.09
c58 22 VSS 0.0179338f $X=0.65 $Y=0.2295
c59 19 VSS 3.14771e-19 $X=0.665 $Y=0.2295
c60 17 VSS 2.67274e-19 $X=0.592 $Y=0.2295
c61 13 VSS 0.0252201f $X=0.594 $Y=0.0405
c62 9 VSS 6.29543e-19 $X=0.611 $Y=0.0405
c63 5 VSS 0.00238279f $X=0.513 $Y=0.09
c64 2 VSS 0.0584396f $X=0.513 $Y=0.0405
r65 53 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.603
+ $Y=0.09 $X2=0.612 $Y2=0.09
r66 52 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.612 $Y2=0.09
r67 51 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.09 $X2=0.603 $Y2=0.09
r68 49 50 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.224 $X2=0.621 $Y2=0.2245
r69 48 49 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.224
r70 47 48 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.203
r71 46 47 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.167
r72 45 46 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r73 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r74 43 44 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.101 $X2=0.621 $Y2=0.122
r75 42 50 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.2245
r76 41 52 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.09
r77 41 43 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.101
r78 36 51 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.09
r79 36 38 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.054
r80 31 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r81 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r82 29 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.09 $X2=0.5805 $Y2=0.09
r83 26 29 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.09 $X2=0.576 $Y2=0.09
r84 24 51 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.594 $Y2=0.09
r85 24 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.5805 $Y2=0.09
r86 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2295 $X2=0.65 $Y2=0.2295
r87 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.592
+ $Y=0.2295 $X2=0.65 $Y2=0.2295
r88 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r89 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r90 13 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.054 $X2=0.594
+ $Y2=0.054
r91 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.594 $Y2=0.0405
r92 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0405 $X2=0.594 $Y2=0.0405
r93 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.09 $X2=0.513
+ $Y2=0.09
r94 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.09 $X2=0.513 $Y2=0.2295
r95 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.09
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%8 2 5 7 9 14 17 21 22 25 27 33 35 37 38 39 41 43
+ 44 45 46 50 52 53 54 55 59 62 65 VSS
c53 65 VSS 2.85958e-19 $X=0.459 $Y=0.131
c54 62 VSS 0.00341346f $X=0.45 $Y=0.036
c55 61 VSS 0.0025252f $X=0.459 $Y=0.036
c56 59 VSS 0.00276391f $X=0.432 $Y=0.036
c57 55 VSS 4.23521e-19 $X=0.5445 $Y=0.131
c58 54 VSS 3.49205e-20 $X=0.522 $Y=0.131
c59 53 VSS 2.00095e-19 $X=0.504 $Y=0.131
c60 52 VSS 0.00133241f $X=0.496 $Y=0.131
c61 50 VSS 2.94642e-19 $X=0.567 $Y=0.131
c62 47 VSS 4.32029e-19 $X=0.459 $Y=0.214
c63 46 VSS 2.06877e-19 $X=0.459 $Y=0.203
c64 45 VSS 6.09344e-21 $X=0.459 $Y=0.167
c65 44 VSS 2.12612e-19 $X=0.459 $Y=0.165
c66 43 VSS 2.51143e-19 $X=0.459 $Y=0.225
c67 41 VSS 3.68971e-19 $X=0.459 $Y=0.114
c68 40 VSS 3.4692e-19 $X=0.459 $Y=0.106
c69 38 VSS 7.88894e-19 $X=0.459 $Y=0.081
c70 37 VSS 2.0833e-19 $X=0.459 $Y=0.122
c71 35 VSS 0.00142907f $X=0.434 $Y=0.234
c72 34 VSS 3.2912e-19 $X=0.418 $Y=0.234
c73 33 VSS 0.00146362f $X=0.414 $Y=0.234
c74 32 VSS 0.00227054f $X=0.396 $Y=0.234
c75 27 VSS 0.00148441f $X=0.378 $Y=0.234
c76 25 VSS 0.00389542f $X=0.45 $Y=0.234
c77 24 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c78 21 VSS 0.00379676f $X=0.378 $Y=0.2025
c79 18 VSS 1.15515e-19 $X=0.3735 $Y=0.216
c80 16 VSS 5.70081e-19 $X=0.432 $Y=0.0405
c81 10 VSS 7.61325e-20 $X=0.4275 $Y=0.054
c82 5 VSS 0.0022736f $X=0.567 $Y=0.1305
c83 2 VSS 0.0591678f $X=0.567 $Y=0.0405
r84 62 63 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r85 61 63 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r86 58 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r87 58 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r88 54 55 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r89 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r90 52 53 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.496
+ $Y=0.131 $X2=0.504 $Y2=0.131
r91 50 55 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r92 48 65 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r93 48 52 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.496 $Y2=0.131
r94 46 47 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.203 $X2=0.459 $Y2=0.214
r95 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.167 $X2=0.459 $Y2=0.203
r96 44 45 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.167
r97 43 47 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r98 42 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r99 42 44 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.165
r100 40 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.106 $X2=0.459 $Y2=0.114
r101 39 40 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.099 $X2=0.459 $Y2=0.106
r102 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.099
r103 37 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r104 37 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.114
r105 36 61 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r106 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.081
r107 34 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.234 $X2=0.434 $Y2=0.234
r108 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.418 $Y2=0.234
r109 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r110 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r111 25 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r112 25 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.434 $Y2=0.234
r113 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r114 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r115 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r116 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r117 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r118 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r119 13 59 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r120 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r121 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r122 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r123 5 50 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.131 $X2=0.567
+ $Y2=0.131
r124 5 7 370.904 $w=2e-08 $l=9.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1305 $X2=0.567 $Y2=0.2295
r125 2 5 337.185 $w=2e-08 $l=9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.1305
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%9 2 5 7 9 14 21 25 26 30 31 32 33 34 39 40 42 43
+ 44 45 46 VSS
c26 46 VSS 1.15795e-19 $X=0.945 $Y=0.171
c27 45 VSS 9.70265e-19 $X=0.945 $Y=0.167
c28 44 VSS 8.8218e-19 $X=0.945 $Y=0.117
c29 43 VSS 0.00183078f $X=0.945 $Y=0.09
c30 42 VSS 0.00237212f $X=0.945 $Y=0.225
c31 40 VSS 0.0018377f $X=0.918 $Y=0.234
c32 39 VSS 0.00568507f $X=0.9 $Y=0.234
c33 34 VSS 0.00462933f $X=0.936 $Y=0.234
c34 33 VSS 0.00189638f $X=0.9 $Y=0.036
c35 32 VSS 0.0035379f $X=0.882 $Y=0.036
c36 31 VSS 0.00146362f $X=0.846 $Y=0.036
c37 30 VSS 0.00510392f $X=0.828 $Y=0.036
c38 26 VSS 0.00226308f $X=0.792 $Y=0.036
c39 25 VSS 0.00657446f $X=0.936 $Y=0.036
c40 21 VSS 0.00122443f $X=0.783 $Y=0.105
c41 17 VSS 0.00481511f $X=0.862 $Y=0.2295
c42 12 VSS 0.00513464f $X=0.862 $Y=0.0405
c43 5 VSS 0.00277722f $X=0.783 $Y=0.1055
c44 2 VSS 0.0590816f $X=0.783 $Y=0.0405
r45 45 46 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.167 $X2=0.945 $Y2=0.171
r46 44 45 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.117 $X2=0.945 $Y2=0.167
r47 43 44 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.09 $X2=0.945 $Y2=0.117
r48 42 46 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.171
r49 41 43 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.09
r50 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.234 $X2=0.918 $Y2=0.234
r51 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.9 $Y2=0.234
r52 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r53 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.918 $Y2=0.234
r54 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r55 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.846 $Y2=0.036
r56 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r57 28 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.846 $Y2=0.036
r58 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.036 $X2=0.828 $Y2=0.036
r59 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r60 25 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.9 $Y2=0.036
r61 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.783 $Y=0.045 $X2=0.792 $Y2=0.036
r62 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.105
r63 17 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234 $X2=0.864
+ $Y2=0.234
r64 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2295 $X2=0.862 $Y2=0.2295
r65 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036 $X2=0.864
+ $Y2=0.036
r66 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.862 $Y2=0.0405
r67 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.105 $X2=0.783
+ $Y2=0.105
r68 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.1055 $X2=0.783 $Y2=0.2295
r69 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.1055
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%10 2 7 10 15 17 18 21 22 23 26 27 32 33 35 37 38
+ 39 40 41 43 44 46 47 50 57 58 66 69 73 76 84 VSS
c57 84 VSS 0.00206151f $X=0.999 $Y=0.135
c58 76 VSS 0.0077122f $X=0.999 $Y=0.153
c59 73 VSS 0.00149995f $X=0.891 $Y=0.153
c60 70 VSS 4.17512e-19 $X=0.837 $Y=0.162
c61 69 VSS 1.52743e-19 $X=0.729 $Y=0.162
c62 66 VSS 0.00357121f $X=0.72 $Y=0.233
c63 65 VSS 0.00257308f $X=0.729 $Y=0.233
c64 58 VSS 4.30636e-19 $X=0.866 $Y=0.162
c65 57 VSS 1.23291e-19 $X=0.85 $Y=0.162
c66 55 VSS 2.75449e-19 $X=0.882 $Y=0.162
c67 50 VSS 3.94906e-19 $X=0.837 $Y=0.135
c68 47 VSS 3.26354e-19 $X=0.792 $Y=0.162
c69 46 VSS 0.00206921f $X=0.774 $Y=0.162
c70 44 VSS 0.00191548f $X=0.828 $Y=0.162
c71 43 VSS 0.00132112f $X=0.729 $Y=0.224
c72 41 VSS 1.52884e-19 $X=0.729 $Y=0.136
c73 40 VSS 2.77769e-19 $X=0.729 $Y=0.119
c74 39 VSS 1.41609e-19 $X=0.729 $Y=0.101
c75 38 VSS 3.52175e-19 $X=0.729 $Y=0.081
c76 37 VSS 2.73935e-19 $X=0.729 $Y=0.153
c77 35 VSS 0.00166757f $X=0.704 $Y=0.036
c78 34 VSS 4.5779e-19 $X=0.688 $Y=0.036
c79 33 VSS 0.00146362f $X=0.684 $Y=0.036
c80 32 VSS 0.00375563f $X=0.666 $Y=0.036
c81 27 VSS 0.00409736f $X=0.72 $Y=0.036
c82 26 VSS 0.00133398f $X=0.702 $Y=0.2295
c83 22 VSS 6.50675e-19 $X=0.719 $Y=0.2295
c84 21 VSS 0.0376609f $X=0.648 $Y=0.0405
c85 17 VSS 5.63046e-19 $X=0.665 $Y=0.0405
c86 13 VSS 0.00322417f $X=0.999 $Y=0.135
c87 10 VSS 0.0656618f $X=0.999 $Y=0.0675
c88 5 VSS 0.00239735f $X=0.837 $Y=0.135
c89 2 VSS 0.0618222f $X=0.837 $Y=0.0405
r90 76 84 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.999 $Y=0.153 $X2=0.999
+ $Y2=0.153
r91 72 76 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.999 $Y2=0.153
r92 72 73 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r93 66 67 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.233 $X2=0.7245 $Y2=0.233
r94 65 67 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.233 $X2=0.7245 $Y2=0.233
r95 62 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.233 $X2=0.72 $Y2=0.233
r96 57 58 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.85
+ $Y=0.162 $X2=0.866 $Y2=0.162
r97 56 70 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.837 $Y2=0.162
r98 56 57 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.85 $Y2=0.162
r99 55 73 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.891 $Y2=0.162
r100 55 58 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.866 $Y2=0.162
r101 48 70 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.162
r102 48 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.135
r103 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.162 $X2=0.792 $Y2=0.162
r104 45 69 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.729 $Y2=0.162
r105 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.774 $Y2=0.162
r106 44 70 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.837 $Y2=0.162
r107 44 47 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.792 $Y2=0.162
r108 43 65 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.224 $X2=0.729 $Y2=0.233
r109 42 69 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.162
r110 42 43 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.224
r111 40 41 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.119 $X2=0.729 $Y2=0.136
r112 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.101 $X2=0.729 $Y2=0.119
r113 38 39 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.081 $X2=0.729 $Y2=0.101
r114 37 69 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.162
r115 37 41 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.136
r116 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.045 $X2=0.729 $Y2=0.081
r117 34 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.036 $X2=0.704 $Y2=0.036
r118 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.688 $Y2=0.036
r119 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.684 $Y2=0.036
r120 29 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.666 $Y2=0.036
r121 27 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.036 $X2=0.729 $Y2=0.045
r122 27 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.704 $Y2=0.036
r123 26 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.233
+ $X2=0.702 $Y2=0.233
r124 23 26 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2295 $X2=0.702 $Y2=0.2295
r125 22 26 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2295 $X2=0.702 $Y2=0.2295
r126 21 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r127 18 21 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0405 $X2=0.648 $Y2=0.0405
r128 17 21 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r129 13 84 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.135 $X2=0.999
+ $Y2=0.135
r130 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.135 $X2=0.999 $Y2=0.2025
r131 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.135
r132 5 50 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.135 $X2=0.837
+ $Y2=0.135
r133 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.2295
r134 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.0405 $X2=0.837 $Y2=0.135
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%QN 1 6 12 14 15 16 19 22 30 VSS
c7 30 VSS 0.00418221f $X=1.044 $Y=0.234
c8 29 VSS 0.00278493f $X=1.053 $Y=0.234
c9 22 VSS 0.00418221f $X=1.044 $Y=0.036
c10 21 VSS 0.00278493f $X=1.053 $Y=0.036
c11 19 VSS 0.00646415f $X=1.026 $Y=0.036
c12 16 VSS 0.00348361f $X=1.053 $Y=0.167
c13 15 VSS 0.00213993f $X=1.053 $Y=0.09
c14 12 VSS 0.00270985f $X=1.053 $Y=0.225
c15 9 VSS 0.00695792f $X=1.024 $Y=0.2025
c16 4 VSS 3.7894e-19 $X=1.024 $Y=0.0675
r17 30 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.234 $X2=1.0485 $Y2=0.234
r18 29 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.234 $X2=1.0485 $Y2=0.234
r19 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.234 $X2=1.044 $Y2=0.234
r20 22 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=1.0485 $Y2=0.036
r21 21 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.036 $X2=1.0485 $Y2=0.036
r22 18 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.036 $X2=1.044 $Y2=0.036
r23 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.036 $X2=1.026
+ $Y2=0.036
r24 15 16 5.22839 $w=1.8e-08 $l=7.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.09 $X2=1.053 $Y2=0.167
r25 14 16 3.80247 $w=1.8e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.223 $X2=1.053 $Y2=0.167
r26 12 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.225 $X2=1.053 $Y2=0.234
r27 12 14 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.225 $X2=1.053 $Y2=0.223
r28 11 21 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.045 $X2=1.053 $Y2=0.036
r29 11 15 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.045 $X2=1.053 $Y2=0.09
r30 9 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.234 $X2=1.026
+ $Y2=0.234
r31 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=1.009
+ $Y=0.2025 $X2=1.024 $Y2=0.2025
r32 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.026
+ $Y=0.0675 $X2=1.026 $Y2=0.036
r33 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.009
+ $Y=0.0675 $X2=1.024 $Y2=0.0675
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%12 1 6 9 VSS
c6 9 VSS 0.0270172f $X=0.38 $Y=0.0675
c7 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c8 4 VSS 3.25039e-19 $X=0.322 $Y=0.0675
r9 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r10 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%13 1 6 9 VSS
c10 9 VSS 0.0209308f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.6182e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%14 1 6 9 VSS
c8 9 VSS 0.0191671f $X=0.758 $Y=0.0405
c9 6 VSS 3.14771e-19 $X=0.773 $Y=0.0405
c10 4 VSS 2.6194e-19 $X=0.7 $Y=0.0405
r11 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r12 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.7
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r13 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.685
+ $Y=0.0405 $X2=0.7 $Y2=0.0405
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%15 1 2 VSS
c0 1 VSS 0.00225696f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%16 1 2 VSS
c3 1 VSS 0.00231486f $X=0.341 $Y=0.2025
r4 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends

.subckt PM_DFFHQNX1_ASAP7_75T_SRAM%17 1 2 VSS
c0 1 VSS 0.00219822f $X=0.773 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2295 $X2=0.739 $Y2=0.2295
.ends


* END of "./DFFHQNx1_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DFFHQNx1_ASAP7_75t_SRAM  VSS VDD CLK D QN
* 
* QN	QN
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_12_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_4_M3_g N_12_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_15_M4_d N_6_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_15_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_10_M7_d N_6_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.611
+ $Y=0.027
M8 N_14_M8_d N_4_M8_g N_10_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M9 VSS N_9_M9_g N_14_M9_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_9_M10_d N_10_M10_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.027
M11 N_QN_M11_d N_10_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M12 VDD N_CLK_M12_g N_4_M12_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M13 N_6_M13_d N_4_M13_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M14 N_16_M14_d N_D_M14_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M15 N_8_M15_d N_6_M15_g N_16_M15_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M16 N_13_M16_d N_4_M16_g N_8_M16_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M17 VDD N_7_M17_g N_13_M17_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M18 N_7_M18_d N_8_M18_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M19 N_10_M19_d N_4_M19_g N_7_M19_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.665 $Y=0.216
M20 N_17_M20_d N_6_M20_g N_10_M20_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.719 $Y=0.216
M21 VDD N_9_M21_g N_17_M21_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M22 N_9_M22_d N_10_M22_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.216
M23 N_QN_M23_d N_10_M23_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
*
* 
* .include "DFFHQNx1_ASAP7_75t_SRAM.pex.sp.DFFHQNX1_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DFFHQNx1_ASAP7_75t_SRAM.pex.sp.DFFHQNX1_ASAP7_75T_SRAM.pxi"
* File: DFFHQNx1_ASAP7_75t_SRAM.pex.sp.DFFHQNX1_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:24:08 2017
* 
x_PM_DFFHQNX1_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_13_p N_CLK_M12_g CLK
+ N_CLK_c_6_p VSS PM_DFFHQNX1_ASAP7_75T_SRAM%CLK
x_PM_DFFHQNX1_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M13_g N_4_M3_g N_4_c_43_p N_4_M16_g
+ N_4_M8_g N_4_c_48_p N_4_M19_g N_4_M0_s N_4_c_22_n N_4_M12_s N_4_c_23_n
+ N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_28_n N_4_c_29_n N_4_c_30_n
+ N_4_c_31_n N_4_c_40_p N_4_c_49_p N_4_c_37_p N_4_c_69_p N_4_c_33_n N_4_c_34_n
+ N_4_c_39_p N_4_c_51_p VSS PM_DFFHQNX1_ASAP7_75T_SRAM%4
x_PM_DFFHQNX1_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_99_n N_D_M14_g N_D_c_113_p D
+ N_D_c_101_n N_D_c_109_p N_D_c_102_n N_D_c_103_n VSS PM_DFFHQNX1_ASAP7_75T_SRAM%D
x_PM_DFFHQNX1_ASAP7_75T_SRAM%6 N_6_c_121_n N_6_M15_g N_6_M4_g N_6_M7_g N_6_c_171_p
+ N_6_c_125_n N_6_M20_g N_6_c_183_p N_6_c_126_n N_6_M1_d N_6_M13_d N_6_c_116_n
+ N_6_c_149_n N_6_c_132_n N_6_c_117_n N_6_c_150_n N_6_c_118_n N_6_c_135_n
+ N_6_c_136_n N_6_c_137_n N_6_c_138_n N_6_c_139_n N_6_c_119_n N_6_c_142_n
+ N_6_c_120_n N_6_c_143_n N_6_c_145_n N_6_c_188_p VSS PM_DFFHQNX1_ASAP7_75T_SRAM%6
x_PM_DFFHQNX1_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_244_p N_7_M17_g N_7_M7_s N_7_M6_d
+ N_7_c_228_n N_7_M18_d N_7_c_229_n N_7_M19_s N_7_c_231_n N_7_c_241_p
+ N_7_c_219_n N_7_c_220_n N_7_c_243_p N_7_c_260_p N_7_c_221_n N_7_c_246_p
+ N_7_c_222_n N_7_c_236_n N_7_c_237_n N_7_c_239_n N_7_c_223_n VSS
+ PM_DFFHQNX1_ASAP7_75T_SRAM%7
x_PM_DFFHQNX1_ASAP7_75T_SRAM%8 N_8_M6_g N_8_c_262_n N_8_M18_g N_8_M3_d N_8_M4_s
+ N_8_M15_d N_8_c_264_n N_8_M16_s N_8_c_310_p N_8_c_276_n N_8_c_265_n
+ N_8_c_311_p N_8_c_267_n N_8_c_283_n N_8_c_284_n N_8_c_268_n N_8_c_312_p
+ N_8_c_269_n N_8_c_286_n N_8_c_288_n N_8_c_302_n N_8_c_271_n N_8_c_303_n
+ N_8_c_272_n N_8_c_295_n N_8_c_273_n N_8_c_274_n N_8_c_275_n VSS
+ PM_DFFHQNX1_ASAP7_75T_SRAM%8
x_PM_DFFHQNX1_ASAP7_75T_SRAM%9 N_9_M9_g N_9_c_320_p N_9_M21_g N_9_M10_d N_9_M22_d
+ N_9_c_319_p N_9_c_331_p N_9_c_318_p N_9_c_323_p N_9_c_317_p N_9_c_327_p
+ N_9_c_329_p N_9_c_338_p N_9_c_328_p N_9_c_332_p N_9_c_322_p N_9_c_336_p
+ N_9_c_334_p N_9_c_330_p N_9_c_335_p VSS PM_DFFHQNX1_ASAP7_75T_SRAM%9
x_PM_DFFHQNX1_ASAP7_75T_SRAM%10 N_10_M10_g N_10_M22_g N_10_M11_g N_10_M23_g
+ N_10_M8_s N_10_M7_d N_10_c_340_n N_10_M20_s N_10_M19_d N_10_c_350_n
+ N_10_c_372_n N_10_c_341_n N_10_c_342_n N_10_c_394_p N_10_c_344_n N_10_c_364_n
+ N_10_c_351_n N_10_c_345_n N_10_c_352_n N_10_c_353_n N_10_c_377_n N_10_c_355_n
+ N_10_c_378_n N_10_c_380_n N_10_c_381_n N_10_c_382_n N_10_c_356_n N_10_c_357_n
+ N_10_c_383_n N_10_c_346_n N_10_c_388_n VSS PM_DFFHQNX1_ASAP7_75T_SRAM%10
x_PM_DFFHQNX1_ASAP7_75T_SRAM%QN N_QN_M11_d N_QN_M23_d N_QN_c_397_n QN N_QN_c_398_n
+ N_QN_c_401_n N_QN_c_403_n N_QN_c_399_n N_QN_c_400_n VSS
+ PM_DFFHQNX1_ASAP7_75T_SRAM%QN
x_PM_DFFHQNX1_ASAP7_75T_SRAM%12 N_12_M2_d N_12_M3_s N_12_c_404_n VSS
+ PM_DFFHQNX1_ASAP7_75T_SRAM%12
x_PM_DFFHQNX1_ASAP7_75T_SRAM%13 N_13_M16_d N_13_M17_s N_13_c_411_n VSS
+ PM_DFFHQNX1_ASAP7_75T_SRAM%13
x_PM_DFFHQNX1_ASAP7_75T_SRAM%14 N_14_M8_d N_14_M9_s N_14_c_420_n VSS
+ PM_DFFHQNX1_ASAP7_75T_SRAM%14
x_PM_DFFHQNX1_ASAP7_75T_SRAM%15 N_15_M5_s N_15_M4_d VSS PM_DFFHQNX1_ASAP7_75T_SRAM%15
x_PM_DFFHQNX1_ASAP7_75T_SRAM%16 N_16_M15_s N_16_M14_d VSS
+ PM_DFFHQNX1_ASAP7_75T_SRAM%16
x_PM_DFFHQNX1_ASAP7_75T_SRAM%17 N_17_M21_s N_17_M20_d VSS
+ PM_DFFHQNX1_ASAP7_75T_SRAM%17
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_22_n 3.57152e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 CLK N_4_c_23_n 0.00136255f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.144
cc_4 CLK N_4_c_24_n 2.75361e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.07
cc_5 CLK N_4_c_25_n 0.00136255f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.107
cc_6 N_CLK_c_6_p N_4_c_26_n 0.00145637f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2
cc_7 N_CLK_c_6_p N_4_c_27_n 2.75361e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2125
cc_8 CLK N_4_c_28_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_6_p N_4_c_29_n 5.03453e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_6_p N_4_c_30_n 0.00123168f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.153
cc_11 CLK N_4_c_31_n 4.93618e-19 $X=0.082 $Y=0.119 $X2=0.175 $Y2=0.153
cc_12 N_CLK_c_6_p N_4_c_31_n 0.00162391f $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_13 N_CLK_c_13_p N_4_c_33_n 0.00115059f $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.135
cc_14 CLK N_4_c_34_n 0.00174864f $X=0.082 $Y=0.119 $X2=0.151 $Y2=0.135
cc_15 N_CLK_c_6_p N_4_c_34_n 3.32041e-19 $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.135
cc_16 CLK N_6_c_116_n 6.37157e-19 $X=0.082 $Y=0.119 $X2=0.027 $Y2=0.234
cc_17 N_CLK_c_6_p N_6_c_117_n 6.45547e-19 $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.153
cc_18 N_CLK_c_6_p N_6_c_118_n 0.00125366f $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_19 N_CLK_c_6_p N_6_c_119_n 4.3806e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_20 CLK N_6_c_120_n 0.00137619f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.153
cc_21 N_4_M3_g N_D_M2_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_22 N_4_c_37_p N_D_c_99_n 2.91747e-19 $X=0.527 $Y=0.153 $X2=0.081 $Y2=0.135
cc_23 N_4_c_33_n N_D_c_99_n 2.1478e-19 $X=0.151 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_4_c_39_p N_D_c_101_n 2.3983e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_25 N_4_c_40_p N_D_c_102_n 8.99815e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_26 N_4_c_40_p N_D_c_103_n 8.75229e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_27 N_4_M3_g N_6_c_121_n 0.00355599f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_28 N_4_c_43_p N_6_c_121_n 0.00126153f $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.054
cc_29 N_4_M3_g N_6_M4_g 0.00355599f $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_4_M8_g N_6_M7_g 0.00355599f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_31 N_4_M8_g N_6_c_125_n 0.00355599f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_32 N_4_M8_g N_6_c_126_n 0.00250257f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_33 N_4_c_48_p N_6_c_126_n 0.00180656f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_34 N_4_c_49_p N_6_c_126_n 6.4075e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_35 N_4_c_37_p N_6_c_126_n 0.00187561f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_36 N_4_c_51_p N_6_c_126_n 0.00123876f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_34_n N_6_c_116_n 2.97444e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_31_n N_6_c_132_n 2.38327e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_34_n N_6_c_117_n 2.85146e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_40_p N_6_c_118_n 2.46239e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_41 N_4_c_31_n N_6_c_135_n 2.31165e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_42 N_4_c_39_p N_6_c_136_n 9.24693e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_43 N_4_c_37_p N_6_c_137_n 3.67557e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_44 N_4_c_37_p N_6_c_138_n 8.06691e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_45 N_4_c_37_p N_6_c_139_n 2.46239e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_46 N_4_c_40_p N_6_c_119_n 0.0299327f $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_39_p N_6_c_119_n 2.98936e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_48 N_4_c_37_p N_6_c_142_n 2.81476e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_49 N_4_c_40_p N_6_c_143_n 8.79704e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_50 N_4_c_34_n N_6_c_143_n 0.00524677f $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_51 N_4_c_37_p N_6_c_145_n 9.92294e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_52 N_4_c_39_p N_6_c_145_n 5.5596e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_53 N_4_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_54 N_4_c_69_p N_7_c_219_n 3.42573e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_55 N_4_c_69_p N_7_c_220_n 5.29207e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_56 N_4_c_51_p N_7_c_221_n 0.00318218f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_57 N_4_c_49_p N_7_c_222_n 0.00115177f $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_58 N_4_c_49_p N_7_c_223_n 3.42573e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_59 N_4_M8_g N_8_M6_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_60 N_4_c_48_p N_8_c_262_n 3.88499e-19 $X=0.675 $Y=0.135 $X2=0.081 $Y2=0.135
cc_61 N_4_c_69_p N_8_c_262_n 3.00379e-19 $X=0.601 $Y=0.153 $X2=0.081 $Y2=0.135
cc_62 N_4_c_39_p N_8_c_264_n 2.36208e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_63 N_4_M3_g N_8_c_265_n 3.49806e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_4_c_39_p N_8_c_265_n 3.83282e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_65 N_4_c_39_p N_8_c_267_n 7.25941e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_66 N_4_c_39_p N_8_c_268_n 7.25941e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_67 N_4_c_37_p N_8_c_269_n 0.00118282f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_68 N_4_c_39_p N_8_c_269_n 8.1935e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_69 N_4_c_37_p N_8_c_271_n 0.00132871f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_70 N_4_c_69_p N_8_c_272_n 0.00132871f $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_71 N_4_c_37_p N_8_c_273_n 2.54113e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_72 N_4_c_37_p N_8_c_274_n 3.92135e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_73 N_4_c_39_p N_8_c_275_n 7.25941e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_74 N_4_M8_g N_9_M9_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_75 N_4_c_49_p N_10_c_340_n 2.24654e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_76 N_4_c_49_p N_10_c_341_n 5.06919e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_77 N_4_M8_g N_10_c_342_n 3.47752e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_78 N_4_c_51_p N_10_c_342_n 5.72565e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_79 N_4_c_49_p N_10_c_344_n 2.46558e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_80 N_4_c_51_p N_10_c_345_n 0.00319993f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_81 N_4_c_49_p N_10_c_346_n 2.9112e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_82 N_4_c_37_p N_12_c_404_n 3.46326e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_83 N_D_M2_g N_6_c_121_n 0.00341068f $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_84 N_D_c_99_n N_6_c_121_n 0.00114686f $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_85 D N_6_c_149_n 0.00215667f $X=0.244 $Y=0.082 $X2=0.0505 $Y2=0.234
cc_86 N_D_c_103_n N_6_c_150_n 0.00215667f $X=0.243 $Y=0.135 $X2=0.405 $Y2=0.153
cc_87 N_D_c_103_n N_6_c_118_n 0.00225008f $X=0.243 $Y=0.135 $X2=0.175 $Y2=0.153
cc_88 N_D_c_109_p N_6_c_137_n 0.00127755f $X=0.281 $Y=0.135 $X2=0.151 $Y2=0.135
cc_89 N_D_c_99_n N_6_c_119_n 2.11668e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_90 N_D_c_103_n N_6_c_119_n 0.00122387f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_91 D N_6_c_120_n 0.00215667f $X=0.244 $Y=0.082 $X2=0.018 $Y2=0.153
cc_92 N_D_c_113_p N_6_c_143_n 0.00215667f $X=0.243 $Y=0.126 $X2=0 $Y2=0
cc_93 N_D_c_103_n N_6_c_145_n 0.00120973f $X=0.243 $Y=0.135 $X2=0.027 $Y2=0.153
cc_94 N_D_c_103_n N_8_c_276_n 2.80198e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_95 N_6_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_96 N_6_M7_g N_7_M5_g 2.13359e-19 $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_97 N_6_c_126_n N_7_M5_g 0.00205997f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_98 N_6_c_142_n N_7_M5_g 3.15189e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_99 N_6_c_126_n N_7_c_228_n 6.55731e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_100 N_6_c_126_n N_7_c_229_n 2.12581e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_101 N_6_c_126_n N_7_M19_s 2.50995e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_102 N_6_M7_g N_7_c_231_n 0.00200065f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_103 N_6_c_126_n N_7_c_231_n 0.00312129f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_104 N_6_c_126_n N_7_c_220_n 3.41745e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_105 N_6_M7_g N_7_c_221_n 3.41702e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_106 N_6_M7_g N_7_c_222_n 2.26424e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_107 N_6_c_142_n N_7_c_236_n 5.75704e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_108 N_6_c_171_p N_7_c_237_n 0.00195059f $X=0.621 $Y=0.178 $X2=0 $Y2=0
cc_109 N_6_c_126_n N_7_c_237_n 0.00191847f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_110 N_6_M7_g N_7_c_239_n 3.8308e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_111 N_6_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_112 N_6_M7_g N_8_M6_g 0.00341068f $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_113 N_6_c_126_n N_8_M6_g 0.00302156f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_114 N_6_c_119_n N_8_c_264_n 3.12535e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_115 N_6_c_145_n N_8_c_264_n 8.9852e-19 $X=0.324 $Y=0.167 $X2=0 $Y2=0
cc_116 N_6_c_119_n N_8_c_276_n 0.0015935f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_117 N_6_M4_g N_8_c_283_n 3.68551e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_118 N_6_M4_g N_8_c_284_n 2.06635e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_119 N_6_M4_g N_8_c_269_n 2.27069e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_120 N_6_c_183_p N_8_c_286_n 4.73369e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_121 N_6_c_142_n N_8_c_286_n 0.00174159f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_122 N_6_c_183_p N_8_c_288_n 0.00171407f $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_123 N_6_c_126_n N_8_c_288_n 5.88593e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_124 N_6_c_119_n N_8_c_288_n 0.00104904f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_125 N_6_c_188_p N_8_c_288_n 2.15173e-19 $X=0.324 $Y=0.178 $X2=0 $Y2=0
cc_126 N_6_c_126_n N_8_c_271_n 8.16411e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_127 N_6_c_126_n N_8_c_272_n 3.32592e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_128 N_6_c_142_n N_8_c_272_n 8.9822e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_129 N_6_c_126_n N_8_c_295_n 4.02972e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_130 N_6_c_125_n N_9_M9_g 0.00341068f $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_131 N_6_c_125_n N_10_M10_g 2.13359e-19 $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_132 N_6_c_126_n N_10_c_340_n 8.27829e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_133 N_6_c_126_n N_10_M20_s 3.37661e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_134 N_6_c_126_n N_10_c_350_n 0.00145548f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_135 N_6_c_125_n N_10_c_351_n 3.03386e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_136 N_6_c_125_n N_10_c_352_n 2.58526e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_137 N_6_c_125_n N_10_c_353_n 0.00228871f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_138 N_6_c_126_n N_10_c_353_n 7.89371e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_139 N_6_c_125_n N_10_c_355_n 4.55487e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_140 N_6_c_126_n N_10_c_356_n 4.54272e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_141 N_6_c_125_n N_10_c_357_n 5.68093e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_142 N_6_c_126_n N_10_c_357_n 2.2968e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_143 N_6_c_121_n N_12_c_404_n 0.00514294f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_144 N_6_c_137_n N_12_c_404_n 0.00114179f $X=0.333 $Y=0.135 $X2=0 $Y2=0
cc_145 N_6_c_126_n N_13_M17_s 2.36286e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.216
cc_146 N_6_M4_g N_13_c_411_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_147 N_6_c_183_p N_13_c_411_n 5.41258e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_148 N_6_c_126_n N_13_c_411_n 0.00230928f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_149 N_6_c_119_n N_13_c_411_n 7.09553e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_150 N_6_c_125_n N_14_c_420_n 0.00198387f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_151 N_6_c_126_n N_14_c_420_n 4.51352e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_152 N_6_c_139_n N_16_M15_s 8.59575e-19 $X=0.324 $Y=0.189 $X2=0.081 $Y2=0.054
cc_153 N_6_c_145_n N_16_M15_s 2.57402e-19 $X=0.324 $Y=0.167 $X2=0.081 $Y2=0.054
cc_154 N_6_c_188_p N_16_M15_s 2.18007e-19 $X=0.324 $Y=0.178 $X2=0.081 $Y2=0.054
cc_155 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_156 N_7_c_241_p N_8_M6_g 3.87418e-19 $X=0.576 $Y=0.09 $X2=0.135 $Y2=0.054
cc_157 N_7_c_221_n N_8_c_262_n 2.20449e-19 $X=0.621 $Y=0.122 $X2=0.135 $Y2=0.135
cc_158 N_7_c_243_p N_8_c_283_n 3.63506e-19 $X=0.594 $Y=0.054 $X2=0.018 $Y2=0.107
cc_159 N_7_c_244_p N_8_c_284_n 3.19692e-19 $X=0.513 $Y=0.09 $X2=0.018 $Y2=0.162
cc_160 N_7_c_241_p N_8_c_284_n 0.00114151f $X=0.576 $Y=0.09 $X2=0.018 $Y2=0.162
cc_161 N_7_c_246_p N_8_c_302_n 7.39815e-19 $X=0.621 $Y=0.14 $X2=0.027 $Y2=0.234
cc_162 N_7_c_241_p N_8_c_303_n 0.0047777f $X=0.576 $Y=0.09 $X2=0.054 $Y2=0.234
cc_163 N_7_M5_g N_8_c_272_n 3.12986e-19 $X=0.513 $Y=0.0405 $X2=0.047 $Y2=0.234
cc_164 N_7_c_244_p N_8_c_273_n 5.2508e-19 $X=0.513 $Y=0.09 $X2=0.033 $Y2=0.153
cc_165 N_7_c_228_n N_10_c_340_n 0.0027803f $X=0.594 $Y=0.0405 $X2=0.675
+ $Y2=0.135
cc_166 N_7_c_243_p N_10_c_340_n 3.72596e-19 $X=0.594 $Y=0.054 $X2=0.675
+ $Y2=0.135
cc_167 N_7_c_239_n N_10_c_340_n 3.30531e-19 $X=0.621 $Y=0.09 $X2=0.675 $Y2=0.135
cc_168 N_7_c_231_n N_10_c_350_n 0.00220898f $X=0.65 $Y=0.2295 $X2=0.056
+ $Y2=0.054
cc_169 N_7_c_228_n N_10_c_341_n 5.23227e-19 $X=0.594 $Y=0.0405 $X2=0 $Y2=0
cc_170 N_7_c_243_p N_10_c_364_n 2.3746e-19 $X=0.594 $Y=0.054 $X2=0.018 $Y2=0.107
cc_171 N_7_c_239_n N_10_c_351_n 4.46294e-19 $X=0.621 $Y=0.09 $X2=0.018 $Y2=0.162
cc_172 N_7_c_237_n N_10_c_353_n 4.46294e-19 $X=0.621 $Y=0.203 $X2=0.027
+ $Y2=0.036
cc_173 N_7_c_231_n N_10_c_356_n 3.64147e-19 $X=0.65 $Y=0.2295 $X2=0.405
+ $Y2=0.153
cc_174 N_7_c_220_n N_10_c_356_n 4.68959e-19 $X=0.612 $Y=0.234 $X2=0.405
+ $Y2=0.153
cc_175 N_7_c_260_p N_10_c_357_n 4.46294e-19 $X=0.621 $Y=0.101 $X2=0.675
+ $Y2=0.153
cc_176 N_8_c_264_n N_12_c_404_n 0.00119486f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_177 N_8_c_273_n N_12_c_404_n 0.00390673f $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_178 N_8_c_274_n N_12_c_404_n 5.36233e-19 $X=0.45 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_179 N_8_c_264_n N_13_c_411_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_180 N_8_c_310_p N_13_c_411_n 0.00209454f $X=0.45 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_181 N_8_c_311_p N_13_c_411_n 0.0013184f $X=0.434 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_182 N_8_c_312_p N_13_c_411_n 0.00119522f $X=0.459 $Y=0.225 $X2=0.405
+ $Y2=0.0675
cc_183 N_8_c_273_n N_13_c_411_n 5.72158e-19 $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_184 N_9_M9_g N_10_M10_g 0.00268443f $X=0.783 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_185 N_9_c_317_p N_10_M10_g 3.74489e-19 $X=0.846 $Y=0.036 $X2=0.135 $Y2=0.054
cc_186 N_9_c_318_p N_10_c_372_n 0.00141609f $X=0.792 $Y=0.036 $X2=0 $Y2=0
cc_187 N_9_c_319_p N_10_c_364_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.018
+ $Y2=0.107
cc_188 N_9_c_320_p N_10_c_351_n 3.34766e-19 $X=0.783 $Y=0.1055 $X2=0.018
+ $Y2=0.162
cc_189 N_9_c_319_p N_10_c_351_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.018
+ $Y2=0.162
cc_190 N_9_c_322_p N_10_c_353_n 2.41112e-19 $X=0.945 $Y=0.225 $X2=0.027
+ $Y2=0.036
cc_191 N_9_c_323_p N_10_c_377_n 2.6154e-19 $X=0.828 $Y=0.036 $X2=0.054 $Y2=0.036
cc_192 N_9_M9_g N_10_c_378_n 6.3699e-19 $X=0.783 $Y=0.0405 $X2=0.047 $Y2=0.036
cc_193 N_9_c_319_p N_10_c_378_n 9.10342e-19 $X=0.783 $Y=0.105 $X2=0.047
+ $Y2=0.036
cc_194 N_9_c_317_p N_10_c_380_n 4.40983e-19 $X=0.846 $Y=0.036 $X2=0.027
+ $Y2=0.234
cc_195 N_9_c_327_p N_10_c_381_n 5.13693e-19 $X=0.882 $Y=0.036 $X2=0.033
+ $Y2=0.153
cc_196 N_9_c_328_p N_10_c_382_n 0.00149072f $X=0.9 $Y=0.234 $X2=0.033 $Y2=0.153
cc_197 N_9_c_329_p N_10_c_383_n 4.52584e-19 $X=0.9 $Y=0.036 $X2=0.601 $Y2=0.153
cc_198 N_9_c_330_p N_10_c_383_n 0.00299476f $X=0.945 $Y=0.167 $X2=0.601
+ $Y2=0.153
cc_199 N_9_c_331_p N_10_c_346_n 2.40515e-19 $X=0.936 $Y=0.036 $X2=0 $Y2=0
cc_200 N_9_c_332_p N_10_c_346_n 7.44774e-19 $X=0.918 $Y=0.234 $X2=0 $Y2=0
cc_201 N_9_c_330_p N_10_c_346_n 9.28741e-19 $X=0.945 $Y=0.167 $X2=0 $Y2=0
cc_202 N_9_c_334_p N_10_c_388_n 0.00322692f $X=0.945 $Y=0.117 $X2=0 $Y2=0
cc_203 N_9_c_335_p N_QN_c_397_n 3.5495e-19 $X=0.945 $Y=0.171 $X2=0.405 $Y2=0.135
cc_204 N_9_c_336_p N_QN_c_398_n 3.5495e-19 $X=0.945 $Y=0.09 $X2=0.405 $Y2=0.2295
cc_205 N_9_c_331_p N_QN_c_399_n 4.40179e-19 $X=0.936 $Y=0.036 $X2=0.675
+ $Y2=0.2295
cc_206 N_9_c_338_p N_QN_c_400_n 4.34861e-19 $X=0.936 $Y=0.234 $X2=0.071
+ $Y2=0.216
cc_207 N_9_c_318_p N_14_c_420_n 7.33799e-19 $X=0.792 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_208 N_10_c_346_n N_QN_c_401_n 2.28166e-19 $X=0.999 $Y=0.153 $X2=0 $Y2=0
cc_209 N_10_c_388_n N_QN_c_401_n 0.00331683f $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_210 N_10_c_388_n N_QN_c_403_n 5.42522e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_211 N_10_c_340_n N_14_c_420_n 0.00182708f $X=0.648 $Y=0.0405 $X2=0.405
+ $Y2=0.0675
cc_212 N_10_c_372_n N_14_c_420_n 0.0020512f $X=0.72 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_213 N_10_c_394_p N_14_c_420_n 0.00131745f $X=0.704 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_214 N_10_c_364_n N_14_c_420_n 0.00103589f $X=0.729 $Y=0.081 $X2=0.405
+ $Y2=0.0675
cc_215 N_10_c_355_n N_14_c_420_n 4.02739e-19 $X=0.774 $Y=0.162 $X2=0.405
+ $Y2=0.0675

* END of "./DFFHQNx1_ASAP7_75t_SRAM.pex.sp.DFFHQNX1_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DFFHQNx2_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:24:31 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DFFHQNx2_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DFFHQNx2_ASAP7_75t_SRAM.pex.sp.pex"
* File: DFFHQNx2_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:24:31 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%CLK 2 5 7 12 14 VSS
c20 14 VSS 0.00674559f $X=0.081 $Y=0.135
c21 12 VSS 0.00682604f $X=0.082 $Y=0.119
c22 5 VSS 0.00206449f $X=0.081 $Y=0.135
c23 2 VSS 0.0629f $X=0.081 $Y=0.054
r24 12 14 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.135
r25 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r26 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r27 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%4 2 7 10 13 15 18 21 23 25 28 30 36 37 38 41 42
+ 45 52 59 67 68 70 72 73 78 79 83 88 VSS
c77 114 VSS 1.06551e-19 $X=0.03 $Y=0.153
c78 113 VSS 6.89947e-19 $X=0.027 $Y=0.153
c79 88 VSS 0.00102973f $X=0.675 $Y=0.135
c80 83 VSS 8.66895e-19 $X=0.405 $Y=0.135
c81 79 VSS 0.00121012f $X=0.151 $Y=0.135
c82 78 VSS 0.00390107f $X=0.151 $Y=0.135
c83 73 VSS 0.00263053f $X=0.601 $Y=0.153
c84 72 VSS 0.00556612f $X=0.527 $Y=0.153
c85 70 VSS 0.00405122f $X=0.675 $Y=0.153
c86 68 VSS 0.00330975f $X=0.29 $Y=0.153
c87 67 VSS 0.00602706f $X=0.175 $Y=0.153
c88 59 VSS 6.74716e-19 $X=0.033 $Y=0.153
c89 55 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c90 54 VSS 0.00180216f $X=0.047 $Y=0.234
c91 52 VSS 0.00250119f $X=0.054 $Y=0.234
c92 50 VSS 0.00305101f $X=0.027 $Y=0.234
c93 48 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c94 47 VSS 0.00199699f $X=0.047 $Y=0.036
c95 45 VSS 0.00250119f $X=0.054 $Y=0.036
c96 43 VSS 0.00305101f $X=0.027 $Y=0.036
c97 42 VSS 4.88707e-19 $X=0.018 $Y=0.2125
c98 41 VSS 0.00180713f $X=0.018 $Y=0.2
c99 40 VSS 4.69158e-19 $X=0.018 $Y=0.225
c100 38 VSS 0.00173342f $X=0.018 $Y=0.107
c101 37 VSS 9.57865e-19 $X=0.018 $Y=0.07
c102 36 VSS 0.00172854f $X=0.018 $Y=0.144
c103 33 VSS 0.00509483f $X=0.056 $Y=0.216
c104 30 VSS 2.98509e-19 $X=0.071 $Y=0.216
c105 28 VSS 0.00497933f $X=0.056 $Y=0.054
c106 25 VSS 2.98509e-19 $X=0.071 $Y=0.054
c107 21 VSS 0.00214819f $X=0.675 $Y=0.135
c108 18 VSS 0.0585656f $X=0.675 $Y=0.0405
c109 13 VSS 0.00214124f $X=0.405 $Y=0.135
c110 10 VSS 0.058827f $X=0.405 $Y=0.0675
c111 2 VSS 0.0628024f $X=0.135 $Y=0.054
r112 113 114 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r113 110 113 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r114 78 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.151 $Y=0.135 $X2=0.151
+ $Y2=0.135
r115 72 73 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.601 $Y2=0.153
r116 70 73 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.675
+ $Y=0.153 $X2=0.601 $Y2=0.153
r117 70 88 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.675 $Y=0.153 $X2=0.675
+ $Y2=0.153
r118 67 68 7.80864 $w=1.8e-08 $l=1.15e-07 $layer=M2 $thickness=3.6e-08 $X=0.175
+ $Y=0.153 $X2=0.29 $Y2=0.153
r119 65 72 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.527 $Y2=0.153
r120 65 68 7.80864 $w=1.8e-08 $l=1.15e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.29 $Y2=0.153
r121 65 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r122 62 67 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.151
+ $Y=0.153 $X2=0.175 $Y2=0.153
r123 62 79 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.151 $Y=0.153 $X2=0.151
+ $Y2=0.153
r124 59 114 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r125 58 62 8.01235 $w=1.8e-08 $l=1.18e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.151 $Y2=0.153
r126 58 59 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r127 54 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r128 52 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r129 50 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r130 47 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r131 45 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r132 43 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r133 41 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r134 40 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r135 40 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r136 39 110 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r137 39 41 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.2
r138 37 38 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.107
r139 36 110 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r140 36 38 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.107
r141 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r142 35 37 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r143 33 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r144 30 33 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r145 28 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r146 25 28 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r147 21 88 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.135 $X2=0.675
+ $Y2=0.135
r148 21 23 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2295
r149 18 21 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.135
r150 13 83 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r151 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2295
r152 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r153 5 78 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.151 $Y2=0.135
r154 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r155 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%D 2 5 7 10 12 14 21 23 28 VSS
c18 28 VSS 0.00931225f $X=0.243 $Y=0.135
c19 24 VSS 2.45662e-20 $X=0.276 $Y=0.135
c20 23 VSS 0.00111822f $X=0.271 $Y=0.135
c21 21 VSS 2.56376e-19 $X=0.281 $Y=0.135
c22 14 VSS 2.7811e-19 $X=0.243 $Y=0.116
c23 12 VSS 0.00925957f $X=0.244 $Y=0.082
c24 10 VSS 2.38113e-19 $X=0.243 $Y=0.126
c25 5 VSS 0.00522238f $X=0.297 $Y=0.135
c26 2 VSS 0.0630392f $X=0.297 $Y=0.0675
r27 23 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.271
+ $Y=0.135 $X2=0.276 $Y2=0.135
r28 21 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.281
+ $Y=0.135 $X2=0.276 $Y2=0.135
r29 21 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.281 $Y=0.135 $X2=0.281
+ $Y2=0.135
r30 19 28 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.243 $Y2=0.135
r31 19 23 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.271 $Y2=0.135
r32 13 14 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.106 $X2=0.243 $Y2=0.116
r33 12 13 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.082 $X2=0.243 $Y2=0.106
r34 10 28 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.135
r35 10 14 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.116
r36 5 22 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.281 $Y2=0.135
r37 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r38 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%6 2 5 8 14 17 20 23 28 35 39 44 50 55 57 61 66
+ 67 68 75 77 78 87 89 105 110 111 113 114 VSS
c102 114 VSS 2.23151e-19 $X=0.324 $Y=0.178
c103 113 VSS 4.08645e-19 $X=0.324 $Y=0.167
c104 111 VSS 7.77947e-19 $X=0.189 $Y=0.167
c105 110 VSS 9.60988e-19 $X=0.189 $Y=0.106
c106 105 VSS 6.81413e-19 $X=0.513 $Y=0.18
c107 89 VSS 0.0113851f $X=0.513 $Y=0.189
c108 87 VSS 0.00141172f $X=0.324 $Y=0.189
c109 78 VSS 4.01771e-19 $X=0.342 $Y=0.135
c110 77 VSS 5.28662e-19 $X=0.333 $Y=0.135
c111 75 VSS 7.4105e-19 $X=0.351 $Y=0.135
c112 68 VSS 0.00169555f $X=0.18 $Y=0.234
c113 67 VSS 9.43175e-19 $X=0.189 $Y=0.225
c114 66 VSS 0.00196236f $X=0.189 $Y=0.234
c115 61 VSS 0.00196921f $X=0.162 $Y=0.234
c116 57 VSS 0.00170883f $X=0.18 $Y=0.036
c117 55 VSS 0.00196236f $X=0.189 $Y=0.036
c118 50 VSS 0.00193426f $X=0.162 $Y=0.036
c119 47 VSS 0.00715944f $X=0.16 $Y=0.216
c120 42 VSS 0.00719538f $X=0.16 $Y=0.054
c121 35 VSS 0.0611368f $X=0.725 $Y=0.178
c122 28 VSS 0.00126548f $X=0.464 $Y=0.178
c123 20 VSS 0.0618767f $X=0.729 $Y=0.178
c124 17 VSS 1.08457e-19 $X=0.621 $Y=0.178
c125 14 VSS 0.0600454f $X=0.621 $Y=0.0405
c126 8 VSS 0.0602427f $X=0.459 $Y=0.0405
c127 2 VSS 0.0623279f $X=0.351 $Y=0.135
r128 113 114 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.324 $Y=0.167 $X2=0.324 $Y2=0.178
r129 110 111 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.106 $X2=0.189 $Y2=0.167
r130 104 105 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r131 89 105 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r132 87 114 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.189 $X2=0.324 $Y2=0.178
r133 86 89 12.8333 $w=1.8e-08 $l=1.89e-07 $layer=M2 $thickness=3.6e-08 $X=0.324
+ $Y=0.189 $X2=0.513 $Y2=0.189
r134 86 87 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.324 $Y=0.189 $X2=0.324
+ $Y2=0.189
r135 83 111 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.167
r136 82 86 9.16667 $w=1.8e-08 $l=1.35e-07 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.324 $Y2=0.189
r137 82 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.189 $X2=0.189
+ $Y2=0.189
r138 77 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.135 $X2=0.342 $Y2=0.135
r139 75 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.342 $Y2=0.135
r140 72 113 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.144 $X2=0.324 $Y2=0.167
r141 71 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.135 $X2=0.333 $Y2=0.135
r142 71 72 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.135 $X2=0.324 $Y2=0.144
r143 68 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r144 67 83 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.189
r145 66 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r146 66 67 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.189 $Y2=0.225
r147 61 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r148 57 58 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r149 56 110 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.106
r150 55 58 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r151 55 56 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r152 50 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r153 47 61 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r154 44 47 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r155 42 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r156 39 42 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r157 28 104 39.0385 $w=2.6e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.178 $X2=0.513 $Y2=0.178
r158 20 35 3.07692 $w=2.6e-08 $l=4e-09 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.178 $X2=0.725 $Y2=0.178
r159 20 23 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.178 $X2=0.729 $Y2=0.2295
r160 17 35 82.8571 $w=2.6e-08 $l=1.04e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.725 $Y2=0.178
r161 17 104 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.513 $Y2=0.178
r162 14 17 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0405 $X2=0.621 $Y2=0.178
r163 11 28 3.84615 $w=2.6e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.178 $X2=0.464 $Y2=0.178
r164 8 11 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.178
r165 2 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r166 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%7 2 5 7 9 10 13 14 17 19 22 29 30 31 38 43 44 45
+ 46 47 48 52 53 VSS
c43 54 VSS 3.52511e-19 $X=0.612 $Y=0.09
c44 53 VSS 1.80704e-19 $X=0.603 $Y=0.09
c45 52 VSS 5.96246e-19 $X=0.621 $Y=0.09
c46 49 VSS 6.86664e-19 $X=0.621 $Y=0.224
c47 48 VSS 4.95788e-19 $X=0.621 $Y=0.203
c48 47 VSS 1.19762e-19 $X=0.621 $Y=0.167
c49 46 VSS 3.19764e-19 $X=0.621 $Y=0.165
c50 45 VSS 3.13056e-19 $X=0.621 $Y=0.14
c51 44 VSS 3.62783e-19 $X=0.621 $Y=0.122
c52 43 VSS 1.48552e-19 $X=0.621 $Y=0.101
c53 38 VSS 0.00113884f $X=0.594 $Y=0.054
c54 31 VSS 0.00668633f $X=0.612 $Y=0.234
c55 30 VSS 3.5821e-19 $X=0.5805 $Y=0.09
c56 29 VSS 0.00257846f $X=0.576 $Y=0.09
c57 24 VSS 1.48201e-19 $X=0.585 $Y=0.09
c58 22 VSS 0.0179338f $X=0.65 $Y=0.2295
c59 19 VSS 3.14771e-19 $X=0.665 $Y=0.2295
c60 17 VSS 2.67274e-19 $X=0.592 $Y=0.2295
c61 13 VSS 0.0252201f $X=0.594 $Y=0.0405
c62 9 VSS 6.29543e-19 $X=0.611 $Y=0.0405
c63 5 VSS 0.00238279f $X=0.513 $Y=0.09
c64 2 VSS 0.0584396f $X=0.513 $Y=0.0405
r65 53 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.603
+ $Y=0.09 $X2=0.612 $Y2=0.09
r66 52 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.612 $Y2=0.09
r67 51 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.09 $X2=0.603 $Y2=0.09
r68 49 50 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.224 $X2=0.621 $Y2=0.2245
r69 48 49 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.224
r70 47 48 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.203
r71 46 47 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.167
r72 45 46 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r73 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r74 43 44 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.101 $X2=0.621 $Y2=0.122
r75 42 50 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.2245
r76 41 52 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.09
r77 41 43 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.101
r78 36 51 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.09
r79 36 38 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.054
r80 31 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r81 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r82 29 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.09 $X2=0.5805 $Y2=0.09
r83 26 29 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.09 $X2=0.576 $Y2=0.09
r84 24 51 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.594 $Y2=0.09
r85 24 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.5805 $Y2=0.09
r86 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2295 $X2=0.65 $Y2=0.2295
r87 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.592
+ $Y=0.2295 $X2=0.65 $Y2=0.2295
r88 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r89 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r90 13 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.054 $X2=0.594
+ $Y2=0.054
r91 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.594 $Y2=0.0405
r92 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0405 $X2=0.594 $Y2=0.0405
r93 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.09 $X2=0.513
+ $Y2=0.09
r94 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.09 $X2=0.513 $Y2=0.2295
r95 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.09
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%8 2 5 7 9 14 17 21 22 25 27 33 35 37 38 39 41 43
+ 44 45 46 50 52 53 54 55 59 62 65 VSS
c53 65 VSS 2.85958e-19 $X=0.459 $Y=0.131
c54 62 VSS 0.00341346f $X=0.45 $Y=0.036
c55 61 VSS 0.0025252f $X=0.459 $Y=0.036
c56 59 VSS 0.00276391f $X=0.432 $Y=0.036
c57 55 VSS 4.23521e-19 $X=0.5445 $Y=0.131
c58 54 VSS 3.49205e-20 $X=0.522 $Y=0.131
c59 53 VSS 2.00095e-19 $X=0.504 $Y=0.131
c60 52 VSS 0.00133241f $X=0.496 $Y=0.131
c61 50 VSS 2.94642e-19 $X=0.567 $Y=0.131
c62 47 VSS 4.32029e-19 $X=0.459 $Y=0.214
c63 46 VSS 2.06877e-19 $X=0.459 $Y=0.203
c64 45 VSS 6.09344e-21 $X=0.459 $Y=0.167
c65 44 VSS 2.12612e-19 $X=0.459 $Y=0.165
c66 43 VSS 2.51143e-19 $X=0.459 $Y=0.225
c67 41 VSS 3.68971e-19 $X=0.459 $Y=0.114
c68 40 VSS 3.4692e-19 $X=0.459 $Y=0.106
c69 38 VSS 7.88894e-19 $X=0.459 $Y=0.081
c70 37 VSS 2.0833e-19 $X=0.459 $Y=0.122
c71 35 VSS 0.00142907f $X=0.434 $Y=0.234
c72 34 VSS 3.2912e-19 $X=0.418 $Y=0.234
c73 33 VSS 0.00146362f $X=0.414 $Y=0.234
c74 32 VSS 0.00227054f $X=0.396 $Y=0.234
c75 27 VSS 0.00148441f $X=0.378 $Y=0.234
c76 25 VSS 0.00389542f $X=0.45 $Y=0.234
c77 24 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c78 21 VSS 0.00379676f $X=0.378 $Y=0.2025
c79 18 VSS 1.15515e-19 $X=0.3735 $Y=0.216
c80 16 VSS 5.70081e-19 $X=0.432 $Y=0.0405
c81 10 VSS 7.61325e-20 $X=0.4275 $Y=0.054
c82 5 VSS 0.0022736f $X=0.567 $Y=0.1305
c83 2 VSS 0.0591678f $X=0.567 $Y=0.0405
r84 62 63 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r85 61 63 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r86 58 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r87 58 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r88 54 55 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r89 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r90 52 53 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.496
+ $Y=0.131 $X2=0.504 $Y2=0.131
r91 50 55 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r92 48 65 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r93 48 52 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.496 $Y2=0.131
r94 46 47 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.203 $X2=0.459 $Y2=0.214
r95 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.167 $X2=0.459 $Y2=0.203
r96 44 45 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.167
r97 43 47 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r98 42 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r99 42 44 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.165
r100 40 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.106 $X2=0.459 $Y2=0.114
r101 39 40 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.099 $X2=0.459 $Y2=0.106
r102 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.099
r103 37 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r104 37 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.114
r105 36 61 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r106 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.081
r107 34 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.234 $X2=0.434 $Y2=0.234
r108 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.418 $Y2=0.234
r109 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r110 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r111 25 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r112 25 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.434 $Y2=0.234
r113 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r114 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r115 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r116 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r117 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r118 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r119 13 59 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r120 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r121 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r122 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r123 5 50 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.131 $X2=0.567
+ $Y2=0.131
r124 5 7 370.904 $w=2e-08 $l=9.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1305 $X2=0.567 $Y2=0.2295
r125 2 5 337.185 $w=2e-08 $l=9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.1305
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%9 2 5 7 9 14 21 25 26 30 31 32 33 39 40 42 45 46
+ 48 VSS
c24 48 VSS 0.0023571f $X=0.945 $Y=0.216
c25 47 VSS 1.87203e-19 $X=0.945 $Y=0.171
c26 46 VSS 0.00102475f $X=0.945 $Y=0.167
c27 45 VSS 8.67706e-19 $X=0.945 $Y=0.117
c28 44 VSS 0.00182154f $X=0.945 $Y=0.09
c29 43 VSS 4.18448e-19 $X=0.945 $Y=0.054
c30 42 VSS 4.22172e-19 $X=0.945 $Y=0.225
c31 40 VSS 0.0018377f $X=0.918 $Y=0.234
c32 39 VSS 0.00568507f $X=0.9 $Y=0.234
c33 34 VSS 0.00474105f $X=0.936 $Y=0.234
c34 33 VSS 0.00189638f $X=0.9 $Y=0.036
c35 32 VSS 0.0035379f $X=0.882 $Y=0.036
c36 31 VSS 0.00146362f $X=0.846 $Y=0.036
c37 30 VSS 0.00510392f $X=0.828 $Y=0.036
c38 26 VSS 0.00226308f $X=0.792 $Y=0.036
c39 25 VSS 0.00668817f $X=0.936 $Y=0.036
c40 21 VSS 0.00122443f $X=0.783 $Y=0.105
c41 17 VSS 0.00481511f $X=0.862 $Y=0.2295
c42 12 VSS 0.00513464f $X=0.862 $Y=0.0405
c43 5 VSS 0.00277722f $X=0.783 $Y=0.1055
c44 2 VSS 0.0590816f $X=0.783 $Y=0.0405
r45 47 48 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.216
r46 46 47 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.167 $X2=0.945 $Y2=0.171
r47 45 46 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.117 $X2=0.945 $Y2=0.167
r48 44 45 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.09 $X2=0.945 $Y2=0.117
r49 43 44 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.054 $X2=0.945 $Y2=0.09
r50 42 48 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.216
r51 41 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.054
r52 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.234 $X2=0.918 $Y2=0.234
r53 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.9 $Y2=0.234
r54 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r55 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.918 $Y2=0.234
r56 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r57 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.846 $Y2=0.036
r58 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r59 28 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.846 $Y2=0.036
r60 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.036 $X2=0.828 $Y2=0.036
r61 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r62 25 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.9 $Y2=0.036
r63 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.783 $Y=0.045 $X2=0.792 $Y2=0.036
r64 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.105
r65 17 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234 $X2=0.864
+ $Y2=0.234
r66 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2295 $X2=0.862 $Y2=0.2295
r67 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036 $X2=0.864
+ $Y2=0.036
r68 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.862 $Y2=0.0405
r69 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.105 $X2=0.783
+ $Y2=0.105
r70 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.1055 $X2=0.783 $Y2=0.2295
r71 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.1055
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%10 2 7 10 15 18 21 23 25 26 29 30 31 34 35 40 41
+ 43 45 46 47 48 49 51 52 54 55 58 65 66 74 77 81 84 92 VSS
c65 92 VSS 0.00214204f $X=0.999 $Y=0.136
c66 84 VSS 0.00791777f $X=0.999 $Y=0.153
c67 81 VSS 0.00149602f $X=0.891 $Y=0.153
c68 78 VSS 4.17512e-19 $X=0.837 $Y=0.162
c69 77 VSS 1.52743e-19 $X=0.729 $Y=0.162
c70 74 VSS 0.00357121f $X=0.72 $Y=0.233
c71 73 VSS 0.00257308f $X=0.729 $Y=0.233
c72 66 VSS 4.30636e-19 $X=0.866 $Y=0.162
c73 65 VSS 1.23291e-19 $X=0.85 $Y=0.162
c74 63 VSS 2.75449e-19 $X=0.882 $Y=0.162
c75 58 VSS 3.94906e-19 $X=0.837 $Y=0.135
c76 55 VSS 3.26354e-19 $X=0.792 $Y=0.162
c77 54 VSS 0.00206921f $X=0.774 $Y=0.162
c78 52 VSS 0.00191548f $X=0.828 $Y=0.162
c79 51 VSS 0.00132112f $X=0.729 $Y=0.224
c80 49 VSS 1.52884e-19 $X=0.729 $Y=0.136
c81 48 VSS 2.77769e-19 $X=0.729 $Y=0.119
c82 47 VSS 1.41609e-19 $X=0.729 $Y=0.101
c83 46 VSS 3.52175e-19 $X=0.729 $Y=0.081
c84 45 VSS 2.73935e-19 $X=0.729 $Y=0.153
c85 43 VSS 0.00166757f $X=0.704 $Y=0.036
c86 42 VSS 4.5779e-19 $X=0.688 $Y=0.036
c87 41 VSS 0.00146362f $X=0.684 $Y=0.036
c88 40 VSS 0.00375563f $X=0.666 $Y=0.036
c89 35 VSS 0.00409736f $X=0.72 $Y=0.036
c90 34 VSS 0.00133398f $X=0.702 $Y=0.2295
c91 30 VSS 6.50675e-19 $X=0.719 $Y=0.2295
c92 29 VSS 0.0376609f $X=0.648 $Y=0.0405
c93 25 VSS 5.63046e-19 $X=0.665 $Y=0.0405
c94 21 VSS 0.00490443f $X=1.053 $Y=0.136
c95 18 VSS 0.0617781f $X=1.053 $Y=0.0675
c96 10 VSS 0.0612321f $X=0.999 $Y=0.0675
c97 5 VSS 0.00239735f $X=0.837 $Y=0.135
c98 2 VSS 0.0618222f $X=0.837 $Y=0.0405
r99 84 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.999 $Y=0.153 $X2=0.999
+ $Y2=0.153
r100 80 84 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.999 $Y2=0.153
r101 80 81 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r102 74 75 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.233 $X2=0.7245 $Y2=0.233
r103 73 75 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.233 $X2=0.7245 $Y2=0.233
r104 70 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.233 $X2=0.72 $Y2=0.233
r105 65 66 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.85
+ $Y=0.162 $X2=0.866 $Y2=0.162
r106 64 78 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.837 $Y2=0.162
r107 64 65 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.85 $Y2=0.162
r108 63 81 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.891 $Y2=0.162
r109 63 66 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.866 $Y2=0.162
r110 56 78 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.162
r111 56 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.135
r112 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.162 $X2=0.792 $Y2=0.162
r113 53 77 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.729 $Y2=0.162
r114 53 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.774 $Y2=0.162
r115 52 78 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.837 $Y2=0.162
r116 52 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.792 $Y2=0.162
r117 51 73 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.224 $X2=0.729 $Y2=0.233
r118 50 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.162
r119 50 51 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.224
r120 48 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.119 $X2=0.729 $Y2=0.136
r121 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.101 $X2=0.729 $Y2=0.119
r122 46 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.081 $X2=0.729 $Y2=0.101
r123 45 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.162
r124 45 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.136
r125 44 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.045 $X2=0.729 $Y2=0.081
r126 42 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.036 $X2=0.704 $Y2=0.036
r127 41 42 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.688 $Y2=0.036
r128 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.684 $Y2=0.036
r129 37 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.666 $Y2=0.036
r130 35 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.036 $X2=0.729 $Y2=0.045
r131 35 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.704 $Y2=0.036
r132 34 70 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.233
+ $X2=0.702 $Y2=0.233
r133 31 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2295 $X2=0.702 $Y2=0.2295
r134 30 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2295 $X2=0.702 $Y2=0.2295
r135 29 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r136 26 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0405 $X2=0.648 $Y2=0.0405
r137 25 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r138 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.136 $X2=1.053 $Y2=0.2025
r139 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.0675 $X2=1.053 $Y2=0.136
r140 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.999
+ $Y=0.136 $X2=1.053 $Y2=0.136
r141 13 92 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.136 $X2=0.999
+ $Y2=0.136
r142 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.136 $X2=0.999 $Y2=0.2025
r143 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.136
r144 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.135 $X2=0.837
+ $Y2=0.135
r145 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.2295
r146 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.0405 $X2=0.837 $Y2=0.135
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%QN 1 2 6 7 10 11 14 16 22 26 VSS
c13 26 VSS 0.00433723f $X=1.108 $Y=0.167
c14 25 VSS 0.00211706f $X=1.108 $Y=0.09
c15 24 VSS 0.00299339f $X=1.108 $Y=0.216
c16 16 VSS 0.0118434f $X=1.099 $Y=0.225
c17 14 VSS 0.00742878f $X=1.026 $Y=0.045
c18 11 VSS 0.0118436f $X=1.099 $Y=0.045
c19 10 VSS 0.00718893f $X=1.026 $Y=0.2025
c20 6 VSS 6.63935e-19 $X=1.043 $Y=0.2025
c21 1 VSS 6.63935e-19 $X=1.043 $Y=0.0675
r22 25 26 5.22839 $w=1.8e-08 $l=7.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.108
+ $Y=0.09 $X2=1.108 $Y2=0.167
r23 24 26 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.108
+ $Y=0.216 $X2=1.108 $Y2=0.167
r24 23 25 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.108
+ $Y=0.054 $X2=1.108 $Y2=0.09
r25 18 22 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.225 $X2=1.085 $Y2=0.225
r26 16 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.099 $Y=0.225 $X2=1.108 $Y2=0.216
r27 16 22 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.099
+ $Y=0.225 $X2=1.085 $Y2=0.225
r28 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.045 $X2=1.026
+ $Y2=0.045
r29 11 23 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.099 $Y=0.045 $X2=1.108 $Y2=0.054
r30 11 13 4.95679 $w=1.8e-08 $l=7.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.099
+ $Y=0.045 $X2=1.026 $Y2=0.045
r31 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.225 $X2=1.026
+ $Y2=0.225
r32 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.2025 $X2=1.026 $Y2=0.2025
r33 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.043 $Y=0.2025 $X2=1.026 $Y2=0.2025
r34 5 14 19.4196 $w=2.4e-08 $l=2.25e-08 $layer=LISD $thickness=2.8e-08 $X=1.026
+ $Y=0.0675 $X2=1.026 $Y2=0.045
r35 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.009
+ $Y=0.0675 $X2=1.026 $Y2=0.0675
r36 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.043
+ $Y=0.0675 $X2=1.026 $Y2=0.0675
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%12 1 6 9 VSS
c6 9 VSS 0.0270172f $X=0.38 $Y=0.0675
c7 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c8 4 VSS 3.25039e-19 $X=0.322 $Y=0.0675
r9 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r10 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%13 1 6 9 VSS
c10 9 VSS 0.0209308f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.6182e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%14 1 6 9 VSS
c8 9 VSS 0.0191671f $X=0.758 $Y=0.0405
c9 6 VSS 3.14771e-19 $X=0.773 $Y=0.0405
c10 4 VSS 2.6194e-19 $X=0.7 $Y=0.0405
r11 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r12 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.7
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r13 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.685
+ $Y=0.0405 $X2=0.7 $Y2=0.0405
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%15 1 2 VSS
c0 1 VSS 0.00225696f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%16 1 2 VSS
c3 1 VSS 0.00231486f $X=0.341 $Y=0.2025
r4 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends

.subckt PM_DFFHQNX2_ASAP7_75T_SRAM%17 1 2 VSS
c0 1 VSS 0.00219822f $X=0.773 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2295 $X2=0.739 $Y2=0.2295
.ends


* END of "./DFFHQNx2_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DFFHQNx2_ASAP7_75t_SRAM  VSS VDD CLK D QN
* 
* QN	QN
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_12_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_4_M3_g N_12_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_15_M4_d N_6_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_15_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_10_M7_d N_6_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.611
+ $Y=0.027
M8 N_14_M8_d N_4_M8_g N_10_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M9 VSS N_9_M9_g N_14_M9_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_9_M10_d N_10_M10_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.027
M11 N_QN_M11_d N_10_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M12 N_QN_M12_d N_10_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.027
M13 VDD N_CLK_M13_g N_4_M13_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M14 N_6_M14_d N_4_M14_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M15 N_16_M15_d N_D_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M16 N_8_M16_d N_6_M16_g N_16_M16_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M17 N_13_M17_d N_4_M17_g N_8_M17_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M18 VDD N_7_M18_g N_13_M18_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M19 N_7_M19_d N_8_M19_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M20 N_10_M20_d N_4_M20_g N_7_M20_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.665 $Y=0.216
M21 N_17_M21_d N_6_M21_g N_10_M21_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.719 $Y=0.216
M22 VDD N_9_M22_g N_17_M22_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M23 N_9_M23_d N_10_M23_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.216
M24 N_QN_M24_d N_10_M24_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
M25 N_QN_M25_d N_10_M25_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.162
*
* 
* .include "DFFHQNx2_ASAP7_75t_SRAM.pex.sp.DFFHQNX2_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DFFHQNx2_ASAP7_75t_SRAM.pex.sp.DFFHQNX2_ASAP7_75T_SRAM.pxi"
* File: DFFHQNx2_ASAP7_75t_SRAM.pex.sp.DFFHQNX2_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:24:31 2017
* 
x_PM_DFFHQNX2_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_13_p N_CLK_M13_g CLK
+ N_CLK_c_6_p VSS PM_DFFHQNX2_ASAP7_75T_SRAM%CLK
x_PM_DFFHQNX2_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M14_g N_4_M3_g N_4_c_43_p N_4_M17_g
+ N_4_M8_g N_4_c_48_p N_4_M20_g N_4_M0_s N_4_c_22_n N_4_M13_s N_4_c_23_n
+ N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_28_n N_4_c_29_n N_4_c_30_n
+ N_4_c_31_n N_4_c_40_p N_4_c_49_p N_4_c_37_p N_4_c_69_p N_4_c_33_n N_4_c_34_n
+ N_4_c_39_p N_4_c_51_p VSS PM_DFFHQNX2_ASAP7_75T_SRAM%4
x_PM_DFFHQNX2_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_99_n N_D_M15_g N_D_c_113_p D
+ N_D_c_101_n N_D_c_109_p N_D_c_102_n N_D_c_103_n VSS PM_DFFHQNX2_ASAP7_75T_SRAM%D
x_PM_DFFHQNX2_ASAP7_75T_SRAM%6 N_6_c_121_n N_6_M16_g N_6_M4_g N_6_M7_g N_6_c_171_p
+ N_6_c_125_n N_6_M21_g N_6_c_183_p N_6_c_126_n N_6_M1_d N_6_M14_d N_6_c_116_n
+ N_6_c_149_n N_6_c_132_n N_6_c_117_n N_6_c_150_n N_6_c_118_n N_6_c_135_n
+ N_6_c_136_n N_6_c_137_n N_6_c_138_n N_6_c_139_n N_6_c_119_n N_6_c_142_n
+ N_6_c_120_n N_6_c_143_n N_6_c_145_n N_6_c_188_p VSS PM_DFFHQNX2_ASAP7_75T_SRAM%6
x_PM_DFFHQNX2_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_244_p N_7_M18_g N_7_M7_s N_7_M6_d
+ N_7_c_228_n N_7_M19_d N_7_c_229_n N_7_M20_s N_7_c_231_n N_7_c_241_p
+ N_7_c_219_n N_7_c_220_n N_7_c_243_p N_7_c_260_p N_7_c_221_n N_7_c_246_p
+ N_7_c_222_n N_7_c_236_n N_7_c_237_n N_7_c_239_n N_7_c_223_n VSS
+ PM_DFFHQNX2_ASAP7_75T_SRAM%7
x_PM_DFFHQNX2_ASAP7_75T_SRAM%8 N_8_M6_g N_8_c_262_n N_8_M19_g N_8_M3_d N_8_M4_s
+ N_8_M16_d N_8_c_264_n N_8_M17_s N_8_c_310_p N_8_c_276_n N_8_c_265_n
+ N_8_c_311_p N_8_c_267_n N_8_c_283_n N_8_c_284_n N_8_c_268_n N_8_c_312_p
+ N_8_c_269_n N_8_c_286_n N_8_c_288_n N_8_c_302_n N_8_c_271_n N_8_c_303_n
+ N_8_c_272_n N_8_c_295_n N_8_c_273_n N_8_c_274_n N_8_c_275_n VSS
+ PM_DFFHQNX2_ASAP7_75T_SRAM%8
x_PM_DFFHQNX2_ASAP7_75T_SRAM%9 N_9_M9_g N_9_c_320_p N_9_M22_g N_9_M10_d N_9_M23_d
+ N_9_c_319_p N_9_c_331_p N_9_c_318_p N_9_c_323_p N_9_c_317_p N_9_c_327_p
+ N_9_c_329_p N_9_c_328_p N_9_c_332_p N_9_c_336_p N_9_c_334_p N_9_c_330_p
+ N_9_c_322_p VSS PM_DFFHQNX2_ASAP7_75T_SRAM%9
x_PM_DFFHQNX2_ASAP7_75T_SRAM%10 N_10_M10_g N_10_M23_g N_10_M11_g N_10_M24_g
+ N_10_M12_g N_10_c_387_p N_10_M25_g N_10_M8_s N_10_M7_d N_10_c_338_n N_10_M21_s
+ N_10_M20_d N_10_c_348_n N_10_c_370_n N_10_c_339_n N_10_c_340_n N_10_c_400_p
+ N_10_c_342_n N_10_c_362_n N_10_c_349_n N_10_c_343_n N_10_c_350_n N_10_c_351_n
+ N_10_c_375_n N_10_c_353_n N_10_c_376_n N_10_c_378_n N_10_c_379_n N_10_c_380_n
+ N_10_c_354_n N_10_c_355_n N_10_c_381_n N_10_c_344_n N_10_c_386_n VSS
+ PM_DFFHQNX2_ASAP7_75T_SRAM%10
x_PM_DFFHQNX2_ASAP7_75T_SRAM%QN N_QN_M12_d N_QN_M11_d N_QN_M25_d N_QN_M24_d
+ N_QN_c_407_n N_QN_c_403_n N_QN_c_410_n N_QN_c_404_n QN N_QN_c_414_n VSS
+ PM_DFFHQNX2_ASAP7_75T_SRAM%QN
x_PM_DFFHQNX2_ASAP7_75T_SRAM%12 N_12_M2_d N_12_M3_s N_12_c_416_n VSS
+ PM_DFFHQNX2_ASAP7_75T_SRAM%12
x_PM_DFFHQNX2_ASAP7_75T_SRAM%13 N_13_M17_d N_13_M18_s N_13_c_423_n VSS
+ PM_DFFHQNX2_ASAP7_75T_SRAM%13
x_PM_DFFHQNX2_ASAP7_75T_SRAM%14 N_14_M8_d N_14_M9_s N_14_c_432_n VSS
+ PM_DFFHQNX2_ASAP7_75T_SRAM%14
x_PM_DFFHQNX2_ASAP7_75T_SRAM%15 N_15_M5_s N_15_M4_d VSS PM_DFFHQNX2_ASAP7_75T_SRAM%15
x_PM_DFFHQNX2_ASAP7_75T_SRAM%16 N_16_M16_s N_16_M15_d VSS
+ PM_DFFHQNX2_ASAP7_75T_SRAM%16
x_PM_DFFHQNX2_ASAP7_75T_SRAM%17 N_17_M22_s N_17_M21_d VSS
+ PM_DFFHQNX2_ASAP7_75T_SRAM%17
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_22_n 3.57152e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 CLK N_4_c_23_n 0.00136255f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.144
cc_4 CLK N_4_c_24_n 2.75361e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.07
cc_5 CLK N_4_c_25_n 0.00136255f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.107
cc_6 N_CLK_c_6_p N_4_c_26_n 0.00145637f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2
cc_7 N_CLK_c_6_p N_4_c_27_n 2.75361e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2125
cc_8 CLK N_4_c_28_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_6_p N_4_c_29_n 5.03453e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_6_p N_4_c_30_n 0.00123168f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.153
cc_11 CLK N_4_c_31_n 4.93618e-19 $X=0.082 $Y=0.119 $X2=0.175 $Y2=0.153
cc_12 N_CLK_c_6_p N_4_c_31_n 0.00162391f $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_13 N_CLK_c_13_p N_4_c_33_n 0.00115059f $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.135
cc_14 CLK N_4_c_34_n 0.00174864f $X=0.082 $Y=0.119 $X2=0.151 $Y2=0.135
cc_15 N_CLK_c_6_p N_4_c_34_n 3.32041e-19 $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.135
cc_16 CLK N_6_c_116_n 6.37157e-19 $X=0.082 $Y=0.119 $X2=0.027 $Y2=0.234
cc_17 N_CLK_c_6_p N_6_c_117_n 6.45547e-19 $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.153
cc_18 N_CLK_c_6_p N_6_c_118_n 0.00125366f $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_19 N_CLK_c_6_p N_6_c_119_n 4.3806e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_20 CLK N_6_c_120_n 0.00137619f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.153
cc_21 N_4_M3_g N_D_M2_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_22 N_4_c_37_p N_D_c_99_n 2.91747e-19 $X=0.527 $Y=0.153 $X2=0.081 $Y2=0.135
cc_23 N_4_c_33_n N_D_c_99_n 2.1478e-19 $X=0.151 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_4_c_39_p N_D_c_101_n 2.3983e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_25 N_4_c_40_p N_D_c_102_n 8.99815e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_26 N_4_c_40_p N_D_c_103_n 8.75229e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_27 N_4_M3_g N_6_c_121_n 0.00355599f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_28 N_4_c_43_p N_6_c_121_n 0.00126153f $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.054
cc_29 N_4_M3_g N_6_M4_g 0.00355599f $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_4_M8_g N_6_M7_g 0.00355599f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_31 N_4_M8_g N_6_c_125_n 0.00355599f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_32 N_4_M8_g N_6_c_126_n 0.00250257f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_33 N_4_c_48_p N_6_c_126_n 0.00180656f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_34 N_4_c_49_p N_6_c_126_n 6.4075e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_35 N_4_c_37_p N_6_c_126_n 0.00187561f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_36 N_4_c_51_p N_6_c_126_n 0.00123876f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_34_n N_6_c_116_n 2.97444e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_31_n N_6_c_132_n 2.38327e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_34_n N_6_c_117_n 2.85146e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_40_p N_6_c_118_n 2.46239e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_41 N_4_c_31_n N_6_c_135_n 2.31165e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_42 N_4_c_39_p N_6_c_136_n 9.24693e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_43 N_4_c_37_p N_6_c_137_n 3.67557e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_44 N_4_c_37_p N_6_c_138_n 8.06691e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_45 N_4_c_37_p N_6_c_139_n 2.46239e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_46 N_4_c_40_p N_6_c_119_n 0.0299327f $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_39_p N_6_c_119_n 2.98936e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_48 N_4_c_37_p N_6_c_142_n 2.81476e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_49 N_4_c_40_p N_6_c_143_n 8.79704e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_50 N_4_c_34_n N_6_c_143_n 0.00524677f $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_51 N_4_c_37_p N_6_c_145_n 9.92294e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_52 N_4_c_39_p N_6_c_145_n 5.5596e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_53 N_4_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_54 N_4_c_69_p N_7_c_219_n 3.42573e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_55 N_4_c_69_p N_7_c_220_n 5.29207e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_56 N_4_c_51_p N_7_c_221_n 0.00318218f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_57 N_4_c_49_p N_7_c_222_n 0.00115177f $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_58 N_4_c_49_p N_7_c_223_n 3.42573e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_59 N_4_M8_g N_8_M6_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_60 N_4_c_48_p N_8_c_262_n 3.88499e-19 $X=0.675 $Y=0.135 $X2=0.081 $Y2=0.135
cc_61 N_4_c_69_p N_8_c_262_n 3.00379e-19 $X=0.601 $Y=0.153 $X2=0.081 $Y2=0.135
cc_62 N_4_c_39_p N_8_c_264_n 2.36208e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_63 N_4_M3_g N_8_c_265_n 3.49806e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_4_c_39_p N_8_c_265_n 3.83282e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_65 N_4_c_39_p N_8_c_267_n 7.25941e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_66 N_4_c_39_p N_8_c_268_n 7.25941e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_67 N_4_c_37_p N_8_c_269_n 0.00118282f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_68 N_4_c_39_p N_8_c_269_n 8.1935e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_69 N_4_c_37_p N_8_c_271_n 0.00132871f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_70 N_4_c_69_p N_8_c_272_n 0.00132871f $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_71 N_4_c_37_p N_8_c_273_n 2.54113e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_72 N_4_c_37_p N_8_c_274_n 3.92135e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_73 N_4_c_39_p N_8_c_275_n 7.25941e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_74 N_4_M8_g N_9_M9_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_75 N_4_c_49_p N_10_c_338_n 2.24654e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_76 N_4_c_49_p N_10_c_339_n 5.06919e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_77 N_4_M8_g N_10_c_340_n 3.47752e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_78 N_4_c_51_p N_10_c_340_n 5.72565e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_79 N_4_c_49_p N_10_c_342_n 2.46558e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_80 N_4_c_51_p N_10_c_343_n 0.00319993f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_81 N_4_c_49_p N_10_c_344_n 2.9112e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_82 N_4_c_37_p N_12_c_416_n 3.46326e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_83 N_D_M2_g N_6_c_121_n 0.00341068f $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_84 N_D_c_99_n N_6_c_121_n 0.00114686f $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_85 D N_6_c_149_n 0.00215667f $X=0.244 $Y=0.082 $X2=0.0505 $Y2=0.234
cc_86 N_D_c_103_n N_6_c_150_n 0.00215667f $X=0.243 $Y=0.135 $X2=0.405 $Y2=0.153
cc_87 N_D_c_103_n N_6_c_118_n 0.00225008f $X=0.243 $Y=0.135 $X2=0.175 $Y2=0.153
cc_88 N_D_c_109_p N_6_c_137_n 0.00127755f $X=0.281 $Y=0.135 $X2=0.151 $Y2=0.135
cc_89 N_D_c_99_n N_6_c_119_n 2.11668e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_90 N_D_c_103_n N_6_c_119_n 0.00122387f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_91 D N_6_c_120_n 0.00215667f $X=0.244 $Y=0.082 $X2=0.018 $Y2=0.153
cc_92 N_D_c_113_p N_6_c_143_n 0.00215667f $X=0.243 $Y=0.126 $X2=0 $Y2=0
cc_93 N_D_c_103_n N_6_c_145_n 0.00120973f $X=0.243 $Y=0.135 $X2=0.027 $Y2=0.153
cc_94 N_D_c_103_n N_8_c_276_n 2.80198e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_95 N_6_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_96 N_6_M7_g N_7_M5_g 2.13359e-19 $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_97 N_6_c_126_n N_7_M5_g 0.00205997f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_98 N_6_c_142_n N_7_M5_g 3.15189e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_99 N_6_c_126_n N_7_c_228_n 6.55731e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_100 N_6_c_126_n N_7_c_229_n 2.12581e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_101 N_6_c_126_n N_7_M20_s 2.50995e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_102 N_6_M7_g N_7_c_231_n 0.00200065f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_103 N_6_c_126_n N_7_c_231_n 0.00312129f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_104 N_6_c_126_n N_7_c_220_n 3.41745e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_105 N_6_M7_g N_7_c_221_n 3.41702e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_106 N_6_M7_g N_7_c_222_n 2.26424e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_107 N_6_c_142_n N_7_c_236_n 5.75704e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_108 N_6_c_171_p N_7_c_237_n 0.00195059f $X=0.621 $Y=0.178 $X2=0 $Y2=0
cc_109 N_6_c_126_n N_7_c_237_n 0.00191847f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_110 N_6_M7_g N_7_c_239_n 3.8308e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_111 N_6_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_112 N_6_M7_g N_8_M6_g 0.00341068f $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_113 N_6_c_126_n N_8_M6_g 0.00302156f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_114 N_6_c_119_n N_8_c_264_n 3.12535e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_115 N_6_c_145_n N_8_c_264_n 8.9852e-19 $X=0.324 $Y=0.167 $X2=0 $Y2=0
cc_116 N_6_c_119_n N_8_c_276_n 0.0015935f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_117 N_6_M4_g N_8_c_283_n 3.68551e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_118 N_6_M4_g N_8_c_284_n 2.06635e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_119 N_6_M4_g N_8_c_269_n 2.27069e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_120 N_6_c_183_p N_8_c_286_n 4.73369e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_121 N_6_c_142_n N_8_c_286_n 0.00174159f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_122 N_6_c_183_p N_8_c_288_n 0.00171407f $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_123 N_6_c_126_n N_8_c_288_n 5.88593e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_124 N_6_c_119_n N_8_c_288_n 0.00104904f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_125 N_6_c_188_p N_8_c_288_n 2.15173e-19 $X=0.324 $Y=0.178 $X2=0 $Y2=0
cc_126 N_6_c_126_n N_8_c_271_n 8.16411e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_127 N_6_c_126_n N_8_c_272_n 3.32592e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_128 N_6_c_142_n N_8_c_272_n 8.9822e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_129 N_6_c_126_n N_8_c_295_n 4.02972e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_130 N_6_c_125_n N_9_M9_g 0.00341068f $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_131 N_6_c_125_n N_10_M10_g 2.13359e-19 $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_132 N_6_c_126_n N_10_c_338_n 8.27829e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_133 N_6_c_126_n N_10_M21_s 3.37661e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_134 N_6_c_126_n N_10_c_348_n 0.00145548f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_135 N_6_c_125_n N_10_c_349_n 3.03386e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_136 N_6_c_125_n N_10_c_350_n 2.58526e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_137 N_6_c_125_n N_10_c_351_n 0.00228871f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_138 N_6_c_126_n N_10_c_351_n 7.89371e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_139 N_6_c_125_n N_10_c_353_n 4.55487e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_140 N_6_c_126_n N_10_c_354_n 4.54272e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_141 N_6_c_125_n N_10_c_355_n 5.68093e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_142 N_6_c_126_n N_10_c_355_n 2.2968e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_143 N_6_c_121_n N_12_c_416_n 0.00514294f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_144 N_6_c_137_n N_12_c_416_n 0.00114179f $X=0.333 $Y=0.135 $X2=0 $Y2=0
cc_145 N_6_c_126_n N_13_M18_s 2.36286e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.216
cc_146 N_6_M4_g N_13_c_423_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_147 N_6_c_183_p N_13_c_423_n 5.41258e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_148 N_6_c_126_n N_13_c_423_n 0.00230928f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_149 N_6_c_119_n N_13_c_423_n 7.09553e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_150 N_6_c_125_n N_14_c_432_n 0.00198387f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_151 N_6_c_126_n N_14_c_432_n 4.51352e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_152 N_6_c_139_n N_16_M16_s 8.59575e-19 $X=0.324 $Y=0.189 $X2=0.081 $Y2=0.054
cc_153 N_6_c_145_n N_16_M16_s 2.57402e-19 $X=0.324 $Y=0.167 $X2=0.081 $Y2=0.054
cc_154 N_6_c_188_p N_16_M16_s 2.18007e-19 $X=0.324 $Y=0.178 $X2=0.081 $Y2=0.054
cc_155 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_156 N_7_c_241_p N_8_M6_g 3.87418e-19 $X=0.576 $Y=0.09 $X2=0.135 $Y2=0.054
cc_157 N_7_c_221_n N_8_c_262_n 2.20449e-19 $X=0.621 $Y=0.122 $X2=0.135 $Y2=0.135
cc_158 N_7_c_243_p N_8_c_283_n 3.63506e-19 $X=0.594 $Y=0.054 $X2=0.018 $Y2=0.107
cc_159 N_7_c_244_p N_8_c_284_n 3.19692e-19 $X=0.513 $Y=0.09 $X2=0.018 $Y2=0.162
cc_160 N_7_c_241_p N_8_c_284_n 0.00114151f $X=0.576 $Y=0.09 $X2=0.018 $Y2=0.162
cc_161 N_7_c_246_p N_8_c_302_n 7.39815e-19 $X=0.621 $Y=0.14 $X2=0.027 $Y2=0.234
cc_162 N_7_c_241_p N_8_c_303_n 0.0047777f $X=0.576 $Y=0.09 $X2=0.054 $Y2=0.234
cc_163 N_7_M5_g N_8_c_272_n 3.12986e-19 $X=0.513 $Y=0.0405 $X2=0.047 $Y2=0.234
cc_164 N_7_c_244_p N_8_c_273_n 5.2508e-19 $X=0.513 $Y=0.09 $X2=0.033 $Y2=0.153
cc_165 N_7_c_228_n N_10_c_338_n 0.0027803f $X=0.594 $Y=0.0405 $X2=0 $Y2=0
cc_166 N_7_c_243_p N_10_c_338_n 3.72596e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_167 N_7_c_239_n N_10_c_338_n 3.30531e-19 $X=0.621 $Y=0.09 $X2=0 $Y2=0
cc_168 N_7_c_231_n N_10_c_348_n 0.00220898f $X=0.65 $Y=0.2295 $X2=0 $Y2=0
cc_169 N_7_c_228_n N_10_c_339_n 5.23227e-19 $X=0.594 $Y=0.0405 $X2=0.018
+ $Y2=0.225
cc_170 N_7_c_243_p N_10_c_362_n 2.3746e-19 $X=0.594 $Y=0.054 $X2=0.054 $Y2=0.036
cc_171 N_7_c_239_n N_10_c_349_n 4.46294e-19 $X=0.621 $Y=0.09 $X2=0.047 $Y2=0.036
cc_172 N_7_c_237_n N_10_c_351_n 4.46294e-19 $X=0.621 $Y=0.203 $X2=0.054
+ $Y2=0.234
cc_173 N_7_c_231_n N_10_c_354_n 3.64147e-19 $X=0.65 $Y=0.2295 $X2=0 $Y2=0
cc_174 N_7_c_220_n N_10_c_354_n 4.68959e-19 $X=0.612 $Y=0.234 $X2=0 $Y2=0
cc_175 N_7_c_260_p N_10_c_355_n 4.46294e-19 $X=0.621 $Y=0.101 $X2=0.151
+ $Y2=0.135
cc_176 N_8_c_264_n N_12_c_416_n 0.00119486f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_177 N_8_c_273_n N_12_c_416_n 0.00390673f $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_178 N_8_c_274_n N_12_c_416_n 5.36233e-19 $X=0.45 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_179 N_8_c_264_n N_13_c_423_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_180 N_8_c_310_p N_13_c_423_n 0.00209454f $X=0.45 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_181 N_8_c_311_p N_13_c_423_n 0.0013184f $X=0.434 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_182 N_8_c_312_p N_13_c_423_n 0.00119522f $X=0.459 $Y=0.225 $X2=0.405
+ $Y2=0.0675
cc_183 N_8_c_273_n N_13_c_423_n 5.72158e-19 $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_184 N_9_M9_g N_10_M10_g 0.00268443f $X=0.783 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_185 N_9_c_317_p N_10_M10_g 3.74489e-19 $X=0.846 $Y=0.036 $X2=0.135 $Y2=0.054
cc_186 N_9_c_318_p N_10_c_370_n 0.00141609f $X=0.792 $Y=0.036 $X2=0.018
+ $Y2=0.045
cc_187 N_9_c_319_p N_10_c_362_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.054
+ $Y2=0.036
cc_188 N_9_c_320_p N_10_c_349_n 3.34766e-19 $X=0.783 $Y=0.1055 $X2=0.047
+ $Y2=0.036
cc_189 N_9_c_319_p N_10_c_349_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.047
+ $Y2=0.036
cc_190 N_9_c_322_p N_10_c_351_n 2.42078e-19 $X=0.945 $Y=0.216 $X2=0.054
+ $Y2=0.234
cc_191 N_9_c_323_p N_10_c_375_n 2.6154e-19 $X=0.828 $Y=0.036 $X2=0.054 $Y2=0.234
cc_192 N_9_M9_g N_10_c_376_n 6.3699e-19 $X=0.783 $Y=0.0405 $X2=0.0505 $Y2=0.234
cc_193 N_9_c_319_p N_10_c_376_n 9.10342e-19 $X=0.783 $Y=0.105 $X2=0.0505
+ $Y2=0.234
cc_194 N_9_c_317_p N_10_c_378_n 4.40983e-19 $X=0.846 $Y=0.036 $X2=0.033
+ $Y2=0.153
cc_195 N_9_c_327_p N_10_c_379_n 5.13693e-19 $X=0.882 $Y=0.036 $X2=0.405
+ $Y2=0.153
cc_196 N_9_c_328_p N_10_c_380_n 0.00149072f $X=0.9 $Y=0.234 $X2=0.405 $Y2=0.153
cc_197 N_9_c_329_p N_10_c_381_n 4.52584e-19 $X=0.9 $Y=0.036 $X2=0 $Y2=0
cc_198 N_9_c_330_p N_10_c_381_n 0.00299425f $X=0.945 $Y=0.167 $X2=0 $Y2=0
cc_199 N_9_c_331_p N_10_c_344_n 2.40515e-19 $X=0.936 $Y=0.036 $X2=0 $Y2=0
cc_200 N_9_c_332_p N_10_c_344_n 7.44774e-19 $X=0.918 $Y=0.234 $X2=0 $Y2=0
cc_201 N_9_c_330_p N_10_c_344_n 8.84468e-19 $X=0.945 $Y=0.167 $X2=0 $Y2=0
cc_202 N_9_c_334_p N_10_c_386_n 0.00323217f $X=0.945 $Y=0.117 $X2=0 $Y2=0
cc_203 N_9_c_331_p N_QN_c_403_n 4.0695e-19 $X=0.936 $Y=0.036 $X2=0 $Y2=0
cc_204 N_9_c_336_p N_QN_c_404_n 4.04283e-19 $X=0.945 $Y=0.225 $X2=0 $Y2=0
cc_205 N_9_c_318_p N_14_c_432_n 7.33799e-19 $X=0.792 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_206 N_10_c_387_p N_QN_M12_d 3.7444e-19 $X=1.053 $Y=0.136 $X2=0.135 $Y2=0.054
cc_207 N_10_c_387_p N_QN_M25_d 3.85232e-19 $X=1.053 $Y=0.136 $X2=0.135 $Y2=0.216
cc_208 N_10_c_387_p N_QN_c_407_n 8.43851e-19 $X=1.053 $Y=0.136 $X2=0.405
+ $Y2=0.0675
cc_209 N_10_M12_g N_QN_c_403_n 4.75199e-19 $X=1.053 $Y=0.0675 $X2=0 $Y2=0
cc_210 N_10_c_387_p N_QN_c_403_n 5.85953e-19 $X=1.053 $Y=0.136 $X2=0 $Y2=0
cc_211 N_10_c_387_p N_QN_c_410_n 7.60428e-19 $X=1.053 $Y=0.136 $X2=0.405
+ $Y2=0.2295
cc_212 N_10_c_386_n N_QN_c_410_n 6.27685e-19 $X=0.999 $Y=0.136 $X2=0.405
+ $Y2=0.2295
cc_213 N_10_M12_g N_QN_c_404_n 4.69796e-19 $X=1.053 $Y=0.0675 $X2=0 $Y2=0
cc_214 N_10_c_387_p N_QN_c_404_n 5.9664e-19 $X=1.053 $Y=0.136 $X2=0 $Y2=0
cc_215 N_10_c_387_p N_QN_c_414_n 3.65635e-19 $X=1.053 $Y=0.136 $X2=0.056
+ $Y2=0.054
cc_216 N_10_c_386_n N_QN_c_414_n 9.88669e-19 $X=0.999 $Y=0.136 $X2=0.056
+ $Y2=0.054
cc_217 N_10_c_338_n N_14_c_432_n 0.00182708f $X=0.648 $Y=0.0405 $X2=0.405
+ $Y2=0.0675
cc_218 N_10_c_370_n N_14_c_432_n 0.0020512f $X=0.72 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_219 N_10_c_400_p N_14_c_432_n 0.00131745f $X=0.704 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_220 N_10_c_362_n N_14_c_432_n 0.00103589f $X=0.729 $Y=0.081 $X2=0.405
+ $Y2=0.0675
cc_221 N_10_c_353_n N_14_c_432_n 4.02739e-19 $X=0.774 $Y=0.162 $X2=0.405
+ $Y2=0.0675

* END of "./DFFHQNx2_ASAP7_75t_SRAM.pex.sp.DFFHQNX2_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DFFHQNx3_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:24:53 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DFFHQNx3_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DFFHQNx3_ASAP7_75t_SRAM.pex.sp.pex"
* File: DFFHQNx3_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:24:53 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%CLK 2 5 7 12 14 VSS
c20 14 VSS 0.00674559f $X=0.081 $Y=0.135
c21 12 VSS 0.00682604f $X=0.082 $Y=0.119
c22 5 VSS 0.00206449f $X=0.081 $Y=0.135
c23 2 VSS 0.0629f $X=0.081 $Y=0.054
r24 12 14 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.135
r25 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r26 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r27 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%4 2 7 10 13 15 18 21 23 25 28 30 36 37 38 41 42
+ 45 52 59 67 68 70 72 73 78 79 83 88 VSS
c77 114 VSS 1.06551e-19 $X=0.03 $Y=0.153
c78 113 VSS 6.89947e-19 $X=0.027 $Y=0.153
c79 88 VSS 0.00102973f $X=0.675 $Y=0.135
c80 83 VSS 8.66895e-19 $X=0.405 $Y=0.135
c81 79 VSS 0.00121012f $X=0.151 $Y=0.135
c82 78 VSS 0.00390107f $X=0.151 $Y=0.135
c83 73 VSS 0.00263053f $X=0.601 $Y=0.153
c84 72 VSS 0.00556612f $X=0.527 $Y=0.153
c85 70 VSS 0.00405122f $X=0.675 $Y=0.153
c86 68 VSS 0.00330975f $X=0.29 $Y=0.153
c87 67 VSS 0.00602706f $X=0.175 $Y=0.153
c88 59 VSS 6.74716e-19 $X=0.033 $Y=0.153
c89 55 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c90 54 VSS 0.00180216f $X=0.047 $Y=0.234
c91 52 VSS 0.00250119f $X=0.054 $Y=0.234
c92 50 VSS 0.00305101f $X=0.027 $Y=0.234
c93 48 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c94 47 VSS 0.00199699f $X=0.047 $Y=0.036
c95 45 VSS 0.00250119f $X=0.054 $Y=0.036
c96 43 VSS 0.00305101f $X=0.027 $Y=0.036
c97 42 VSS 4.88707e-19 $X=0.018 $Y=0.2125
c98 41 VSS 0.00180713f $X=0.018 $Y=0.2
c99 40 VSS 4.69158e-19 $X=0.018 $Y=0.225
c100 38 VSS 0.00173342f $X=0.018 $Y=0.107
c101 37 VSS 9.57865e-19 $X=0.018 $Y=0.07
c102 36 VSS 0.00172854f $X=0.018 $Y=0.144
c103 33 VSS 0.00509483f $X=0.056 $Y=0.216
c104 30 VSS 2.98509e-19 $X=0.071 $Y=0.216
c105 28 VSS 0.00497933f $X=0.056 $Y=0.054
c106 25 VSS 2.98509e-19 $X=0.071 $Y=0.054
c107 21 VSS 0.00214819f $X=0.675 $Y=0.135
c108 18 VSS 0.0585656f $X=0.675 $Y=0.0405
c109 13 VSS 0.00214124f $X=0.405 $Y=0.135
c110 10 VSS 0.058827f $X=0.405 $Y=0.0675
c111 2 VSS 0.0628024f $X=0.135 $Y=0.054
r112 113 114 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r113 110 113 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r114 78 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.151 $Y=0.135 $X2=0.151
+ $Y2=0.135
r115 72 73 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.601 $Y2=0.153
r116 70 73 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.675
+ $Y=0.153 $X2=0.601 $Y2=0.153
r117 70 88 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.675 $Y=0.153 $X2=0.675
+ $Y2=0.153
r118 67 68 7.80864 $w=1.8e-08 $l=1.15e-07 $layer=M2 $thickness=3.6e-08 $X=0.175
+ $Y=0.153 $X2=0.29 $Y2=0.153
r119 65 72 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.527 $Y2=0.153
r120 65 68 7.80864 $w=1.8e-08 $l=1.15e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.29 $Y2=0.153
r121 65 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r122 62 67 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.151
+ $Y=0.153 $X2=0.175 $Y2=0.153
r123 62 79 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.151 $Y=0.153 $X2=0.151
+ $Y2=0.153
r124 59 114 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r125 58 62 8.01235 $w=1.8e-08 $l=1.18e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.151 $Y2=0.153
r126 58 59 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r127 54 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r128 52 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r129 50 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r130 47 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r131 45 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r132 43 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r133 41 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r134 40 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r135 40 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r136 39 110 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r137 39 41 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.2
r138 37 38 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.107
r139 36 110 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r140 36 38 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.107
r141 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r142 35 37 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r143 33 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r144 30 33 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r145 28 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r146 25 28 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r147 21 88 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.135 $X2=0.675
+ $Y2=0.135
r148 21 23 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2295
r149 18 21 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.135
r150 13 83 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r151 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2295
r152 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r153 5 78 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.151 $Y2=0.135
r154 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r155 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%D 2 5 7 10 12 14 21 23 28 VSS
c18 28 VSS 0.00931225f $X=0.243 $Y=0.135
c19 24 VSS 2.45662e-20 $X=0.276 $Y=0.135
c20 23 VSS 0.00111822f $X=0.271 $Y=0.135
c21 21 VSS 2.56376e-19 $X=0.281 $Y=0.135
c22 14 VSS 2.7811e-19 $X=0.243 $Y=0.116
c23 12 VSS 0.00925957f $X=0.244 $Y=0.082
c24 10 VSS 2.38113e-19 $X=0.243 $Y=0.126
c25 5 VSS 0.00522238f $X=0.297 $Y=0.135
c26 2 VSS 0.0630392f $X=0.297 $Y=0.0675
r27 23 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.271
+ $Y=0.135 $X2=0.276 $Y2=0.135
r28 21 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.281
+ $Y=0.135 $X2=0.276 $Y2=0.135
r29 21 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.281 $Y=0.135 $X2=0.281
+ $Y2=0.135
r30 19 28 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.243 $Y2=0.135
r31 19 23 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.271 $Y2=0.135
r32 13 14 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.106 $X2=0.243 $Y2=0.116
r33 12 13 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.082 $X2=0.243 $Y2=0.106
r34 10 28 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.135
r35 10 14 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.116
r36 5 22 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.281 $Y2=0.135
r37 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r38 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%6 2 5 8 14 17 20 23 28 35 39 44 50 55 57 61 66
+ 67 68 75 77 78 87 89 105 110 111 113 114 VSS
c102 114 VSS 2.23151e-19 $X=0.324 $Y=0.178
c103 113 VSS 4.08645e-19 $X=0.324 $Y=0.167
c104 111 VSS 7.77947e-19 $X=0.189 $Y=0.167
c105 110 VSS 9.60988e-19 $X=0.189 $Y=0.106
c106 105 VSS 6.81413e-19 $X=0.513 $Y=0.18
c107 89 VSS 0.0113851f $X=0.513 $Y=0.189
c108 87 VSS 0.00141172f $X=0.324 $Y=0.189
c109 78 VSS 4.01771e-19 $X=0.342 $Y=0.135
c110 77 VSS 5.28662e-19 $X=0.333 $Y=0.135
c111 75 VSS 7.4105e-19 $X=0.351 $Y=0.135
c112 68 VSS 0.00169555f $X=0.18 $Y=0.234
c113 67 VSS 9.43175e-19 $X=0.189 $Y=0.225
c114 66 VSS 0.00196236f $X=0.189 $Y=0.234
c115 61 VSS 0.00196921f $X=0.162 $Y=0.234
c116 57 VSS 0.00170883f $X=0.18 $Y=0.036
c117 55 VSS 0.00196236f $X=0.189 $Y=0.036
c118 50 VSS 0.00193426f $X=0.162 $Y=0.036
c119 47 VSS 0.00715944f $X=0.16 $Y=0.216
c120 42 VSS 0.00719538f $X=0.16 $Y=0.054
c121 35 VSS 0.0611368f $X=0.725 $Y=0.178
c122 28 VSS 0.00126548f $X=0.464 $Y=0.178
c123 20 VSS 0.0618767f $X=0.729 $Y=0.178
c124 17 VSS 1.08457e-19 $X=0.621 $Y=0.178
c125 14 VSS 0.0600454f $X=0.621 $Y=0.0405
c126 8 VSS 0.0602427f $X=0.459 $Y=0.0405
c127 2 VSS 0.0623279f $X=0.351 $Y=0.135
r128 113 114 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.324 $Y=0.167 $X2=0.324 $Y2=0.178
r129 110 111 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.106 $X2=0.189 $Y2=0.167
r130 104 105 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r131 89 105 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r132 87 114 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.189 $X2=0.324 $Y2=0.178
r133 86 89 12.8333 $w=1.8e-08 $l=1.89e-07 $layer=M2 $thickness=3.6e-08 $X=0.324
+ $Y=0.189 $X2=0.513 $Y2=0.189
r134 86 87 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.324 $Y=0.189 $X2=0.324
+ $Y2=0.189
r135 83 111 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.167
r136 82 86 9.16667 $w=1.8e-08 $l=1.35e-07 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.324 $Y2=0.189
r137 82 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.189 $X2=0.189
+ $Y2=0.189
r138 77 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.135 $X2=0.342 $Y2=0.135
r139 75 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.342 $Y2=0.135
r140 72 113 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.144 $X2=0.324 $Y2=0.167
r141 71 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.135 $X2=0.333 $Y2=0.135
r142 71 72 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.135 $X2=0.324 $Y2=0.144
r143 68 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r144 67 83 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.189
r145 66 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r146 66 67 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.189 $Y2=0.225
r147 61 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r148 57 58 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r149 56 110 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.106
r150 55 58 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r151 55 56 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r152 50 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r153 47 61 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r154 44 47 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r155 42 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r156 39 42 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r157 28 104 39.0385 $w=2.6e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.178 $X2=0.513 $Y2=0.178
r158 20 35 3.07692 $w=2.6e-08 $l=4e-09 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.178 $X2=0.725 $Y2=0.178
r159 20 23 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.178 $X2=0.729 $Y2=0.2295
r160 17 35 82.8571 $w=2.6e-08 $l=1.04e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.725 $Y2=0.178
r161 17 104 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.513 $Y2=0.178
r162 14 17 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0405 $X2=0.621 $Y2=0.178
r163 11 28 3.84615 $w=2.6e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.178 $X2=0.464 $Y2=0.178
r164 8 11 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.178
r165 2 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r166 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%7 2 5 7 9 10 13 14 17 19 22 29 30 31 38 43 44 45
+ 46 47 48 52 53 VSS
c43 54 VSS 3.52511e-19 $X=0.612 $Y=0.09
c44 53 VSS 1.80704e-19 $X=0.603 $Y=0.09
c45 52 VSS 5.96246e-19 $X=0.621 $Y=0.09
c46 49 VSS 6.86664e-19 $X=0.621 $Y=0.224
c47 48 VSS 4.95788e-19 $X=0.621 $Y=0.203
c48 47 VSS 1.19762e-19 $X=0.621 $Y=0.167
c49 46 VSS 3.19764e-19 $X=0.621 $Y=0.165
c50 45 VSS 3.13056e-19 $X=0.621 $Y=0.14
c51 44 VSS 3.62783e-19 $X=0.621 $Y=0.122
c52 43 VSS 1.48552e-19 $X=0.621 $Y=0.101
c53 38 VSS 0.00113884f $X=0.594 $Y=0.054
c54 31 VSS 0.00668633f $X=0.612 $Y=0.234
c55 30 VSS 3.5821e-19 $X=0.5805 $Y=0.09
c56 29 VSS 0.00257846f $X=0.576 $Y=0.09
c57 24 VSS 1.48201e-19 $X=0.585 $Y=0.09
c58 22 VSS 0.0179338f $X=0.65 $Y=0.2295
c59 19 VSS 3.14771e-19 $X=0.665 $Y=0.2295
c60 17 VSS 2.67274e-19 $X=0.592 $Y=0.2295
c61 13 VSS 0.0252201f $X=0.594 $Y=0.0405
c62 9 VSS 6.29543e-19 $X=0.611 $Y=0.0405
c63 5 VSS 0.00238279f $X=0.513 $Y=0.09
c64 2 VSS 0.0584396f $X=0.513 $Y=0.0405
r65 53 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.603
+ $Y=0.09 $X2=0.612 $Y2=0.09
r66 52 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.612 $Y2=0.09
r67 51 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.09 $X2=0.603 $Y2=0.09
r68 49 50 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.224 $X2=0.621 $Y2=0.2245
r69 48 49 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.224
r70 47 48 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.203
r71 46 47 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.167
r72 45 46 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r73 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r74 43 44 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.101 $X2=0.621 $Y2=0.122
r75 42 50 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.2245
r76 41 52 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.09
r77 41 43 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.101
r78 36 51 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.09
r79 36 38 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.054
r80 31 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r81 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r82 29 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.09 $X2=0.5805 $Y2=0.09
r83 26 29 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.09 $X2=0.576 $Y2=0.09
r84 24 51 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.594 $Y2=0.09
r85 24 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.5805 $Y2=0.09
r86 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2295 $X2=0.65 $Y2=0.2295
r87 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.592
+ $Y=0.2295 $X2=0.65 $Y2=0.2295
r88 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r89 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r90 13 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.054 $X2=0.594
+ $Y2=0.054
r91 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.594 $Y2=0.0405
r92 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0405 $X2=0.594 $Y2=0.0405
r93 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.09 $X2=0.513
+ $Y2=0.09
r94 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.09 $X2=0.513 $Y2=0.2295
r95 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.09
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%8 2 5 7 9 14 17 21 22 25 27 33 35 37 38 39 41 43
+ 44 45 46 50 52 53 54 55 59 62 65 VSS
c53 65 VSS 2.85958e-19 $X=0.459 $Y=0.131
c54 62 VSS 0.00341346f $X=0.45 $Y=0.036
c55 61 VSS 0.0025252f $X=0.459 $Y=0.036
c56 59 VSS 0.00276391f $X=0.432 $Y=0.036
c57 55 VSS 4.23521e-19 $X=0.5445 $Y=0.131
c58 54 VSS 3.49205e-20 $X=0.522 $Y=0.131
c59 53 VSS 2.00095e-19 $X=0.504 $Y=0.131
c60 52 VSS 0.00133241f $X=0.496 $Y=0.131
c61 50 VSS 2.94642e-19 $X=0.567 $Y=0.131
c62 47 VSS 4.32029e-19 $X=0.459 $Y=0.214
c63 46 VSS 2.06877e-19 $X=0.459 $Y=0.203
c64 45 VSS 6.09344e-21 $X=0.459 $Y=0.167
c65 44 VSS 2.12612e-19 $X=0.459 $Y=0.165
c66 43 VSS 2.51143e-19 $X=0.459 $Y=0.225
c67 41 VSS 3.68971e-19 $X=0.459 $Y=0.114
c68 40 VSS 3.4692e-19 $X=0.459 $Y=0.106
c69 38 VSS 7.88894e-19 $X=0.459 $Y=0.081
c70 37 VSS 2.0833e-19 $X=0.459 $Y=0.122
c71 35 VSS 0.00142907f $X=0.434 $Y=0.234
c72 34 VSS 3.2912e-19 $X=0.418 $Y=0.234
c73 33 VSS 0.00146362f $X=0.414 $Y=0.234
c74 32 VSS 0.00227054f $X=0.396 $Y=0.234
c75 27 VSS 0.00148441f $X=0.378 $Y=0.234
c76 25 VSS 0.00389542f $X=0.45 $Y=0.234
c77 24 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c78 21 VSS 0.00379676f $X=0.378 $Y=0.2025
c79 18 VSS 1.15515e-19 $X=0.3735 $Y=0.216
c80 16 VSS 5.70081e-19 $X=0.432 $Y=0.0405
c81 10 VSS 7.61325e-20 $X=0.4275 $Y=0.054
c82 5 VSS 0.0022736f $X=0.567 $Y=0.1305
c83 2 VSS 0.0591678f $X=0.567 $Y=0.0405
r84 62 63 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r85 61 63 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r86 58 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r87 58 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r88 54 55 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r89 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r90 52 53 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.496
+ $Y=0.131 $X2=0.504 $Y2=0.131
r91 50 55 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r92 48 65 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r93 48 52 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.496 $Y2=0.131
r94 46 47 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.203 $X2=0.459 $Y2=0.214
r95 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.167 $X2=0.459 $Y2=0.203
r96 44 45 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.167
r97 43 47 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r98 42 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r99 42 44 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.165
r100 40 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.106 $X2=0.459 $Y2=0.114
r101 39 40 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.099 $X2=0.459 $Y2=0.106
r102 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.099
r103 37 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r104 37 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.114
r105 36 61 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r106 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.081
r107 34 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.234 $X2=0.434 $Y2=0.234
r108 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.418 $Y2=0.234
r109 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r110 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r111 25 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r112 25 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.434 $Y2=0.234
r113 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r114 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r115 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r116 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r117 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r118 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r119 13 59 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r120 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r121 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r122 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r123 5 50 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.131 $X2=0.567
+ $Y2=0.131
r124 5 7 370.904 $w=2e-08 $l=9.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1305 $X2=0.567 $Y2=0.2295
r125 2 5 337.185 $w=2e-08 $l=9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.1305
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%9 2 5 7 9 14 21 25 26 30 31 32 33 34 39 40 42 44
+ 45 VSS
c24 46 VSS 2.31795e-19 $X=0.945 $Y=0.171
c25 45 VSS 0.0010039f $X=0.945 $Y=0.167
c26 44 VSS 2.58105e-19 $X=0.945 $Y=0.122
c27 43 VSS 0.00381805f $X=0.945 $Y=0.117
c28 42 VSS 0.00298997f $X=0.945 $Y=0.225
c29 40 VSS 0.0018377f $X=0.918 $Y=0.234
c30 39 VSS 0.00568507f $X=0.9 $Y=0.234
c31 34 VSS 0.00462933f $X=0.936 $Y=0.234
c32 33 VSS 0.00189638f $X=0.9 $Y=0.036
c33 32 VSS 0.0035379f $X=0.882 $Y=0.036
c34 31 VSS 0.00146362f $X=0.846 $Y=0.036
c35 30 VSS 0.00510392f $X=0.828 $Y=0.036
c36 26 VSS 0.00226308f $X=0.792 $Y=0.036
c37 25 VSS 0.00657446f $X=0.936 $Y=0.036
c38 21 VSS 0.00122443f $X=0.783 $Y=0.105
c39 17 VSS 0.00481511f $X=0.862 $Y=0.2295
c40 12 VSS 0.00513464f $X=0.862 $Y=0.0405
c41 5 VSS 0.00277722f $X=0.783 $Y=0.1055
c42 2 VSS 0.0590816f $X=0.783 $Y=0.0405
r43 45 46 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.167 $X2=0.945 $Y2=0.171
r44 44 45 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.122 $X2=0.945 $Y2=0.167
r45 43 44 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.117 $X2=0.945 $Y2=0.122
r46 42 46 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.171
r47 41 43 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.117
r48 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.234 $X2=0.918 $Y2=0.234
r49 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.9 $Y2=0.234
r50 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r51 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.918 $Y2=0.234
r52 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r53 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.846 $Y2=0.036
r54 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r55 28 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.846 $Y2=0.036
r56 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.036 $X2=0.828 $Y2=0.036
r57 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r58 25 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.9 $Y2=0.036
r59 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.783 $Y=0.045 $X2=0.792 $Y2=0.036
r60 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.105
r61 17 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234 $X2=0.864
+ $Y2=0.234
r62 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2295 $X2=0.862 $Y2=0.2295
r63 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036 $X2=0.864
+ $Y2=0.036
r64 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.862 $Y2=0.0405
r65 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.105 $X2=0.783
+ $Y2=0.105
r66 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.1055 $X2=0.783 $Y2=0.2295
r67 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.1055
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%10 2 7 10 15 18 23 26 29 31 33 34 37 38 39 42 43
+ 48 49 51 53 54 55 56 57 59 60 62 63 66 73 74 82 85 89 92 100 VSS
c66 100 VSS 0.00121049f $X=0.999 $Y=0.136
c67 92 VSS 0.0079578f $X=0.999 $Y=0.153
c68 89 VSS 0.00168283f $X=0.891 $Y=0.153
c69 86 VSS 4.17512e-19 $X=0.837 $Y=0.162
c70 85 VSS 1.52743e-19 $X=0.729 $Y=0.162
c71 82 VSS 0.00357121f $X=0.72 $Y=0.233
c72 81 VSS 0.00257308f $X=0.729 $Y=0.233
c73 74 VSS 4.30636e-19 $X=0.866 $Y=0.162
c74 73 VSS 1.23291e-19 $X=0.85 $Y=0.162
c75 71 VSS 2.75449e-19 $X=0.882 $Y=0.162
c76 66 VSS 3.94906e-19 $X=0.837 $Y=0.135
c77 63 VSS 3.26354e-19 $X=0.792 $Y=0.162
c78 62 VSS 0.00206921f $X=0.774 $Y=0.162
c79 60 VSS 0.00191548f $X=0.828 $Y=0.162
c80 59 VSS 0.00132112f $X=0.729 $Y=0.224
c81 57 VSS 1.52884e-19 $X=0.729 $Y=0.136
c82 56 VSS 2.77769e-19 $X=0.729 $Y=0.119
c83 55 VSS 1.41609e-19 $X=0.729 $Y=0.101
c84 54 VSS 3.52175e-19 $X=0.729 $Y=0.081
c85 53 VSS 2.73935e-19 $X=0.729 $Y=0.153
c86 51 VSS 0.00166757f $X=0.704 $Y=0.036
c87 50 VSS 4.5779e-19 $X=0.688 $Y=0.036
c88 49 VSS 0.00146362f $X=0.684 $Y=0.036
c89 48 VSS 0.00375563f $X=0.666 $Y=0.036
c90 43 VSS 0.00409736f $X=0.72 $Y=0.036
c91 42 VSS 0.00133398f $X=0.702 $Y=0.2295
c92 38 VSS 6.50675e-19 $X=0.719 $Y=0.2295
c93 37 VSS 0.0376609f $X=0.648 $Y=0.0405
c94 33 VSS 5.63046e-19 $X=0.665 $Y=0.0405
c95 29 VSS 0.0129248f $X=1.107 $Y=0.136
c96 26 VSS 0.0647964f $X=1.107 $Y=0.0675
c97 18 VSS 0.0617066f $X=1.053 $Y=0.0675
c98 10 VSS 0.0615046f $X=0.999 $Y=0.0675
c99 5 VSS 0.00239735f $X=0.837 $Y=0.135
c100 2 VSS 0.0618222f $X=0.837 $Y=0.0405
r101 92 100 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.999 $Y=0.153 $X2=0.999
+ $Y2=0.153
r102 88 92 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.999 $Y2=0.153
r103 88 89 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r104 82 83 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.233 $X2=0.7245 $Y2=0.233
r105 81 83 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.233 $X2=0.7245 $Y2=0.233
r106 78 82 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.233 $X2=0.72 $Y2=0.233
r107 73 74 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.85
+ $Y=0.162 $X2=0.866 $Y2=0.162
r108 72 86 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.837 $Y2=0.162
r109 72 73 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.85 $Y2=0.162
r110 71 89 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.891 $Y2=0.162
r111 71 74 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.866 $Y2=0.162
r112 64 86 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.162
r113 64 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.135
r114 62 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.162 $X2=0.792 $Y2=0.162
r115 61 85 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.729 $Y2=0.162
r116 61 62 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.774 $Y2=0.162
r117 60 86 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.837 $Y2=0.162
r118 60 63 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.792 $Y2=0.162
r119 59 81 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.224 $X2=0.729 $Y2=0.233
r120 58 85 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.162
r121 58 59 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.224
r122 56 57 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.119 $X2=0.729 $Y2=0.136
r123 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.101 $X2=0.729 $Y2=0.119
r124 54 55 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.081 $X2=0.729 $Y2=0.101
r125 53 85 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.162
r126 53 57 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.136
r127 52 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.045 $X2=0.729 $Y2=0.081
r128 50 51 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.036 $X2=0.704 $Y2=0.036
r129 49 50 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.688 $Y2=0.036
r130 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.684 $Y2=0.036
r131 45 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.666 $Y2=0.036
r132 43 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.036 $X2=0.729 $Y2=0.045
r133 43 51 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.704 $Y2=0.036
r134 42 78 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.233
+ $X2=0.702 $Y2=0.233
r135 39 42 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2295 $X2=0.702 $Y2=0.2295
r136 38 42 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2295 $X2=0.702 $Y2=0.2295
r137 37 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r138 34 37 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0405 $X2=0.648 $Y2=0.0405
r139 33 37 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r140 29 31 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.136 $X2=1.107 $Y2=0.2025
r141 26 29 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.0675 $X2=1.107 $Y2=0.136
r142 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.053
+ $Y=0.136 $X2=1.107 $Y2=0.136
r143 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.136 $X2=1.053 $Y2=0.2025
r144 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.0675 $X2=1.053 $Y2=0.136
r145 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.999
+ $Y=0.136 $X2=1.053 $Y2=0.136
r146 13 100 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.136
+ $X2=0.999 $Y2=0.136
r147 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.136 $X2=0.999 $Y2=0.2025
r148 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.136
r149 5 66 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.135 $X2=0.837
+ $Y2=0.135
r150 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.2295
r151 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.0405 $X2=0.837 $Y2=0.135
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%QN 1 2 6 11 12 15 16 21 24 29 40 42 VSS
c14 44 VSS 0.00147594f $X=1.162 $Y=0.196
c15 42 VSS 6.36985e-19 $X=1.162 $Y=0.1355
c16 41 VSS 0.0040149f $X=1.162 $Y=0.122
c17 40 VSS 0.00181756f $X=1.166 $Y=0.149
c18 38 VSS 0.00144174f $X=1.162 $Y=0.225
c19 29 VSS 0.0196895f $X=1.153 $Y=0.234
c20 28 VSS 0.00635401f $X=1.134 $Y=0.036
c21 24 VSS 0.00903278f $X=1.026 $Y=0.036
c22 21 VSS 0.0196989f $X=1.153 $Y=0.036
c23 19 VSS 0.00662347f $X=1.132 $Y=0.2025
c24 15 VSS 0.00940513f $X=1.026 $Y=0.2025
c25 11 VSS 5.72268e-19 $X=1.043 $Y=0.2025
c26 9 VSS 2.69461e-19 $X=1.132 $Y=0.0675
c27 1 VSS 5.72268e-19 $X=1.043 $Y=0.0675
r28 43 44 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.167 $X2=1.162 $Y2=0.196
r29 41 42 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.122 $X2=1.162 $Y2=0.1355
r30 40 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.149 $X2=1.162 $Y2=0.167
r31 40 42 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.149 $X2=1.162 $Y2=0.1355
r32 38 44 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.225 $X2=1.162 $Y2=0.196
r33 37 41 5.22839 $w=1.8e-08 $l=7.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.045 $X2=1.162 $Y2=0.122
r34 31 35 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.234 $X2=1.134 $Y2=0.234
r35 29 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.153 $Y=0.234 $X2=1.162 $Y2=0.225
r36 29 35 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.153
+ $Y=0.234 $X2=1.134 $Y2=0.234
r37 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.134 $Y=0.036 $X2=1.134
+ $Y2=0.036
r38 23 27 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.036 $X2=1.134 $Y2=0.036
r39 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.036 $X2=1.026
+ $Y2=0.036
r40 21 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.153 $Y=0.036 $X2=1.162 $Y2=0.045
r41 21 27 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.153
+ $Y=0.036 $X2=1.134 $Y2=0.036
r42 19 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.134 $Y=0.234 $X2=1.134
+ $Y2=0.234
r43 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.117 $Y=0.2025 $X2=1.132 $Y2=0.2025
r44 15 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.234 $X2=1.026
+ $Y2=0.234
r45 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.2025 $X2=1.026 $Y2=0.2025
r46 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.043 $Y=0.2025 $X2=1.026 $Y2=0.2025
r47 9 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.134
+ $Y=0.0675 $X2=1.134 $Y2=0.036
r48 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.117
+ $Y=0.0675 $X2=1.132 $Y2=0.0675
r49 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.026
+ $Y=0.0675 $X2=1.026 $Y2=0.036
r50 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.009
+ $Y=0.0675 $X2=1.026 $Y2=0.0675
r51 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.043
+ $Y=0.0675 $X2=1.026 $Y2=0.0675
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%12 1 6 9 VSS
c6 9 VSS 0.0270172f $X=0.38 $Y=0.0675
c7 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c8 4 VSS 3.25039e-19 $X=0.322 $Y=0.0675
r9 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r10 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%13 1 6 9 VSS
c10 9 VSS 0.0209308f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.6182e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%14 1 6 9 VSS
c8 9 VSS 0.0191671f $X=0.758 $Y=0.0405
c9 6 VSS 3.14771e-19 $X=0.773 $Y=0.0405
c10 4 VSS 2.6194e-19 $X=0.7 $Y=0.0405
r11 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r12 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.7
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r13 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.685
+ $Y=0.0405 $X2=0.7 $Y2=0.0405
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%15 1 2 VSS
c0 1 VSS 0.00225696f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%16 1 2 VSS
c3 1 VSS 0.00231486f $X=0.341 $Y=0.2025
r4 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends

.subckt PM_DFFHQNX3_ASAP7_75T_SRAM%17 1 2 VSS
c0 1 VSS 0.00219822f $X=0.773 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2295 $X2=0.739 $Y2=0.2295
.ends


* END of "./DFFHQNx3_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DFFHQNx3_ASAP7_75t_SRAM  VSS VDD CLK D QN
* 
* QN	QN
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_12_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_4_M3_g N_12_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_15_M4_d N_6_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_15_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_10_M7_d N_6_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.611
+ $Y=0.027
M8 N_14_M8_d N_4_M8_g N_10_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M9 VSS N_9_M9_g N_14_M9_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_9_M10_d N_10_M10_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.027
M11 N_QN_M11_d N_10_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M12 N_QN_M12_d N_10_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.027
M13 N_QN_M13_d N_10_M13_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.027
M14 VDD N_CLK_M14_g N_4_M14_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M15 N_6_M15_d N_4_M15_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M16 N_16_M16_d N_D_M16_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M17 N_8_M17_d N_6_M17_g N_16_M17_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M18 N_13_M18_d N_4_M18_g N_8_M18_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M19 VDD N_7_M19_g N_13_M19_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M20 N_7_M20_d N_8_M20_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M21 N_10_M21_d N_4_M21_g N_7_M21_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.665 $Y=0.216
M22 N_17_M22_d N_6_M22_g N_10_M22_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.719 $Y=0.216
M23 VDD N_9_M23_g N_17_M23_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M24 N_9_M24_d N_10_M24_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.216
M25 N_QN_M25_d N_10_M25_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
M26 N_QN_M26_d N_10_M26_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.162
M27 N_QN_M27_d N_10_M27_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.162
*
* 
* .include "DFFHQNx3_ASAP7_75t_SRAM.pex.sp.DFFHQNX3_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DFFHQNx3_ASAP7_75t_SRAM.pex.sp.DFFHQNX3_ASAP7_75T_SRAM.pxi"
* File: DFFHQNx3_ASAP7_75t_SRAM.pex.sp.DFFHQNX3_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:24:53 2017
* 
x_PM_DFFHQNX3_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_13_p N_CLK_M14_g CLK
+ N_CLK_c_6_p VSS PM_DFFHQNX3_ASAP7_75T_SRAM%CLK
x_PM_DFFHQNX3_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M15_g N_4_M3_g N_4_c_43_p N_4_M18_g
+ N_4_M8_g N_4_c_48_p N_4_M21_g N_4_M0_s N_4_c_22_n N_4_M14_s N_4_c_23_n
+ N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_28_n N_4_c_29_n N_4_c_30_n
+ N_4_c_31_n N_4_c_40_p N_4_c_49_p N_4_c_37_p N_4_c_69_p N_4_c_33_n N_4_c_34_n
+ N_4_c_39_p N_4_c_51_p VSS PM_DFFHQNX3_ASAP7_75T_SRAM%4
x_PM_DFFHQNX3_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_99_n N_D_M16_g N_D_c_113_p D
+ N_D_c_101_n N_D_c_109_p N_D_c_102_n N_D_c_103_n VSS PM_DFFHQNX3_ASAP7_75T_SRAM%D
x_PM_DFFHQNX3_ASAP7_75T_SRAM%6 N_6_c_121_n N_6_M17_g N_6_M4_g N_6_M7_g N_6_c_171_p
+ N_6_c_125_n N_6_M22_g N_6_c_183_p N_6_c_126_n N_6_M1_d N_6_M15_d N_6_c_116_n
+ N_6_c_149_n N_6_c_132_n N_6_c_117_n N_6_c_150_n N_6_c_118_n N_6_c_135_n
+ N_6_c_136_n N_6_c_137_n N_6_c_138_n N_6_c_139_n N_6_c_119_n N_6_c_142_n
+ N_6_c_120_n N_6_c_143_n N_6_c_145_n N_6_c_188_p VSS PM_DFFHQNX3_ASAP7_75T_SRAM%6
x_PM_DFFHQNX3_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_244_p N_7_M19_g N_7_M7_s N_7_M6_d
+ N_7_c_228_n N_7_M20_d N_7_c_229_n N_7_M21_s N_7_c_231_n N_7_c_241_p
+ N_7_c_219_n N_7_c_220_n N_7_c_243_p N_7_c_260_p N_7_c_221_n N_7_c_246_p
+ N_7_c_222_n N_7_c_236_n N_7_c_237_n N_7_c_239_n N_7_c_223_n VSS
+ PM_DFFHQNX3_ASAP7_75T_SRAM%7
x_PM_DFFHQNX3_ASAP7_75T_SRAM%8 N_8_M6_g N_8_c_262_n N_8_M20_g N_8_M3_d N_8_M4_s
+ N_8_M17_d N_8_c_264_n N_8_M18_s N_8_c_310_p N_8_c_276_n N_8_c_265_n
+ N_8_c_311_p N_8_c_267_n N_8_c_283_n N_8_c_284_n N_8_c_268_n N_8_c_312_p
+ N_8_c_269_n N_8_c_286_n N_8_c_288_n N_8_c_302_n N_8_c_271_n N_8_c_303_n
+ N_8_c_272_n N_8_c_295_n N_8_c_273_n N_8_c_274_n N_8_c_275_n VSS
+ PM_DFFHQNX3_ASAP7_75T_SRAM%8
x_PM_DFFHQNX3_ASAP7_75T_SRAM%9 N_9_M9_g N_9_c_320_p N_9_M23_g N_9_M10_d N_9_M24_d
+ N_9_c_319_p N_9_c_331_p N_9_c_318_p N_9_c_323_p N_9_c_317_p N_9_c_327_p
+ N_9_c_329_p N_9_c_336_p N_9_c_328_p N_9_c_332_p N_9_c_322_p N_9_c_330_p
+ N_9_c_333_p VSS PM_DFFHQNX3_ASAP7_75T_SRAM%9
x_PM_DFFHQNX3_ASAP7_75T_SRAM%10 N_10_M10_g N_10_M24_g N_10_M11_g N_10_M25_g
+ N_10_M12_g N_10_M26_g N_10_M13_g N_10_c_387_p N_10_M27_g N_10_M8_s N_10_M7_d
+ N_10_c_338_n N_10_M22_s N_10_M21_d N_10_c_348_n N_10_c_370_n N_10_c_339_n
+ N_10_c_340_n N_10_c_401_p N_10_c_342_n N_10_c_362_n N_10_c_349_n N_10_c_343_n
+ N_10_c_350_n N_10_c_351_n N_10_c_375_n N_10_c_353_n N_10_c_376_n N_10_c_378_n
+ N_10_c_379_n N_10_c_380_n N_10_c_354_n N_10_c_355_n N_10_c_381_n N_10_c_344_n
+ N_10_c_386_n VSS PM_DFFHQNX3_ASAP7_75T_SRAM%10
x_PM_DFFHQNX3_ASAP7_75T_SRAM%QN N_QN_M12_d N_QN_M11_d N_QN_M13_d N_QN_M26_d
+ N_QN_M25_d N_QN_c_408_n N_QN_M27_d N_QN_c_404_n N_QN_c_412_n N_QN_c_405_n QN
+ N_QN_c_416_n VSS PM_DFFHQNX3_ASAP7_75T_SRAM%QN
x_PM_DFFHQNX3_ASAP7_75T_SRAM%12 N_12_M2_d N_12_M3_s N_12_c_418_n VSS
+ PM_DFFHQNX3_ASAP7_75T_SRAM%12
x_PM_DFFHQNX3_ASAP7_75T_SRAM%13 N_13_M18_d N_13_M19_s N_13_c_425_n VSS
+ PM_DFFHQNX3_ASAP7_75T_SRAM%13
x_PM_DFFHQNX3_ASAP7_75T_SRAM%14 N_14_M8_d N_14_M9_s N_14_c_434_n VSS
+ PM_DFFHQNX3_ASAP7_75T_SRAM%14
x_PM_DFFHQNX3_ASAP7_75T_SRAM%15 N_15_M5_s N_15_M4_d VSS PM_DFFHQNX3_ASAP7_75T_SRAM%15
x_PM_DFFHQNX3_ASAP7_75T_SRAM%16 N_16_M17_s N_16_M16_d VSS
+ PM_DFFHQNX3_ASAP7_75T_SRAM%16
x_PM_DFFHQNX3_ASAP7_75T_SRAM%17 N_17_M23_s N_17_M22_d VSS
+ PM_DFFHQNX3_ASAP7_75T_SRAM%17
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_22_n 3.57152e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 CLK N_4_c_23_n 0.00136255f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.144
cc_4 CLK N_4_c_24_n 2.75361e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.07
cc_5 CLK N_4_c_25_n 0.00136255f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.107
cc_6 N_CLK_c_6_p N_4_c_26_n 0.00145637f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2
cc_7 N_CLK_c_6_p N_4_c_27_n 2.75361e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2125
cc_8 CLK N_4_c_28_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_6_p N_4_c_29_n 5.03453e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_6_p N_4_c_30_n 0.00123168f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.153
cc_11 CLK N_4_c_31_n 4.93618e-19 $X=0.082 $Y=0.119 $X2=0.175 $Y2=0.153
cc_12 N_CLK_c_6_p N_4_c_31_n 0.00162391f $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_13 N_CLK_c_13_p N_4_c_33_n 0.00115059f $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.135
cc_14 CLK N_4_c_34_n 0.00174864f $X=0.082 $Y=0.119 $X2=0.151 $Y2=0.135
cc_15 N_CLK_c_6_p N_4_c_34_n 3.32041e-19 $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.135
cc_16 CLK N_6_c_116_n 6.37157e-19 $X=0.082 $Y=0.119 $X2=0.027 $Y2=0.234
cc_17 N_CLK_c_6_p N_6_c_117_n 6.45547e-19 $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.153
cc_18 N_CLK_c_6_p N_6_c_118_n 0.00125366f $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_19 N_CLK_c_6_p N_6_c_119_n 4.3806e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_20 CLK N_6_c_120_n 0.00137619f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.153
cc_21 N_4_M3_g N_D_M2_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_22 N_4_c_37_p N_D_c_99_n 2.91747e-19 $X=0.527 $Y=0.153 $X2=0.081 $Y2=0.135
cc_23 N_4_c_33_n N_D_c_99_n 2.1478e-19 $X=0.151 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_4_c_39_p N_D_c_101_n 2.3983e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_25 N_4_c_40_p N_D_c_102_n 8.99815e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_26 N_4_c_40_p N_D_c_103_n 8.75229e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_27 N_4_M3_g N_6_c_121_n 0.00355599f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_28 N_4_c_43_p N_6_c_121_n 0.00126153f $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.054
cc_29 N_4_M3_g N_6_M4_g 0.00355599f $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_4_M8_g N_6_M7_g 0.00355599f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_31 N_4_M8_g N_6_c_125_n 0.00355599f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_32 N_4_M8_g N_6_c_126_n 0.00250257f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_33 N_4_c_48_p N_6_c_126_n 0.00180656f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_34 N_4_c_49_p N_6_c_126_n 6.4075e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_35 N_4_c_37_p N_6_c_126_n 0.00187561f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_36 N_4_c_51_p N_6_c_126_n 0.00123876f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_34_n N_6_c_116_n 2.97444e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_31_n N_6_c_132_n 2.38327e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_34_n N_6_c_117_n 2.85146e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_40_p N_6_c_118_n 2.46239e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_41 N_4_c_31_n N_6_c_135_n 2.31165e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_42 N_4_c_39_p N_6_c_136_n 9.24693e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_43 N_4_c_37_p N_6_c_137_n 3.67557e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_44 N_4_c_37_p N_6_c_138_n 8.06691e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_45 N_4_c_37_p N_6_c_139_n 2.46239e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_46 N_4_c_40_p N_6_c_119_n 0.0299327f $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_39_p N_6_c_119_n 2.98936e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_48 N_4_c_37_p N_6_c_142_n 2.81476e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_49 N_4_c_40_p N_6_c_143_n 8.79704e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_50 N_4_c_34_n N_6_c_143_n 0.00524677f $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_51 N_4_c_37_p N_6_c_145_n 9.92294e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_52 N_4_c_39_p N_6_c_145_n 5.5596e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_53 N_4_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_54 N_4_c_69_p N_7_c_219_n 3.42573e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_55 N_4_c_69_p N_7_c_220_n 5.29207e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_56 N_4_c_51_p N_7_c_221_n 0.00318218f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_57 N_4_c_49_p N_7_c_222_n 0.00115177f $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_58 N_4_c_49_p N_7_c_223_n 3.42573e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_59 N_4_M8_g N_8_M6_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_60 N_4_c_48_p N_8_c_262_n 3.88499e-19 $X=0.675 $Y=0.135 $X2=0.081 $Y2=0.135
cc_61 N_4_c_69_p N_8_c_262_n 3.00379e-19 $X=0.601 $Y=0.153 $X2=0.081 $Y2=0.135
cc_62 N_4_c_39_p N_8_c_264_n 2.36208e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_63 N_4_M3_g N_8_c_265_n 3.49806e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_4_c_39_p N_8_c_265_n 3.83282e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_65 N_4_c_39_p N_8_c_267_n 7.25941e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_66 N_4_c_39_p N_8_c_268_n 7.25941e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_67 N_4_c_37_p N_8_c_269_n 0.00118282f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_68 N_4_c_39_p N_8_c_269_n 8.1935e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_69 N_4_c_37_p N_8_c_271_n 0.00132871f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_70 N_4_c_69_p N_8_c_272_n 0.00132871f $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_71 N_4_c_37_p N_8_c_273_n 2.54113e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_72 N_4_c_37_p N_8_c_274_n 3.92135e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_73 N_4_c_39_p N_8_c_275_n 7.25941e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_74 N_4_M8_g N_9_M9_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_75 N_4_c_49_p N_10_c_338_n 2.24654e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_76 N_4_c_49_p N_10_c_339_n 5.06919e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_77 N_4_M8_g N_10_c_340_n 3.47752e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_78 N_4_c_51_p N_10_c_340_n 5.72565e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_79 N_4_c_49_p N_10_c_342_n 2.46558e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_80 N_4_c_51_p N_10_c_343_n 0.00319993f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_81 N_4_c_49_p N_10_c_344_n 2.9112e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_82 N_4_c_37_p N_12_c_418_n 3.46326e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_83 N_D_M2_g N_6_c_121_n 0.00341068f $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_84 N_D_c_99_n N_6_c_121_n 0.00114686f $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_85 D N_6_c_149_n 0.00215667f $X=0.244 $Y=0.082 $X2=0.0505 $Y2=0.234
cc_86 N_D_c_103_n N_6_c_150_n 0.00215667f $X=0.243 $Y=0.135 $X2=0.405 $Y2=0.153
cc_87 N_D_c_103_n N_6_c_118_n 0.00225008f $X=0.243 $Y=0.135 $X2=0.175 $Y2=0.153
cc_88 N_D_c_109_p N_6_c_137_n 0.00127755f $X=0.281 $Y=0.135 $X2=0.151 $Y2=0.135
cc_89 N_D_c_99_n N_6_c_119_n 2.11668e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_90 N_D_c_103_n N_6_c_119_n 0.00122387f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_91 D N_6_c_120_n 0.00215667f $X=0.244 $Y=0.082 $X2=0.018 $Y2=0.153
cc_92 N_D_c_113_p N_6_c_143_n 0.00215667f $X=0.243 $Y=0.126 $X2=0 $Y2=0
cc_93 N_D_c_103_n N_6_c_145_n 0.00120973f $X=0.243 $Y=0.135 $X2=0.027 $Y2=0.153
cc_94 N_D_c_103_n N_8_c_276_n 2.80198e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_95 N_6_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_96 N_6_M7_g N_7_M5_g 2.13359e-19 $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_97 N_6_c_126_n N_7_M5_g 0.00205997f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_98 N_6_c_142_n N_7_M5_g 3.15189e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_99 N_6_c_126_n N_7_c_228_n 6.55731e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_100 N_6_c_126_n N_7_c_229_n 2.12581e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_101 N_6_c_126_n N_7_M21_s 2.50995e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_102 N_6_M7_g N_7_c_231_n 0.00200065f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_103 N_6_c_126_n N_7_c_231_n 0.00312129f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_104 N_6_c_126_n N_7_c_220_n 3.41745e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_105 N_6_M7_g N_7_c_221_n 3.41702e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_106 N_6_M7_g N_7_c_222_n 2.26424e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_107 N_6_c_142_n N_7_c_236_n 5.75704e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_108 N_6_c_171_p N_7_c_237_n 0.00195059f $X=0.621 $Y=0.178 $X2=0 $Y2=0
cc_109 N_6_c_126_n N_7_c_237_n 0.00191847f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_110 N_6_M7_g N_7_c_239_n 3.8308e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_111 N_6_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_112 N_6_M7_g N_8_M6_g 0.00341068f $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_113 N_6_c_126_n N_8_M6_g 0.00302156f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_114 N_6_c_119_n N_8_c_264_n 3.12535e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_115 N_6_c_145_n N_8_c_264_n 8.9852e-19 $X=0.324 $Y=0.167 $X2=0 $Y2=0
cc_116 N_6_c_119_n N_8_c_276_n 0.0015935f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_117 N_6_M4_g N_8_c_283_n 3.68551e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_118 N_6_M4_g N_8_c_284_n 2.06635e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_119 N_6_M4_g N_8_c_269_n 2.27069e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_120 N_6_c_183_p N_8_c_286_n 4.73369e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_121 N_6_c_142_n N_8_c_286_n 0.00174159f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_122 N_6_c_183_p N_8_c_288_n 0.00171407f $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_123 N_6_c_126_n N_8_c_288_n 5.88593e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_124 N_6_c_119_n N_8_c_288_n 0.00104904f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_125 N_6_c_188_p N_8_c_288_n 2.15173e-19 $X=0.324 $Y=0.178 $X2=0 $Y2=0
cc_126 N_6_c_126_n N_8_c_271_n 8.16411e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_127 N_6_c_126_n N_8_c_272_n 3.32592e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_128 N_6_c_142_n N_8_c_272_n 8.9822e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_129 N_6_c_126_n N_8_c_295_n 4.02972e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_130 N_6_c_125_n N_9_M9_g 0.00341068f $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_131 N_6_c_125_n N_10_M10_g 2.13359e-19 $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_132 N_6_c_126_n N_10_c_338_n 8.27829e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_133 N_6_c_126_n N_10_M22_s 3.37661e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_134 N_6_c_126_n N_10_c_348_n 0.00145548f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_135 N_6_c_125_n N_10_c_349_n 3.03386e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_136 N_6_c_125_n N_10_c_350_n 2.58526e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_137 N_6_c_125_n N_10_c_351_n 0.00228871f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_138 N_6_c_126_n N_10_c_351_n 7.89371e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_139 N_6_c_125_n N_10_c_353_n 4.55487e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_140 N_6_c_126_n N_10_c_354_n 4.54272e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_141 N_6_c_125_n N_10_c_355_n 5.68093e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_142 N_6_c_126_n N_10_c_355_n 2.2968e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_143 N_6_c_121_n N_12_c_418_n 0.00514294f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_144 N_6_c_137_n N_12_c_418_n 0.00114179f $X=0.333 $Y=0.135 $X2=0 $Y2=0
cc_145 N_6_c_126_n N_13_M19_s 2.36286e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.216
cc_146 N_6_M4_g N_13_c_425_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_147 N_6_c_183_p N_13_c_425_n 5.41258e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_148 N_6_c_126_n N_13_c_425_n 0.00230928f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_149 N_6_c_119_n N_13_c_425_n 7.09553e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_150 N_6_c_125_n N_14_c_434_n 0.00198387f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_151 N_6_c_126_n N_14_c_434_n 4.51352e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_152 N_6_c_139_n N_16_M17_s 8.59575e-19 $X=0.324 $Y=0.189 $X2=0.081 $Y2=0.054
cc_153 N_6_c_145_n N_16_M17_s 2.57402e-19 $X=0.324 $Y=0.167 $X2=0.081 $Y2=0.054
cc_154 N_6_c_188_p N_16_M17_s 2.18007e-19 $X=0.324 $Y=0.178 $X2=0.081 $Y2=0.054
cc_155 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_156 N_7_c_241_p N_8_M6_g 3.87418e-19 $X=0.576 $Y=0.09 $X2=0.135 $Y2=0.054
cc_157 N_7_c_221_n N_8_c_262_n 2.20449e-19 $X=0.621 $Y=0.122 $X2=0.135 $Y2=0.135
cc_158 N_7_c_243_p N_8_c_283_n 3.63506e-19 $X=0.594 $Y=0.054 $X2=0.018 $Y2=0.107
cc_159 N_7_c_244_p N_8_c_284_n 3.19692e-19 $X=0.513 $Y=0.09 $X2=0.018 $Y2=0.162
cc_160 N_7_c_241_p N_8_c_284_n 0.00114151f $X=0.576 $Y=0.09 $X2=0.018 $Y2=0.162
cc_161 N_7_c_246_p N_8_c_302_n 7.39815e-19 $X=0.621 $Y=0.14 $X2=0.027 $Y2=0.234
cc_162 N_7_c_241_p N_8_c_303_n 0.0047777f $X=0.576 $Y=0.09 $X2=0.054 $Y2=0.234
cc_163 N_7_M5_g N_8_c_272_n 3.12986e-19 $X=0.513 $Y=0.0405 $X2=0.047 $Y2=0.234
cc_164 N_7_c_244_p N_8_c_273_n 5.2508e-19 $X=0.513 $Y=0.09 $X2=0.033 $Y2=0.153
cc_165 N_7_c_228_n N_10_c_338_n 0.0027803f $X=0.594 $Y=0.0405 $X2=0.018 $Y2=0.07
cc_166 N_7_c_243_p N_10_c_338_n 3.72596e-19 $X=0.594 $Y=0.054 $X2=0.018 $Y2=0.07
cc_167 N_7_c_239_n N_10_c_338_n 3.30531e-19 $X=0.621 $Y=0.09 $X2=0.018 $Y2=0.07
cc_168 N_7_c_231_n N_10_c_348_n 0.00220898f $X=0.65 $Y=0.2295 $X2=0.018
+ $Y2=0.2125
cc_169 N_7_c_228_n N_10_c_339_n 5.23227e-19 $X=0.594 $Y=0.0405 $X2=0.0505
+ $Y2=0.036
cc_170 N_7_c_243_p N_10_c_362_n 2.3746e-19 $X=0.594 $Y=0.054 $X2=0.047 $Y2=0.234
cc_171 N_7_c_239_n N_10_c_349_n 4.46294e-19 $X=0.621 $Y=0.09 $X2=0.0505
+ $Y2=0.234
cc_172 N_7_c_237_n N_10_c_351_n 4.46294e-19 $X=0.621 $Y=0.203 $X2=0.033
+ $Y2=0.153
cc_173 N_7_c_231_n N_10_c_354_n 3.64147e-19 $X=0.65 $Y=0.2295 $X2=0.405
+ $Y2=0.135
cc_174 N_7_c_220_n N_10_c_354_n 4.68959e-19 $X=0.612 $Y=0.234 $X2=0.405
+ $Y2=0.135
cc_175 N_7_c_260_p N_10_c_355_n 4.46294e-19 $X=0.621 $Y=0.101 $X2=0 $Y2=0
cc_176 N_8_c_264_n N_12_c_418_n 0.00119486f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_177 N_8_c_273_n N_12_c_418_n 0.00390673f $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_178 N_8_c_274_n N_12_c_418_n 5.36233e-19 $X=0.45 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_179 N_8_c_264_n N_13_c_425_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_180 N_8_c_310_p N_13_c_425_n 0.00209454f $X=0.45 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_181 N_8_c_311_p N_13_c_425_n 0.0013184f $X=0.434 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_182 N_8_c_312_p N_13_c_425_n 0.00119522f $X=0.459 $Y=0.225 $X2=0.405
+ $Y2=0.0675
cc_183 N_8_c_273_n N_13_c_425_n 5.72158e-19 $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_184 N_9_M9_g N_10_M10_g 0.00268443f $X=0.783 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_185 N_9_c_317_p N_10_M10_g 3.74489e-19 $X=0.846 $Y=0.036 $X2=0.135 $Y2=0.054
cc_186 N_9_c_318_p N_10_c_370_n 0.00141609f $X=0.792 $Y=0.036 $X2=0.027
+ $Y2=0.036
cc_187 N_9_c_319_p N_10_c_362_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.047
+ $Y2=0.234
cc_188 N_9_c_320_p N_10_c_349_n 3.34766e-19 $X=0.783 $Y=0.1055 $X2=0.0505
+ $Y2=0.234
cc_189 N_9_c_319_p N_10_c_349_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.0505
+ $Y2=0.234
cc_190 N_9_c_322_p N_10_c_351_n 2.41112e-19 $X=0.945 $Y=0.225 $X2=0.033
+ $Y2=0.153
cc_191 N_9_c_323_p N_10_c_375_n 2.6154e-19 $X=0.828 $Y=0.036 $X2=0 $Y2=0
cc_192 N_9_M9_g N_10_c_376_n 6.3699e-19 $X=0.783 $Y=0.0405 $X2=0.151 $Y2=0.153
cc_193 N_9_c_319_p N_10_c_376_n 9.10342e-19 $X=0.783 $Y=0.105 $X2=0.151
+ $Y2=0.153
cc_194 N_9_c_317_p N_10_c_378_n 4.40983e-19 $X=0.846 $Y=0.036 $X2=0.405
+ $Y2=0.153
cc_195 N_9_c_327_p N_10_c_379_n 5.13693e-19 $X=0.882 $Y=0.036 $X2=0.601
+ $Y2=0.153
cc_196 N_9_c_328_p N_10_c_380_n 0.00149072f $X=0.9 $Y=0.234 $X2=0 $Y2=0
cc_197 N_9_c_329_p N_10_c_381_n 4.52584e-19 $X=0.9 $Y=0.036 $X2=0 $Y2=0
cc_198 N_9_c_330_p N_10_c_381_n 0.00280794f $X=0.945 $Y=0.122 $X2=0 $Y2=0
cc_199 N_9_c_331_p N_10_c_344_n 2.40515e-19 $X=0.936 $Y=0.036 $X2=0 $Y2=0
cc_200 N_9_c_332_p N_10_c_344_n 7.44774e-19 $X=0.918 $Y=0.234 $X2=0 $Y2=0
cc_201 N_9_c_333_p N_10_c_344_n 8.84468e-19 $X=0.945 $Y=0.167 $X2=0 $Y2=0
cc_202 N_9_c_333_p N_10_c_386_n 0.00213033f $X=0.945 $Y=0.167 $X2=0 $Y2=0
cc_203 N_9_c_331_p N_QN_c_404_n 4.76361e-19 $X=0.936 $Y=0.036 $X2=0.675
+ $Y2=0.135
cc_204 N_9_c_336_p N_QN_c_405_n 4.61952e-19 $X=0.936 $Y=0.234 $X2=0 $Y2=0
cc_205 N_9_c_318_p N_14_c_434_n 7.33799e-19 $X=0.792 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_206 N_10_c_387_p N_QN_M12_d 3.7444e-19 $X=1.107 $Y=0.136 $X2=0.135 $Y2=0.054
cc_207 N_10_c_387_p N_QN_M26_d 3.85232e-19 $X=1.107 $Y=0.136 $X2=0 $Y2=0
cc_208 N_10_c_387_p N_QN_c_408_n 8.43851e-19 $X=1.107 $Y=0.136 $X2=0.405
+ $Y2=0.2295
cc_209 N_10_M12_g N_QN_c_404_n 4.61823e-19 $X=1.053 $Y=0.0675 $X2=0.675
+ $Y2=0.135
cc_210 N_10_M13_g N_QN_c_404_n 4.61823e-19 $X=1.107 $Y=0.0675 $X2=0.675
+ $Y2=0.135
cc_211 N_10_c_387_p N_QN_c_404_n 0.00131663f $X=1.107 $Y=0.136 $X2=0.675
+ $Y2=0.135
cc_212 N_10_c_387_p N_QN_c_412_n 7.60428e-19 $X=1.107 $Y=0.136 $X2=0 $Y2=0
cc_213 N_10_M12_g N_QN_c_405_n 4.56718e-19 $X=1.053 $Y=0.0675 $X2=0 $Y2=0
cc_214 N_10_M13_g N_QN_c_405_n 4.56718e-19 $X=1.107 $Y=0.0675 $X2=0 $Y2=0
cc_215 N_10_c_387_p N_QN_c_405_n 0.00134222f $X=1.107 $Y=0.136 $X2=0 $Y2=0
cc_216 N_10_c_387_p N_QN_c_416_n 3.48867e-19 $X=1.107 $Y=0.136 $X2=0.018
+ $Y2=0.2125
cc_217 N_10_c_386_n N_QN_c_416_n 2.87084e-19 $X=0.999 $Y=0.136 $X2=0.018
+ $Y2=0.2125
cc_218 N_10_c_338_n N_14_c_434_n 0.00182708f $X=0.648 $Y=0.0405 $X2=0.405
+ $Y2=0.0675
cc_219 N_10_c_370_n N_14_c_434_n 0.0020512f $X=0.72 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_220 N_10_c_401_p N_14_c_434_n 0.00131745f $X=0.704 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_221 N_10_c_362_n N_14_c_434_n 0.00103589f $X=0.729 $Y=0.081 $X2=0.405
+ $Y2=0.0675
cc_222 N_10_c_353_n N_14_c_434_n 4.02739e-19 $X=0.774 $Y=0.162 $X2=0.405
+ $Y2=0.0675

* END of "./DFFHQNx3_ASAP7_75t_SRAM.pex.sp.DFFHQNX3_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DFFHQx4_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:25:16 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DFFHQx4_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DFFHQx4_ASAP7_75t_SRAM.pex.sp.pex"
* File: DFFHQx4_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:25:16 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DFFHQX4_ASAP7_75T_SRAM%CLK 2 5 7 12 14 VSS
c20 14 VSS 0.00665223f $X=0.081 $Y=0.135
c21 12 VSS 0.00671818f $X=0.082 $Y=0.119
c22 5 VSS 0.00212887f $X=0.081 $Y=0.135
c23 2 VSS 0.0629f $X=0.081 $Y=0.054
r24 12 14 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.135
r25 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r26 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r27 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%4 2 7 10 13 15 18 21 23 25 28 30 36 37 38 41 42
+ 45 52 59 67 68 70 72 73 78 79 83 88 VSS
c80 114 VSS 1.06551e-19 $X=0.03 $Y=0.153
c81 113 VSS 6.89947e-19 $X=0.027 $Y=0.153
c82 88 VSS 0.00102973f $X=0.675 $Y=0.135
c83 83 VSS 8.77298e-19 $X=0.405 $Y=0.135
c84 79 VSS 0.00121012f $X=0.151 $Y=0.135
c85 78 VSS 0.00388356f $X=0.151 $Y=0.135
c86 73 VSS 0.00260015f $X=0.601 $Y=0.153
c87 72 VSS 0.00550417f $X=0.527 $Y=0.153
c88 70 VSS 0.0040358f $X=0.675 $Y=0.153
c89 68 VSS 0.00327616f $X=0.29 $Y=0.153
c90 67 VSS 0.00599408f $X=0.175 $Y=0.153
c91 59 VSS 6.74612e-19 $X=0.033 $Y=0.153
c92 55 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c93 54 VSS 0.00180216f $X=0.047 $Y=0.234
c94 52 VSS 0.00250119f $X=0.054 $Y=0.234
c95 50 VSS 0.00305101f $X=0.027 $Y=0.234
c96 48 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c97 47 VSS 0.00199699f $X=0.047 $Y=0.036
c98 45 VSS 0.00250119f $X=0.054 $Y=0.036
c99 43 VSS 0.00305101f $X=0.027 $Y=0.036
c100 42 VSS 4.88707e-19 $X=0.018 $Y=0.2125
c101 41 VSS 0.00180713f $X=0.018 $Y=0.2
c102 40 VSS 4.69158e-19 $X=0.018 $Y=0.225
c103 38 VSS 0.00173342f $X=0.018 $Y=0.107
c104 37 VSS 9.57865e-19 $X=0.018 $Y=0.07
c105 36 VSS 0.00172854f $X=0.018 $Y=0.144
c106 33 VSS 0.00565775f $X=0.056 $Y=0.216
c107 30 VSS 2.98509e-19 $X=0.071 $Y=0.216
c108 28 VSS 0.00554224f $X=0.056 $Y=0.054
c109 25 VSS 2.98509e-19 $X=0.071 $Y=0.054
c110 21 VSS 0.00207437f $X=0.675 $Y=0.135
c111 18 VSS 0.0585656f $X=0.675 $Y=0.0405
c112 13 VSS 0.00211542f $X=0.405 $Y=0.135
c113 10 VSS 0.058827f $X=0.405 $Y=0.0675
c114 2 VSS 0.0628024f $X=0.135 $Y=0.054
r115 113 114 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r116 110 113 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r117 78 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.151 $Y=0.135 $X2=0.151
+ $Y2=0.135
r118 72 73 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.601 $Y2=0.153
r119 70 73 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.675
+ $Y=0.153 $X2=0.601 $Y2=0.153
r120 70 88 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.675 $Y=0.153 $X2=0.675
+ $Y2=0.153
r121 67 68 7.80864 $w=1.8e-08 $l=1.15e-07 $layer=M2 $thickness=3.6e-08 $X=0.175
+ $Y=0.153 $X2=0.29 $Y2=0.153
r122 65 72 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.527 $Y2=0.153
r123 65 68 7.80864 $w=1.8e-08 $l=1.15e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.29 $Y2=0.153
r124 65 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r125 62 67 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.151
+ $Y=0.153 $X2=0.175 $Y2=0.153
r126 62 79 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.151 $Y=0.153 $X2=0.151
+ $Y2=0.153
r127 59 114 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r128 58 62 8.01235 $w=1.8e-08 $l=1.18e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.151 $Y2=0.153
r129 58 59 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r130 54 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r131 52 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r132 50 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r133 47 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r134 45 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r135 43 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r136 41 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r137 40 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r138 40 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r139 39 110 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r140 39 41 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.2
r141 37 38 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.107
r142 36 110 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r143 36 38 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.107
r144 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r145 35 37 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r146 33 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r147 30 33 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r148 28 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r149 25 28 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r150 21 88 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.135 $X2=0.675
+ $Y2=0.135
r151 21 23 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2295
r152 18 21 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.135
r153 13 83 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r154 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2295
r155 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r156 5 78 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.151 $Y2=0.135
r157 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r158 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%D 2 5 7 10 12 14 21 23 28 VSS
c18 28 VSS 0.00931082f $X=0.243 $Y=0.135
c19 24 VSS 2.45662e-20 $X=0.276 $Y=0.135
c20 23 VSS 0.00111822f $X=0.271 $Y=0.135
c21 21 VSS 2.56376e-19 $X=0.281 $Y=0.135
c22 14 VSS 2.7811e-19 $X=0.243 $Y=0.116
c23 12 VSS 0.00925957f $X=0.244 $Y=0.082
c24 10 VSS 2.38113e-19 $X=0.243 $Y=0.126
c25 5 VSS 0.00529812f $X=0.297 $Y=0.135
c26 2 VSS 0.0630392f $X=0.297 $Y=0.0675
r27 23 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.271
+ $Y=0.135 $X2=0.276 $Y2=0.135
r28 21 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.281
+ $Y=0.135 $X2=0.276 $Y2=0.135
r29 21 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.281 $Y=0.135 $X2=0.281
+ $Y2=0.135
r30 19 28 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.243 $Y2=0.135
r31 19 23 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.271 $Y2=0.135
r32 13 14 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.106 $X2=0.243 $Y2=0.116
r33 12 13 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.082 $X2=0.243 $Y2=0.106
r34 10 28 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.135
r35 10 14 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.116
r36 5 22 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.281 $Y2=0.135
r37 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r38 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%6 2 5 8 14 17 20 23 28 35 39 44 50 55 57 61 66 67
+ 68 75 77 78 87 89 105 110 111 113 114 VSS
c101 114 VSS 2.23151e-19 $X=0.324 $Y=0.178
c102 113 VSS 4.08645e-19 $X=0.324 $Y=0.167
c103 111 VSS 7.77947e-19 $X=0.189 $Y=0.167
c104 110 VSS 9.60988e-19 $X=0.189 $Y=0.106
c105 105 VSS 6.81413e-19 $X=0.513 $Y=0.18
c106 89 VSS 0.0113851f $X=0.513 $Y=0.189
c107 87 VSS 0.00137981f $X=0.324 $Y=0.189
c108 78 VSS 4.01595e-19 $X=0.342 $Y=0.135
c109 77 VSS 5.2076e-19 $X=0.333 $Y=0.135
c110 75 VSS 7.41013e-19 $X=0.351 $Y=0.135
c111 68 VSS 0.00169555f $X=0.18 $Y=0.234
c112 67 VSS 9.43175e-19 $X=0.189 $Y=0.225
c113 66 VSS 0.00196236f $X=0.189 $Y=0.234
c114 61 VSS 0.00196921f $X=0.162 $Y=0.234
c115 57 VSS 0.00170883f $X=0.18 $Y=0.036
c116 55 VSS 0.00196236f $X=0.189 $Y=0.036
c117 50 VSS 0.00193426f $X=0.162 $Y=0.036
c118 47 VSS 0.00754879f $X=0.16 $Y=0.216
c119 42 VSS 0.00764528f $X=0.16 $Y=0.054
c120 35 VSS 0.0610442f $X=0.725 $Y=0.178
c121 28 VSS 0.00134228f $X=0.464 $Y=0.178
c122 20 VSS 0.0613962f $X=0.729 $Y=0.178
c123 17 VSS 1.08457e-19 $X=0.621 $Y=0.178
c124 14 VSS 0.0600374f $X=0.621 $Y=0.0405
c125 8 VSS 0.0601849f $X=0.459 $Y=0.0405
c126 2 VSS 0.0623471f $X=0.351 $Y=0.135
r127 113 114 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.324 $Y=0.167 $X2=0.324 $Y2=0.178
r128 110 111 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.106 $X2=0.189 $Y2=0.167
r129 104 105 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r130 89 105 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r131 87 114 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.189 $X2=0.324 $Y2=0.178
r132 86 89 12.8333 $w=1.8e-08 $l=1.89e-07 $layer=M2 $thickness=3.6e-08 $X=0.324
+ $Y=0.189 $X2=0.513 $Y2=0.189
r133 86 87 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.324 $Y=0.189 $X2=0.324
+ $Y2=0.189
r134 83 111 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.167
r135 82 86 9.16667 $w=1.8e-08 $l=1.35e-07 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.324 $Y2=0.189
r136 82 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.189 $X2=0.189
+ $Y2=0.189
r137 77 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.135 $X2=0.342 $Y2=0.135
r138 75 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.342 $Y2=0.135
r139 72 113 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.144 $X2=0.324 $Y2=0.167
r140 71 77 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.135 $X2=0.333 $Y2=0.135
r141 71 72 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.135 $X2=0.324 $Y2=0.144
r142 68 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r143 67 83 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.189
r144 66 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r145 66 67 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.189 $Y2=0.225
r146 61 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r147 57 58 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r148 56 110 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.106
r149 55 58 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r150 55 56 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r151 50 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r152 47 61 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r153 44 47 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r154 42 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r155 39 42 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r156 28 104 39.0385 $w=2.6e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.178 $X2=0.513 $Y2=0.178
r157 20 35 3.07692 $w=2.6e-08 $l=4e-09 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.178 $X2=0.725 $Y2=0.178
r158 20 23 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.178 $X2=0.729 $Y2=0.2295
r159 17 35 82.8571 $w=2.6e-08 $l=1.04e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.725 $Y2=0.178
r160 17 104 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.513 $Y2=0.178
r161 14 17 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0405 $X2=0.621 $Y2=0.178
r162 11 28 3.84615 $w=2.6e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.178 $X2=0.464 $Y2=0.178
r163 8 11 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.178
r164 2 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r165 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%7 2 5 7 9 10 13 14 17 19 22 29 30 31 33 40 45 46
+ 47 48 49 50 54 55 VSS
c43 56 VSS 3.52511e-19 $X=0.612 $Y=0.09
c44 55 VSS 1.80704e-19 $X=0.603 $Y=0.09
c45 54 VSS 5.96246e-19 $X=0.621 $Y=0.09
c46 51 VSS 6.85462e-19 $X=0.621 $Y=0.224
c47 50 VSS 4.95788e-19 $X=0.621 $Y=0.203
c48 49 VSS 1.19762e-19 $X=0.621 $Y=0.167
c49 48 VSS 3.47205e-19 $X=0.621 $Y=0.165
c50 47 VSS 2.82671e-19 $X=0.621 $Y=0.14
c51 46 VSS 4.86366e-19 $X=0.621 $Y=0.122
c52 45 VSS 1.45036e-19 $X=0.621 $Y=0.101
c53 40 VSS 0.00113884f $X=0.594 $Y=0.054
c54 33 VSS 0.00266679f $X=0.594 $Y=0.234
c55 31 VSS 0.00427836f $X=0.612 $Y=0.234
c56 30 VSS 1.97343e-19 $X=0.583 $Y=0.09
c57 29 VSS 0.00268203f $X=0.581 $Y=0.09
c58 24 VSS 4.90193e-20 $X=0.585 $Y=0.09
c59 22 VSS 0.0185872f $X=0.65 $Y=0.2295
c60 19 VSS 3.14771e-19 $X=0.665 $Y=0.2295
c61 17 VSS 2.5391e-19 $X=0.592 $Y=0.2295
c62 13 VSS 0.00396424f $X=0.594 $Y=0.0405
c63 9 VSS 6.29543e-19 $X=0.611 $Y=0.0405
c64 5 VSS 0.00255452f $X=0.513 $Y=0.09
c65 2 VSS 0.0583002f $X=0.513 $Y=0.0405
r66 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.603
+ $Y=0.09 $X2=0.612 $Y2=0.09
r67 54 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.612 $Y2=0.09
r68 53 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.09 $X2=0.603 $Y2=0.09
r69 51 52 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.224 $X2=0.621 $Y2=0.2245
r70 50 51 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.224
r71 49 50 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.203
r72 48 49 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.167
r73 47 48 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r74 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r75 45 46 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.101 $X2=0.621 $Y2=0.122
r76 44 52 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.2245
r77 43 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.09
r78 43 45 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.101
r79 38 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.09
r80 38 40 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.054
r81 31 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r82 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r83 29 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.581
+ $Y=0.09 $X2=0.583 $Y2=0.09
r84 26 29 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.09 $X2=0.581 $Y2=0.09
r85 24 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.594 $Y2=0.09
r86 24 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.583 $Y2=0.09
r87 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2295 $X2=0.65 $Y2=0.2295
r88 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.592
+ $Y=0.2295 $X2=0.65 $Y2=0.2295
r89 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r90 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r91 13 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.054 $X2=0.594
+ $Y2=0.054
r92 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.594 $Y2=0.0405
r93 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0405 $X2=0.594 $Y2=0.0405
r94 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.09 $X2=0.513
+ $Y2=0.09
r95 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.09 $X2=0.513 $Y2=0.2295
r96 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.09
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%8 2 5 7 9 14 17 21 22 25 27 33 35 37 38 39 41 43
+ 44 45 46 50 52 53 54 55 60 63 66 VSS
c54 66 VSS 2.86012e-19 $X=0.459 $Y=0.131
c55 63 VSS 0.00343707f $X=0.45 $Y=0.036
c56 62 VSS 0.0025237f $X=0.459 $Y=0.036
c57 60 VSS 0.00424264f $X=0.432 $Y=0.036
c58 55 VSS 4.23511e-19 $X=0.5445 $Y=0.131
c59 54 VSS 3.49205e-20 $X=0.522 $Y=0.131
c60 53 VSS 2.0008e-19 $X=0.504 $Y=0.131
c61 52 VSS 0.00133205f $X=0.496 $Y=0.131
c62 50 VSS 5.30081e-19 $X=0.567 $Y=0.131
c63 47 VSS 4.30827e-19 $X=0.459 $Y=0.214
c64 46 VSS 2.06877e-19 $X=0.459 $Y=0.203
c65 45 VSS 6.09344e-21 $X=0.459 $Y=0.167
c66 44 VSS 2.1141e-19 $X=0.459 $Y=0.165
c67 43 VSS 2.51143e-19 $X=0.459 $Y=0.225
c68 41 VSS 3.66085e-19 $X=0.459 $Y=0.114
c69 40 VSS 3.44034e-19 $X=0.459 $Y=0.106
c70 38 VSS 7.88894e-19 $X=0.459 $Y=0.081
c71 37 VSS 2.0833e-19 $X=0.459 $Y=0.122
c72 35 VSS 0.00142907f $X=0.434 $Y=0.234
c73 34 VSS 3.33033e-19 $X=0.418 $Y=0.234
c74 33 VSS 0.00146362f $X=0.414 $Y=0.234
c75 32 VSS 0.00227837f $X=0.396 $Y=0.234
c76 27 VSS 0.00148441f $X=0.378 $Y=0.234
c77 25 VSS 0.00389542f $X=0.45 $Y=0.234
c78 24 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c79 21 VSS 0.00449633f $X=0.378 $Y=0.2025
c80 18 VSS 1.15515e-19 $X=0.3735 $Y=0.216
c81 16 VSS 5.70081e-19 $X=0.432 $Y=0.0405
c82 10 VSS 7.61325e-20 $X=0.4275 $Y=0.054
c83 5 VSS 0.00216437f $X=0.567 $Y=0.1305
c84 2 VSS 0.0591864f $X=0.567 $Y=0.0405
r85 63 64 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r86 62 64 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r87 59 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r88 59 60 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r89 54 55 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r90 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r91 52 53 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.496
+ $Y=0.131 $X2=0.504 $Y2=0.131
r92 50 55 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r93 48 66 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r94 48 52 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.496 $Y2=0.131
r95 46 47 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.203 $X2=0.459 $Y2=0.214
r96 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.167 $X2=0.459 $Y2=0.203
r97 44 45 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.167
r98 43 47 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r99 42 66 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r100 42 44 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.165
r101 40 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.106 $X2=0.459 $Y2=0.114
r102 39 40 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.099 $X2=0.459 $Y2=0.106
r103 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.099
r104 37 66 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r105 37 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.114
r106 36 62 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r107 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.081
r108 34 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.234 $X2=0.434 $Y2=0.234
r109 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.418 $Y2=0.234
r110 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r111 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r112 25 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r113 25 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.434 $Y2=0.234
r114 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r115 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r116 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r117 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r118 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r119 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r120 13 60 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r121 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r122 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r123 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r124 5 50 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.131 $X2=0.567
+ $Y2=0.131
r125 5 7 370.904 $w=2e-08 $l=9.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1305 $X2=0.567 $Y2=0.2295
r126 2 5 337.185 $w=2e-08 $l=9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.1305
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%9 2 5 7 9 14 21 25 26 30 31 32 33 34 39 40 42 44
+ 45 VSS
c24 46 VSS 2.95823e-19 $X=0.945 $Y=0.171
c25 45 VSS 9.82796e-19 $X=0.945 $Y=0.167
c26 44 VSS 3.06877e-19 $X=0.945 $Y=0.122
c27 43 VSS 0.00344802f $X=0.945 $Y=0.117
c28 42 VSS 0.00284656f $X=0.945 $Y=0.225
c29 40 VSS 0.0018377f $X=0.918 $Y=0.234
c30 39 VSS 0.00568507f $X=0.9 $Y=0.234
c31 34 VSS 0.00462933f $X=0.936 $Y=0.234
c32 33 VSS 0.00189638f $X=0.9 $Y=0.036
c33 32 VSS 0.0035379f $X=0.882 $Y=0.036
c34 31 VSS 0.00146362f $X=0.846 $Y=0.036
c35 30 VSS 0.00480249f $X=0.828 $Y=0.036
c36 26 VSS 0.00226308f $X=0.792 $Y=0.036
c37 25 VSS 0.00657446f $X=0.936 $Y=0.036
c38 21 VSS 0.00135803f $X=0.783 $Y=0.105
c39 17 VSS 0.00535489f $X=0.862 $Y=0.2295
c40 12 VSS 0.00569943f $X=0.862 $Y=0.0405
c41 5 VSS 0.00257499f $X=0.783 $Y=0.1055
c42 2 VSS 0.0589361f $X=0.783 $Y=0.0405
r43 45 46 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.167 $X2=0.945 $Y2=0.171
r44 44 45 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.122 $X2=0.945 $Y2=0.167
r45 43 44 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.117 $X2=0.945 $Y2=0.122
r46 42 46 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.171
r47 41 43 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.117
r48 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.234 $X2=0.918 $Y2=0.234
r49 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.9 $Y2=0.234
r50 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r51 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.918 $Y2=0.234
r52 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r53 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.846 $Y2=0.036
r54 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r55 28 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.846 $Y2=0.036
r56 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.036 $X2=0.828 $Y2=0.036
r57 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r58 25 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.9 $Y2=0.036
r59 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.783 $Y=0.045 $X2=0.792 $Y2=0.036
r60 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.105
r61 17 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234 $X2=0.864
+ $Y2=0.234
r62 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2295 $X2=0.862 $Y2=0.2295
r63 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036 $X2=0.864
+ $Y2=0.036
r64 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.862 $Y2=0.0405
r65 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.105 $X2=0.783
+ $Y2=0.105
r66 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.1055 $X2=0.783 $Y2=0.2295
r67 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.1055
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%10 2 5 7 10 15 18 21 23 25 26 29 30 31 34 35 40
+ 41 43 45 46 47 48 49 51 52 54 55 58 65 66 74 77 81 84 92 VSS
c69 92 VSS 0.00121551f $X=0.999 $Y=0.136
c70 84 VSS 0.00773455f $X=0.999 $Y=0.153
c71 81 VSS 0.00168283f $X=0.891 $Y=0.153
c72 78 VSS 4.17512e-19 $X=0.837 $Y=0.162
c73 77 VSS 1.52743e-19 $X=0.729 $Y=0.162
c74 74 VSS 0.00357422f $X=0.72 $Y=0.233
c75 73 VSS 0.00244813f $X=0.729 $Y=0.233
c76 66 VSS 4.13886e-19 $X=0.866 $Y=0.162
c77 65 VSS 1.21361e-19 $X=0.85 $Y=0.162
c78 63 VSS 2.72392e-19 $X=0.882 $Y=0.162
c79 58 VSS 3.90416e-19 $X=0.837 $Y=0.135
c80 55 VSS 3.26354e-19 $X=0.792 $Y=0.162
c81 54 VSS 0.00200395f $X=0.774 $Y=0.162
c82 52 VSS 0.00182633f $X=0.828 $Y=0.162
c83 51 VSS 0.00126232f $X=0.729 $Y=0.224
c84 49 VSS 1.52219e-19 $X=0.729 $Y=0.136
c85 48 VSS 2.77769e-19 $X=0.729 $Y=0.119
c86 47 VSS 1.41609e-19 $X=0.729 $Y=0.101
c87 46 VSS 3.47341e-19 $X=0.729 $Y=0.081
c88 45 VSS 2.73935e-19 $X=0.729 $Y=0.153
c89 43 VSS 0.00166747f $X=0.704 $Y=0.036
c90 42 VSS 4.5912e-19 $X=0.688 $Y=0.036
c91 41 VSS 0.00146362f $X=0.684 $Y=0.036
c92 40 VSS 0.00375499f $X=0.666 $Y=0.036
c93 35 VSS 0.00402292f $X=0.72 $Y=0.036
c94 34 VSS 0.00153815f $X=0.702 $Y=0.2295
c95 30 VSS 6.50675e-19 $X=0.719 $Y=0.2295
c96 29 VSS 0.0322408f $X=0.648 $Y=0.0405
c97 25 VSS 5.63046e-19 $X=0.665 $Y=0.0405
c98 21 VSS 0.00425984f $X=1.053 $Y=0.136
c99 18 VSS 0.0584171f $X=1.053 $Y=0.0675
c100 10 VSS 0.0615046f $X=0.999 $Y=0.0675
c101 5 VSS 0.00238412f $X=0.837 $Y=0.135
c102 2 VSS 0.0618222f $X=0.837 $Y=0.0405
r103 84 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.999 $Y=0.153 $X2=0.999
+ $Y2=0.153
r104 80 84 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.999 $Y2=0.153
r105 80 81 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r106 74 75 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.233 $X2=0.7245 $Y2=0.233
r107 73 75 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.233 $X2=0.7245 $Y2=0.233
r108 70 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.233 $X2=0.72 $Y2=0.233
r109 65 66 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.85
+ $Y=0.162 $X2=0.866 $Y2=0.162
r110 64 78 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.837 $Y2=0.162
r111 64 65 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.85 $Y2=0.162
r112 63 81 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.891 $Y2=0.162
r113 63 66 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.866 $Y2=0.162
r114 56 78 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.162
r115 56 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.135
r116 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.162 $X2=0.792 $Y2=0.162
r117 53 77 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.729 $Y2=0.162
r118 53 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.774 $Y2=0.162
r119 52 78 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.837 $Y2=0.162
r120 52 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.792 $Y2=0.162
r121 51 73 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.224 $X2=0.729 $Y2=0.233
r122 50 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.162
r123 50 51 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.224
r124 48 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.119 $X2=0.729 $Y2=0.136
r125 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.101 $X2=0.729 $Y2=0.119
r126 46 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.081 $X2=0.729 $Y2=0.101
r127 45 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.162
r128 45 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.136
r129 44 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.045 $X2=0.729 $Y2=0.081
r130 42 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.036 $X2=0.704 $Y2=0.036
r131 41 42 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.688 $Y2=0.036
r132 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.684 $Y2=0.036
r133 37 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.666 $Y2=0.036
r134 35 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.036 $X2=0.729 $Y2=0.045
r135 35 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.704 $Y2=0.036
r136 34 70 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.233
+ $X2=0.702 $Y2=0.233
r137 31 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2295 $X2=0.702 $Y2=0.2295
r138 30 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2295 $X2=0.702 $Y2=0.2295
r139 29 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r140 26 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0405 $X2=0.648 $Y2=0.0405
r141 25 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r142 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.136 $X2=1.053 $Y2=0.2025
r143 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.0675 $X2=1.053 $Y2=0.136
r144 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.999
+ $Y=0.136 $X2=1.053 $Y2=0.136
r145 13 92 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.136 $X2=0.999
+ $Y2=0.136
r146 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.136 $X2=0.999 $Y2=0.2025
r147 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.136
r148 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.135 $X2=0.837
+ $Y2=0.135
r149 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.2295
r150 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.0405 $X2=0.837 $Y2=0.135
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%11 2 7 10 15 18 23 26 29 31 33 34 38 39 42 43 46
+ 48 54 55 58 59 63 66 68 VSS
c43 68 VSS 3.78938e-19 $X=1.089 $Y=0.136
c44 66 VSS 4.82002e-21 $X=1.143 $Y=0.136
c45 65 VSS 7.16275e-19 $X=1.125 $Y=0.136
c46 63 VSS 1.52274e-19 $X=1.161 $Y=0.136
c47 60 VSS 0.00141149f $X=1.089 $Y=0.201
c48 59 VSS 8.53779e-19 $X=1.089 $Y=0.167
c49 58 VSS 6.05349e-19 $X=1.089 $Y=0.225
c50 56 VSS 0.00227099f $X=1.089 $Y=0.122
c51 55 VSS 7.78235e-19 $X=1.089 $Y=0.069
c52 54 VSS 3.06947e-19 $X=1.089 $Y=0.127
c53 48 VSS 0.0110409f $X=1.08 $Y=0.234
c54 46 VSS 0.00899572f $X=1.026 $Y=0.036
c55 43 VSS 0.0110409f $X=1.08 $Y=0.036
c56 42 VSS 0.00937164f $X=1.026 $Y=0.2025
c57 38 VSS 5.72268e-19 $X=1.043 $Y=0.2025
c58 33 VSS 5.72268e-19 $X=1.043 $Y=0.0675
c59 29 VSS 0.0143997f $X=1.269 $Y=0.136
c60 26 VSS 0.0615048f $X=1.269 $Y=0.0675
c61 18 VSS 0.0615873f $X=1.215 $Y=0.0675
c62 10 VSS 0.061355f $X=1.161 $Y=0.0675
c63 2 VSS 0.0588241f $X=1.107 $Y=0.0675
r64 65 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.125
+ $Y=0.136 $X2=1.143 $Y2=0.136
r65 63 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.136 $X2=1.143 $Y2=0.136
r66 61 68 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.136 $X2=1.089 $Y2=0.136
r67 61 65 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.136 $X2=1.125 $Y2=0.136
r68 59 60 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.167 $X2=1.089 $Y2=0.201
r69 58 60 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.225 $X2=1.089 $Y2=0.201
r70 57 68 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.145 $X2=1.089 $Y2=0.136
r71 57 59 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.145 $X2=1.089 $Y2=0.167
r72 55 56 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.069 $X2=1.089 $Y2=0.122
r73 54 68 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.127 $X2=1.089 $Y2=0.136
r74 54 56 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.127 $X2=1.089 $Y2=0.122
r75 53 55 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.045 $X2=1.089 $Y2=0.069
r76 48 58 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.08 $Y=0.234 $X2=1.089 $Y2=0.225
r77 48 50 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.026 $Y2=0.234
r78 45 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.036 $X2=1.026
+ $Y2=0.036
r79 43 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.08 $Y=0.036 $X2=1.089 $Y2=0.045
r80 43 45 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.036 $X2=1.026 $Y2=0.036
r81 42 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.234 $X2=1.026
+ $Y2=0.234
r82 39 42 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.2025 $X2=1.026 $Y2=0.2025
r83 38 42 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.043 $Y=0.2025 $X2=1.026 $Y2=0.2025
r84 37 46 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.026
+ $Y=0.0675 $X2=1.026 $Y2=0.036
r85 34 37 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.0675 $X2=1.026 $Y2=0.0675
r86 33 37 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.043 $Y=0.0675 $X2=1.026 $Y2=0.0675
r87 29 31 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.269
+ $Y=0.136 $X2=1.269 $Y2=0.2025
r88 26 29 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.269
+ $Y=0.0675 $X2=1.269 $Y2=0.136
r89 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.215
+ $Y=0.136 $X2=1.269 $Y2=0.136
r90 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.215
+ $Y=0.136 $X2=1.215 $Y2=0.2025
r91 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.215
+ $Y=0.0675 $X2=1.215 $Y2=0.136
r92 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.161
+ $Y=0.136 $X2=1.215 $Y2=0.136
r93 13 63 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.161 $Y=0.136 $X2=1.161
+ $Y2=0.136
r94 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.161
+ $Y=0.136 $X2=1.161 $Y2=0.2025
r95 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.161
+ $Y=0.0675 $X2=1.161 $Y2=0.136
r96 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.107
+ $Y=0.136 $X2=1.161 $Y2=0.136
r97 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.107
+ $Y=0.136 $X2=1.107 $Y2=0.2025
r98 2 5 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.107
+ $Y=0.0675 $X2=1.107 $Y2=0.136
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%Q 1 2 5 6 7 11 12 15 16 17 20 21 25 26 28 33 38
+ 40 43 46 49 52 VSS
c27 55 VSS 0.00197453f $X=1.134 $Y=0.234
c28 52 VSS 8.50672e-19 $X=1.134 $Y=0.216
c29 49 VSS 1.39487e-19 $X=1.134 $Y=0.0495
c30 46 VSS 6.94854e-19 $X=1.134 $Y=0.054
c31 43 VSS 0.00199537f $X=1.134 $Y=0.036
c32 42 VSS 0.00435712f $X=1.323 $Y=0.201
c33 40 VSS 0.0045092f $X=1.323 $Y=0.127
c34 39 VSS 0.0010981f $X=1.323 $Y=0.069
c35 38 VSS 9.20903e-19 $X=1.329 $Y=0.134
c36 36 VSS 0.0010981f $X=1.323 $Y=0.225
c37 34 VSS 0.00545672f $X=1.2085 $Y=0.234
c38 33 VSS 0.00256929f $X=1.175 $Y=0.234
c39 28 VSS 0.0155121f $X=1.313 $Y=0.234
c40 27 VSS 0.0054658f $X=1.2085 $Y=0.036
c41 26 VSS 0.0025515f $X=1.175 $Y=0.036
c42 25 VSS 0.00926069f $X=1.242 $Y=0.036
c43 21 VSS 0.0155121f $X=1.313 $Y=0.036
c44 20 VSS 0.00929505f $X=1.242 $Y=0.2025
c45 16 VSS 5.38922e-19 $X=1.259 $Y=0.2025
c46 15 VSS 0.0105438f $X=1.134 $Y=0.2025
c47 11 VSS 5.945e-19 $X=1.151 $Y=0.2025
c48 6 VSS 5.38922e-19 $X=1.259 $Y=0.0675
c49 5 VSS 0.010566f $X=1.134 $Y=0.0675
c50 1 VSS 5.945e-19 $X=1.151 $Y=0.0675
r51 56 57 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.225 $X2=1.134 $Y2=0.2295
r52 55 57 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.234 $X2=1.134 $Y2=0.2295
r53 52 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.216 $X2=1.134 $Y2=0.225
r54 48 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.045 $X2=1.134 $Y2=0.0495
r55 46 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.054 $X2=1.134 $Y2=0.0495
r56 43 48 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.036 $X2=1.134 $Y2=0.045
r57 41 42 3.3358 $w=2e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.145 $X2=1.323 $Y2=0.201
r58 39 40 3.45494 $w=2e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.069 $X2=1.323 $Y2=0.127
r59 38 41 0.655247 $w=2e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.134 $X2=1.323 $Y2=0.145
r60 38 40 0.416975 $w=2e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.134 $X2=1.323 $Y2=0.127
r61 36 42 1.42963 $w=2e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.225 $X2=1.323 $Y2=0.201
r62 35 39 1.42963 $w=2e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.045 $X2=1.323 $Y2=0.069
r63 33 34 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.175
+ $Y=0.234 $X2=1.2085 $Y2=0.234
r64 31 34 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.242
+ $Y=0.234 $X2=1.2085 $Y2=0.234
r65 29 55 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.143
+ $Y=0.234 $X2=1.134 $Y2=0.234
r66 29 33 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.143
+ $Y=0.234 $X2=1.175 $Y2=0.234
r67 28 36 0.685354 $w=2e-08 $l=1.3784e-08 $layer=M1 $thickness=3.6e-08 $X=1.313
+ $Y=0.234 $X2=1.323 $Y2=0.225
r68 28 31 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.313
+ $Y=0.234 $X2=1.242 $Y2=0.234
r69 26 27 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.175
+ $Y=0.036 $X2=1.2085 $Y2=0.036
r70 24 27 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.242
+ $Y=0.036 $X2=1.2085 $Y2=0.036
r71 24 25 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.242 $Y=0.036 $X2=1.242
+ $Y2=0.036
r72 22 43 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.143
+ $Y=0.036 $X2=1.134 $Y2=0.036
r73 22 26 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.143
+ $Y=0.036 $X2=1.175 $Y2=0.036
r74 21 35 0.685354 $w=2e-08 $l=1.3784e-08 $layer=M1 $thickness=3.6e-08 $X=1.313
+ $Y=0.036 $X2=1.323 $Y2=0.045
r75 21 24 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.313
+ $Y=0.036 $X2=1.242 $Y2=0.036
r76 20 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.242 $Y=0.234 $X2=1.242
+ $Y2=0.234
r77 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.225 $Y=0.2025 $X2=1.242 $Y2=0.2025
r78 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.259 $Y=0.2025 $X2=1.242 $Y2=0.2025
r79 15 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.134 $Y=0.216 $X2=1.134
+ $Y2=0.216
r80 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.117 $Y=0.2025 $X2=1.134 $Y2=0.2025
r81 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.151 $Y=0.2025 $X2=1.134 $Y2=0.2025
r82 10 25 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.242
+ $Y=0.0675 $X2=1.242 $Y2=0.036
r83 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.225 $Y=0.0675 $X2=1.242 $Y2=0.0675
r84 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.259 $Y=0.0675 $X2=1.242 $Y2=0.0675
r85 5 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.134 $Y=0.054 $X2=1.134
+ $Y2=0.054
r86 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.117
+ $Y=0.0675 $X2=1.134 $Y2=0.0675
r87 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.151
+ $Y=0.0675 $X2=1.134 $Y2=0.0675
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%13 1 6 9 VSS
c6 9 VSS 0.0268266f $X=0.38 $Y=0.0675
c7 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c8 4 VSS 3.25039e-19 $X=0.322 $Y=0.0675
r9 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r10 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%14 1 6 9 VSS
c10 9 VSS 0.0221513f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.6182e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%15 1 6 9 VSS
c8 9 VSS 0.0223778f $X=0.758 $Y=0.0405
c9 6 VSS 3.14771e-19 $X=0.773 $Y=0.0405
c10 4 VSS 2.6194e-19 $X=0.7 $Y=0.0405
r11 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r12 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.7
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r13 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.685
+ $Y=0.0405 $X2=0.7 $Y2=0.0405
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%16 1 2 VSS
c0 1 VSS 0.00225696f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%17 1 2 VSS
c3 1 VSS 0.00231486f $X=0.341 $Y=0.2025
r4 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends

.subckt PM_DFFHQX4_ASAP7_75T_SRAM%18 1 2 VSS
c0 1 VSS 0.00219822f $X=0.773 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2295 $X2=0.739 $Y2=0.2295
.ends


* END of "./DFFHQx4_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DFFHQx4_ASAP7_75t_SRAM  VSS VDD CLK D Q
* 
* Q	Q
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_13_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_4_M3_g N_13_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_16_M4_d N_6_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_16_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_10_M7_d N_6_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.611
+ $Y=0.027
M8 N_15_M8_d N_4_M8_g N_10_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M9 VSS N_9_M9_g N_15_M9_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_9_M10_d N_10_M10_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.027
M11 N_11_M11_d N_10_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M12 N_11_M12_d N_10_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.027
M13 N_Q_M13_d N_11_M13_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.027
M14 N_Q_M14_d N_11_M14_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.151
+ $Y=0.027
M15 N_Q_M15_d N_11_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.027
M16 N_Q_M16_d N_11_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M17 VDD N_CLK_M17_g N_4_M17_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M18 N_6_M18_d N_4_M18_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M19 N_17_M19_d N_D_M19_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M20 N_8_M20_d N_6_M20_g N_17_M20_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M21 N_14_M21_d N_4_M21_g N_8_M21_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M22 VDD N_7_M22_g N_14_M22_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M23 N_7_M23_d N_8_M23_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M24 N_10_M24_d N_4_M24_g N_7_M24_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.665 $Y=0.216
M25 N_18_M25_d N_6_M25_g N_10_M25_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.719 $Y=0.216
M26 VDD N_9_M26_g N_18_M26_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M27 N_9_M27_d N_10_M27_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.216
M28 N_11_M28_d N_10_M28_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
M29 N_11_M29_d N_10_M29_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.162
M30 N_Q_M30_d N_11_M30_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.162
M31 N_Q_M31_d N_11_M31_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.151
+ $Y=0.162
M32 N_Q_M32_d N_11_M32_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.162
M33 N_Q_M33_d N_11_M33_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
*
* 
* .include "DFFHQx4_ASAP7_75t_SRAM.pex.sp.DFFHQX4_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DFFHQx4_ASAP7_75t_SRAM.pex.sp.DFFHQX4_ASAP7_75T_SRAM.pxi"
* File: DFFHQx4_ASAP7_75t_SRAM.pex.sp.DFFHQX4_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:25:16 2017
* 
x_PM_DFFHQX4_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_13_p N_CLK_M17_g CLK N_CLK_c_6_p
+ VSS PM_DFFHQX4_ASAP7_75T_SRAM%CLK
x_PM_DFFHQX4_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M18_g N_4_M3_g N_4_c_43_p N_4_M21_g
+ N_4_M8_g N_4_c_48_p N_4_M24_g N_4_M0_s N_4_c_22_n N_4_M17_s N_4_c_23_n
+ N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_28_n N_4_c_29_n N_4_c_30_n
+ N_4_c_31_n N_4_c_40_p N_4_c_49_p N_4_c_37_p N_4_c_69_p N_4_c_33_n N_4_c_34_n
+ N_4_c_39_p N_4_c_51_p VSS PM_DFFHQX4_ASAP7_75T_SRAM%4
x_PM_DFFHQX4_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_102_n N_D_M19_g N_D_c_116_p D
+ N_D_c_104_n N_D_c_112_p N_D_c_105_n N_D_c_106_n VSS PM_DFFHQX4_ASAP7_75T_SRAM%D
x_PM_DFFHQX4_ASAP7_75T_SRAM%6 N_6_c_124_n N_6_M20_g N_6_M4_g N_6_M7_g N_6_c_173_p
+ N_6_c_128_n N_6_M25_g N_6_c_185_p N_6_c_129_n N_6_M1_d N_6_M18_d N_6_c_119_n
+ N_6_c_152_n N_6_c_135_n N_6_c_120_n N_6_c_153_n N_6_c_121_n N_6_c_138_n
+ N_6_c_139_n N_6_c_140_n N_6_c_141_n N_6_c_142_n N_6_c_122_n N_6_c_145_n
+ N_6_c_123_n N_6_c_146_n N_6_c_148_n N_6_c_190_p VSS PM_DFFHQX4_ASAP7_75T_SRAM%6
x_PM_DFFHQX4_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_245_p N_7_M22_g N_7_M7_s N_7_M6_d
+ N_7_c_231_n N_7_M23_d N_7_c_232_n N_7_M24_s N_7_c_234_n N_7_c_243_p
+ N_7_c_221_n N_7_c_261_p N_7_c_222_n N_7_c_244_p N_7_c_262_p N_7_c_224_n
+ N_7_c_247_p N_7_c_225_n N_7_c_238_n N_7_c_239_n N_7_c_241_n N_7_c_226_n VSS
+ PM_DFFHQX4_ASAP7_75T_SRAM%7
x_PM_DFFHQX4_ASAP7_75T_SRAM%8 N_8_M6_g N_8_c_264_n N_8_M23_g N_8_M3_d N_8_M4_s
+ N_8_M20_d N_8_c_267_n N_8_M21_s N_8_c_313_p N_8_c_279_n N_8_c_268_n
+ N_8_c_314_p N_8_c_270_n N_8_c_286_n N_8_c_287_n N_8_c_271_n N_8_c_315_p
+ N_8_c_272_n N_8_c_289_n N_8_c_291_n N_8_c_304_n N_8_c_274_n N_8_c_305_n
+ N_8_c_296_n N_8_c_275_n N_8_c_276_n N_8_c_277_n N_8_c_278_n VSS
+ PM_DFFHQX4_ASAP7_75T_SRAM%8
x_PM_DFFHQX4_ASAP7_75T_SRAM%9 N_9_M9_g N_9_c_323_p N_9_M26_g N_9_M10_d N_9_M27_d
+ N_9_c_322_p N_9_c_334_p N_9_c_321_p N_9_c_326_p N_9_c_320_p N_9_c_330_p
+ N_9_c_332_p N_9_c_339_p N_9_c_331_p N_9_c_335_p N_9_c_325_p N_9_c_333_p
+ N_9_c_336_p VSS PM_DFFHQX4_ASAP7_75T_SRAM%9
x_PM_DFFHQX4_ASAP7_75T_SRAM%10 N_10_M10_g N_10_c_341_n N_10_M27_g N_10_M11_g
+ N_10_M28_g N_10_M12_g N_10_c_394_p N_10_M29_g N_10_M8_s N_10_M7_d N_10_c_342_n
+ N_10_M25_s N_10_M24_d N_10_c_352_n N_10_c_374_n N_10_c_343_n N_10_c_344_n
+ N_10_c_407_p N_10_c_346_n N_10_c_366_n N_10_c_353_n N_10_c_347_n N_10_c_354_n
+ N_10_c_355_n N_10_c_379_n N_10_c_357_n N_10_c_380_n N_10_c_382_n N_10_c_383_n
+ N_10_c_384_n N_10_c_358_n N_10_c_359_n N_10_c_385_n N_10_c_348_n N_10_c_390_n
+ VSS PM_DFFHQX4_ASAP7_75T_SRAM%10
x_PM_DFFHQX4_ASAP7_75T_SRAM%11 N_11_M13_g N_11_M30_g N_11_M14_g N_11_M31_g
+ N_11_M15_g N_11_M32_g N_11_M16_g N_11_c_415_n N_11_M33_g N_11_M12_d N_11_M11_d
+ N_11_M29_d N_11_M28_d N_11_c_418_n N_11_c_410_n N_11_c_421_n N_11_c_411_n
+ N_11_c_424_n N_11_c_450_p N_11_c_451_p N_11_c_432_p N_11_c_440_p N_11_c_449_p
+ N_11_c_425_n VSS PM_DFFHQX4_ASAP7_75T_SRAM%11
x_PM_DFFHQX4_ASAP7_75T_SRAM%Q N_Q_M14_d N_Q_M13_d N_Q_c_454_n N_Q_M16_d N_Q_M15_d
+ N_Q_M31_d N_Q_M30_d N_Q_c_458_n N_Q_M33_d N_Q_M32_d N_Q_c_461_n N_Q_c_462_n
+ N_Q_c_464_n N_Q_c_465_n N_Q_c_468_n N_Q_c_470_n Q N_Q_c_474_n N_Q_c_475_n
+ N_Q_c_476_n N_Q_c_477_n N_Q_c_478_n VSS PM_DFFHQX4_ASAP7_75T_SRAM%Q
x_PM_DFFHQX4_ASAP7_75T_SRAM%13 N_13_M2_d N_13_M3_s N_13_c_480_n VSS
+ PM_DFFHQX4_ASAP7_75T_SRAM%13
x_PM_DFFHQX4_ASAP7_75T_SRAM%14 N_14_M21_d N_14_M22_s N_14_c_487_n VSS
+ PM_DFFHQX4_ASAP7_75T_SRAM%14
x_PM_DFFHQX4_ASAP7_75T_SRAM%15 N_15_M8_d N_15_M9_s N_15_c_496_n VSS
+ PM_DFFHQX4_ASAP7_75T_SRAM%15
x_PM_DFFHQX4_ASAP7_75T_SRAM%16 N_16_M5_s N_16_M4_d VSS PM_DFFHQX4_ASAP7_75T_SRAM%16
x_PM_DFFHQX4_ASAP7_75T_SRAM%17 N_17_M20_s N_17_M19_d VSS PM_DFFHQX4_ASAP7_75T_SRAM%17
x_PM_DFFHQX4_ASAP7_75T_SRAM%18 N_18_M26_s N_18_M25_d VSS PM_DFFHQX4_ASAP7_75T_SRAM%18
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_22_n 3.57152e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 CLK N_4_c_23_n 0.00136255f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.144
cc_4 CLK N_4_c_24_n 2.75361e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.07
cc_5 CLK N_4_c_25_n 0.00136255f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.107
cc_6 N_CLK_c_6_p N_4_c_26_n 0.00145637f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2
cc_7 N_CLK_c_6_p N_4_c_27_n 2.75361e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2125
cc_8 CLK N_4_c_28_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_6_p N_4_c_29_n 5.03453e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_6_p N_4_c_30_n 0.00123168f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.153
cc_11 CLK N_4_c_31_n 4.93618e-19 $X=0.082 $Y=0.119 $X2=0.175 $Y2=0.153
cc_12 N_CLK_c_6_p N_4_c_31_n 0.00162391f $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_13 N_CLK_c_13_p N_4_c_33_n 0.00109779f $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.135
cc_14 CLK N_4_c_34_n 0.00174841f $X=0.082 $Y=0.119 $X2=0.151 $Y2=0.135
cc_15 N_CLK_c_6_p N_4_c_34_n 3.29534e-19 $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.135
cc_16 CLK N_6_c_119_n 6.37157e-19 $X=0.082 $Y=0.119 $X2=0.027 $Y2=0.234
cc_17 N_CLK_c_6_p N_6_c_120_n 6.45547e-19 $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.153
cc_18 N_CLK_c_6_p N_6_c_121_n 0.00124695f $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_19 N_CLK_c_6_p N_6_c_122_n 3.64822e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_20 CLK N_6_c_123_n 0.00136827f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.153
cc_21 N_4_M3_g N_D_M2_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_22 N_4_c_37_p N_D_c_102_n 2.91747e-19 $X=0.527 $Y=0.153 $X2=0.081 $Y2=0.135
cc_23 N_4_c_33_n N_D_c_102_n 2.04625e-19 $X=0.151 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_4_c_39_p N_D_c_104_n 2.3983e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_25 N_4_c_40_p N_D_c_105_n 8.99815e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_26 N_4_c_40_p N_D_c_106_n 8.75229e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_27 N_4_M3_g N_6_c_124_n 0.00355599f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_28 N_4_c_43_p N_6_c_124_n 0.00125076f $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.054
cc_29 N_4_M3_g N_6_M4_g 0.00355599f $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_4_M8_g N_6_M7_g 0.00355599f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_31 N_4_M8_g N_6_c_128_n 0.00355599f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_32 N_4_M8_g N_6_c_129_n 0.00250099f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_33 N_4_c_48_p N_6_c_129_n 0.00180656f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_34 N_4_c_49_p N_6_c_129_n 6.63386e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_35 N_4_c_37_p N_6_c_129_n 0.00187561f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_36 N_4_c_51_p N_6_c_129_n 0.00123876f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_34_n N_6_c_119_n 2.97444e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_31_n N_6_c_135_n 2.38327e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_34_n N_6_c_120_n 2.85146e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_40_p N_6_c_121_n 2.46239e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_41 N_4_c_31_n N_6_c_138_n 2.31165e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_42 N_4_c_39_p N_6_c_139_n 9.24693e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_43 N_4_c_37_p N_6_c_140_n 3.67557e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_44 N_4_c_37_p N_6_c_141_n 8.06691e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_45 N_4_c_37_p N_6_c_142_n 2.46239e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_46 N_4_c_40_p N_6_c_122_n 0.0299327f $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_39_p N_6_c_122_n 2.98936e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_48 N_4_c_37_p N_6_c_145_n 2.81476e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_49 N_4_c_40_p N_6_c_146_n 8.79704e-19 $X=0.29 $Y=0.153 $X2=0 $Y2=0
cc_50 N_4_c_34_n N_6_c_146_n 0.00524677f $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_51 N_4_c_37_p N_6_c_148_n 9.92294e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_52 N_4_c_39_p N_6_c_148_n 5.5596e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_53 N_4_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_54 N_4_c_69_p N_7_c_221_n 2.95658e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_55 N_4_c_49_p N_7_c_222_n 2.61213e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_56 N_4_c_69_p N_7_c_222_n 2.61213e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_57 N_4_c_51_p N_7_c_224_n 0.0031817f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_58 N_4_c_49_p N_7_c_225_n 0.00115177f $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_59 N_4_c_49_p N_7_c_226_n 2.95658e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_60 N_4_M8_g N_8_M6_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_61 N_4_c_43_p N_8_c_264_n 2.07716e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_62 N_4_c_48_p N_8_c_264_n 4.17807e-19 $X=0.675 $Y=0.135 $X2=0.081 $Y2=0.135
cc_63 N_4_c_69_p N_8_c_264_n 2.88013e-19 $X=0.601 $Y=0.153 $X2=0.081 $Y2=0.135
cc_64 N_4_c_39_p N_8_c_267_n 2.36208e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_65 N_4_M3_g N_8_c_268_n 3.49806e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_66 N_4_c_39_p N_8_c_268_n 3.83282e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_67 N_4_c_39_p N_8_c_270_n 7.28732e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_68 N_4_c_39_p N_8_c_271_n 7.28732e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_69 N_4_c_37_p N_8_c_272_n 0.00118282f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_70 N_4_c_39_p N_8_c_272_n 8.2214e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_71 N_4_c_37_p N_8_c_274_n 0.00138591f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_72 N_4_c_69_p N_8_c_275_n 0.00138591f $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_73 N_4_c_37_p N_8_c_276_n 2.54113e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_74 N_4_c_37_p N_8_c_277_n 3.92135e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_75 N_4_c_39_p N_8_c_278_n 7.28732e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_76 N_4_M8_g N_9_M9_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_77 N_4_c_48_p N_10_c_341_n 2.7571e-19 $X=0.675 $Y=0.135 $X2=0.081 $Y2=0.135
cc_78 N_4_c_49_p N_10_c_342_n 2.24654e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_79 N_4_c_49_p N_10_c_343_n 5.06919e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_80 N_4_M8_g N_10_c_344_n 3.47752e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_81 N_4_c_51_p N_10_c_344_n 5.72565e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_82 N_4_c_49_p N_10_c_346_n 2.46558e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_83 N_4_c_51_p N_10_c_347_n 0.00319931f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_84 N_4_c_49_p N_10_c_348_n 2.9112e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_85 N_4_c_37_p N_13_c_480_n 3.46326e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_86 N_D_M2_g N_6_c_124_n 0.00341068f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_87 N_D_c_102_n N_6_c_124_n 0.00113998f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.054
cc_88 D N_6_c_152_n 0.00215667f $X=0.244 $Y=0.082 $X2=0 $Y2=0
cc_89 N_D_c_106_n N_6_c_153_n 0.00215667f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_90 N_D_c_106_n N_6_c_121_n 0.00225008f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_91 N_D_c_112_p N_6_c_140_n 0.00127755f $X=0.281 $Y=0.135 $X2=0 $Y2=0
cc_92 N_D_c_102_n N_6_c_122_n 2.11668e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_93 N_D_c_106_n N_6_c_122_n 0.00122387f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_94 D N_6_c_123_n 0.00215667f $X=0.244 $Y=0.082 $X2=0 $Y2=0
cc_95 N_D_c_116_p N_6_c_146_n 0.00215667f $X=0.243 $Y=0.126 $X2=0 $Y2=0
cc_96 N_D_c_106_n N_6_c_148_n 0.00120973f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_97 N_D_c_106_n N_8_c_279_n 2.80198e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_98 N_6_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_99 N_6_M7_g N_7_M5_g 2.13359e-19 $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_100 N_6_c_129_n N_7_M5_g 0.00205839f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_101 N_6_c_145_n N_7_M5_g 3.15189e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_102 N_6_c_129_n N_7_c_231_n 5.5606e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_103 N_6_c_129_n N_7_c_232_n 2.12581e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_104 N_6_c_129_n N_7_M24_s 2.50995e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_105 N_6_M7_g N_7_c_234_n 0.00200088f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_106 N_6_c_129_n N_7_c_234_n 0.00303373f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_107 N_6_M7_g N_7_c_224_n 3.34915e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_108 N_6_M7_g N_7_c_225_n 2.25102e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_109 N_6_c_145_n N_7_c_238_n 5.75704e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_110 N_6_c_173_p N_7_c_239_n 0.00195059f $X=0.621 $Y=0.178 $X2=0 $Y2=0
cc_111 N_6_c_129_n N_7_c_239_n 0.00191847f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_112 N_6_M7_g N_7_c_241_n 3.80981e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_113 N_6_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_114 N_6_M7_g N_8_M6_g 0.00341068f $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_115 N_6_c_129_n N_8_M6_g 0.00303187f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_116 N_6_c_122_n N_8_c_267_n 3.12535e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_117 N_6_c_148_n N_8_c_267_n 8.9852e-19 $X=0.324 $Y=0.167 $X2=0 $Y2=0
cc_118 N_6_c_122_n N_8_c_279_n 0.0015935f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_119 N_6_M4_g N_8_c_286_n 3.68551e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_120 N_6_M4_g N_8_c_287_n 2.06635e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_121 N_6_M4_g N_8_c_272_n 2.25747e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_122 N_6_c_185_p N_8_c_289_n 2.70413e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_123 N_6_c_145_n N_8_c_289_n 0.00174159f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_124 N_6_c_185_p N_8_c_291_n 0.00171407f $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_125 N_6_c_129_n N_8_c_291_n 5.88593e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_126 N_6_c_122_n N_8_c_291_n 0.00104904f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_127 N_6_c_190_p N_8_c_291_n 2.15173e-19 $X=0.324 $Y=0.178 $X2=0 $Y2=0
cc_128 N_6_c_129_n N_8_c_274_n 8.16411e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_129 N_6_c_129_n N_8_c_296_n 3.32592e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_130 N_6_c_145_n N_8_c_296_n 8.9822e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_131 N_6_c_129_n N_8_c_275_n 4.52853e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_132 N_6_c_128_n N_9_M9_g 0.00341068f $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_133 N_6_c_128_n N_10_M10_g 2.13359e-19 $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_134 N_6_c_129_n N_10_c_342_n 8.28378e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_135 N_6_c_129_n N_10_M25_s 3.37661e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_136 N_6_c_129_n N_10_c_352_n 0.00134523f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_137 N_6_c_128_n N_10_c_353_n 3.01068e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_138 N_6_c_128_n N_10_c_354_n 2.58474e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_139 N_6_c_128_n N_10_c_355_n 0.00228871f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_140 N_6_c_129_n N_10_c_355_n 7.89371e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_141 N_6_c_128_n N_10_c_357_n 3.99306e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_142 N_6_c_129_n N_10_c_358_n 4.54272e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_143 N_6_c_128_n N_10_c_359_n 4.71808e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_144 N_6_c_129_n N_10_c_359_n 2.2968e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_145 N_6_c_124_n N_13_c_480_n 0.00515096f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_146 N_6_c_140_n N_13_c_480_n 0.00114179f $X=0.333 $Y=0.135 $X2=0 $Y2=0
cc_147 N_6_c_129_n N_14_M22_s 2.36286e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.216
cc_148 N_6_M4_g N_14_c_487_n 0.00200088f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_149 N_6_c_185_p N_14_c_487_n 5.41258e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_150 N_6_c_129_n N_14_c_487_n 0.00230928f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_151 N_6_c_122_n N_14_c_487_n 7.09553e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_152 N_6_c_128_n N_15_c_496_n 0.0019841f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_153 N_6_c_129_n N_15_c_496_n 4.3039e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_154 N_6_c_142_n N_17_M20_s 8.51186e-19 $X=0.324 $Y=0.189 $X2=0.081 $Y2=0.054
cc_155 N_6_c_148_n N_17_M20_s 2.57402e-19 $X=0.324 $Y=0.167 $X2=0.081 $Y2=0.054
cc_156 N_6_c_190_p N_17_M20_s 2.18007e-19 $X=0.324 $Y=0.178 $X2=0.081 $Y2=0.054
cc_157 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_158 N_7_c_243_p N_8_M6_g 3.91159e-19 $X=0.581 $Y=0.09 $X2=0.135 $Y2=0.054
cc_159 N_7_c_244_p N_8_c_286_n 3.48522e-19 $X=0.594 $Y=0.054 $X2=0.018 $Y2=0.107
cc_160 N_7_c_245_p N_8_c_287_n 3.19692e-19 $X=0.513 $Y=0.09 $X2=0.018 $Y2=0.162
cc_161 N_7_c_243_p N_8_c_287_n 0.00114151f $X=0.581 $Y=0.09 $X2=0.018 $Y2=0.162
cc_162 N_7_c_247_p N_8_c_304_n 9.68907e-19 $X=0.621 $Y=0.14 $X2=0.027 $Y2=0.234
cc_163 N_7_c_243_p N_8_c_305_n 0.00506529f $X=0.581 $Y=0.09 $X2=0.054 $Y2=0.234
cc_164 N_7_M5_g N_8_c_296_n 3.12986e-19 $X=0.513 $Y=0.0405 $X2=0.047 $Y2=0.234
cc_165 N_7_c_245_p N_8_c_276_n 5.2508e-19 $X=0.513 $Y=0.09 $X2=0 $Y2=0
cc_166 N_7_c_231_n N_8_c_276_n 3.32985e-19 $X=0.594 $Y=0.0405 $X2=0 $Y2=0
cc_167 N_7_c_231_n N_10_c_342_n 0.00265056f $X=0.594 $Y=0.0405 $X2=0 $Y2=0
cc_168 N_7_c_244_p N_10_c_342_n 3.2755e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_169 N_7_c_241_n N_10_c_342_n 2.52634e-19 $X=0.621 $Y=0.09 $X2=0 $Y2=0
cc_170 N_7_c_234_n N_10_c_352_n 0.00205649f $X=0.65 $Y=0.2295 $X2=0 $Y2=0
cc_171 N_7_c_231_n N_10_c_343_n 5.23227e-19 $X=0.594 $Y=0.0405 $X2=0.018
+ $Y2=0.225
cc_172 N_7_c_244_p N_10_c_366_n 2.3746e-19 $X=0.594 $Y=0.054 $X2=0.054 $Y2=0.036
cc_173 N_7_c_241_n N_10_c_353_n 4.4424e-19 $X=0.621 $Y=0.09 $X2=0.047 $Y2=0.036
cc_174 N_7_c_239_n N_10_c_355_n 4.4424e-19 $X=0.621 $Y=0.203 $X2=0.054 $Y2=0.234
cc_175 N_7_c_234_n N_10_c_358_n 3.64729e-19 $X=0.65 $Y=0.2295 $X2=0 $Y2=0
cc_176 N_7_c_261_p N_10_c_358_n 4.68959e-19 $X=0.612 $Y=0.234 $X2=0 $Y2=0
cc_177 N_7_c_262_p N_10_c_359_n 4.4424e-19 $X=0.621 $Y=0.101 $X2=0.151 $Y2=0.135
cc_178 N_8_c_267_n N_13_c_480_n 0.00119486f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_179 N_8_c_276_n N_13_c_480_n 0.00362439f $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_180 N_8_c_277_n N_13_c_480_n 5.36233e-19 $X=0.45 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_181 N_8_c_267_n N_14_c_487_n 0.0018138f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_182 N_8_c_313_p N_14_c_487_n 0.00209454f $X=0.45 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_183 N_8_c_314_p N_14_c_487_n 0.0013184f $X=0.434 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_184 N_8_c_315_p N_14_c_487_n 0.00119497f $X=0.459 $Y=0.225 $X2=0.405
+ $Y2=0.0675
cc_185 N_8_c_276_n N_14_c_487_n 6.06615e-19 $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_186 N_9_M9_g N_10_M10_g 0.00268443f $X=0.783 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_187 N_9_c_320_p N_10_M10_g 3.74489e-19 $X=0.846 $Y=0.036 $X2=0.135 $Y2=0.054
cc_188 N_9_c_321_p N_10_c_374_n 0.00141609f $X=0.792 $Y=0.036 $X2=0.018
+ $Y2=0.045
cc_189 N_9_c_322_p N_10_c_366_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.054
+ $Y2=0.036
cc_190 N_9_c_323_p N_10_c_353_n 3.34766e-19 $X=0.783 $Y=0.1055 $X2=0.047
+ $Y2=0.036
cc_191 N_9_c_322_p N_10_c_353_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.047
+ $Y2=0.036
cc_192 N_9_c_325_p N_10_c_355_n 2.26874e-19 $X=0.945 $Y=0.225 $X2=0.054
+ $Y2=0.234
cc_193 N_9_c_326_p N_10_c_379_n 2.56938e-19 $X=0.828 $Y=0.036 $X2=0.054
+ $Y2=0.234
cc_194 N_9_M9_g N_10_c_380_n 6.3699e-19 $X=0.783 $Y=0.0405 $X2=0.0505 $Y2=0.234
cc_195 N_9_c_322_p N_10_c_380_n 9.0998e-19 $X=0.783 $Y=0.105 $X2=0.0505
+ $Y2=0.234
cc_196 N_9_c_320_p N_10_c_382_n 4.40983e-19 $X=0.846 $Y=0.036 $X2=0.033
+ $Y2=0.153
cc_197 N_9_c_330_p N_10_c_383_n 5.04796e-19 $X=0.882 $Y=0.036 $X2=0.405
+ $Y2=0.153
cc_198 N_9_c_331_p N_10_c_384_n 0.00148937f $X=0.9 $Y=0.234 $X2=0.405 $Y2=0.153
cc_199 N_9_c_332_p N_10_c_385_n 4.52584e-19 $X=0.9 $Y=0.036 $X2=0 $Y2=0
cc_200 N_9_c_333_p N_10_c_385_n 0.00280793f $X=0.945 $Y=0.122 $X2=0 $Y2=0
cc_201 N_9_c_334_p N_10_c_348_n 2.40515e-19 $X=0.936 $Y=0.036 $X2=0 $Y2=0
cc_202 N_9_c_335_p N_10_c_348_n 7.44774e-19 $X=0.918 $Y=0.234 $X2=0 $Y2=0
cc_203 N_9_c_336_p N_10_c_348_n 8.84468e-19 $X=0.945 $Y=0.167 $X2=0 $Y2=0
cc_204 N_9_c_336_p N_10_c_390_n 0.00213032f $X=0.945 $Y=0.167 $X2=0 $Y2=0
cc_205 N_9_c_334_p N_11_c_410_n 4.57392e-19 $X=0.936 $Y=0.036 $X2=0.027
+ $Y2=0.036
cc_206 N_9_c_339_p N_11_c_411_n 4.495e-19 $X=0.936 $Y=0.234 $X2=0.0505 $Y2=0.036
cc_207 N_9_c_321_p N_15_c_496_n 7.33799e-19 $X=0.792 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_208 N_10_M11_g N_11_M13_g 2.13359e-19 $X=0.999 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_209 N_10_M12_g N_11_M13_g 0.00268443f $X=1.053 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_210 N_10_M12_g N_11_M14_g 2.13359e-19 $X=1.053 $Y=0.0675 $X2=0.405 $Y2=0.0675
cc_211 N_10_c_394_p N_11_c_415_n 0.00102658f $X=1.053 $Y=0.136 $X2=0 $Y2=0
cc_212 N_10_c_394_p N_11_M12_d 3.7444e-19 $X=1.053 $Y=0.136 $X2=0.056 $Y2=0.216
cc_213 N_10_c_394_p N_11_M29_d 3.85232e-19 $X=1.053 $Y=0.136 $X2=0.018 $Y2=0.107
cc_214 N_10_c_394_p N_11_c_418_n 8.43851e-19 $X=1.053 $Y=0.136 $X2=0.018
+ $Y2=0.2125
cc_215 N_10_M12_g N_11_c_410_n 4.61823e-19 $X=1.053 $Y=0.0675 $X2=0.027
+ $Y2=0.036
cc_216 N_10_c_394_p N_11_c_410_n 5.30021e-19 $X=1.053 $Y=0.136 $X2=0.027
+ $Y2=0.036
cc_217 N_10_c_394_p N_11_c_421_n 7.60428e-19 $X=1.053 $Y=0.136 $X2=0.054
+ $Y2=0.036
cc_218 N_10_M12_g N_11_c_411_n 4.56718e-19 $X=1.053 $Y=0.0675 $X2=0.0505
+ $Y2=0.036
cc_219 N_10_c_394_p N_11_c_411_n 5.38938e-19 $X=1.053 $Y=0.136 $X2=0.0505
+ $Y2=0.036
cc_220 N_10_c_390_n N_11_c_424_n 0.00103215f $X=0.999 $Y=0.136 $X2=0.047
+ $Y2=0.234
cc_221 N_10_c_348_n N_11_c_425_n 3.06386e-19 $X=0.999 $Y=0.153 $X2=0.29
+ $Y2=0.153
cc_222 N_10_c_342_n N_15_c_496_n 0.0018138f $X=0.648 $Y=0.0405 $X2=0.405
+ $Y2=0.0675
cc_223 N_10_c_374_n N_15_c_496_n 0.0020512f $X=0.72 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_224 N_10_c_407_p N_15_c_496_n 0.00131745f $X=0.704 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_225 N_10_c_366_n N_15_c_496_n 0.00103564f $X=0.729 $Y=0.081 $X2=0.405
+ $Y2=0.0675
cc_226 N_10_c_357_n N_15_c_496_n 4.47528e-19 $X=0.774 $Y=0.162 $X2=0.405
+ $Y2=0.0675
cc_227 N_11_c_415_n N_Q_M14_d 3.73731e-19 $X=1.269 $Y=0.136 $X2=0.783 $Y2=0.0405
cc_228 N_11_c_410_n N_Q_c_454_n 0.00118764f $X=1.08 $Y=0.036 $X2=0.783
+ $Y2=0.1055
cc_229 N_11_c_421_n N_Q_c_454_n 2.62013e-19 $X=1.026 $Y=0.036 $X2=0.783
+ $Y2=0.1055
cc_230 N_11_c_415_n N_Q_M16_d 3.7444e-19 $X=1.269 $Y=0.136 $X2=0.783 $Y2=0.2295
cc_231 N_11_c_415_n N_Q_M31_d 3.8685e-19 $X=1.269 $Y=0.136 $X2=0 $Y2=0
cc_232 N_11_c_418_n N_Q_c_458_n 2.68378e-19 $X=1.026 $Y=0.2025 $X2=0.862
+ $Y2=0.2295
cc_233 N_11_c_432_p N_Q_c_458_n 0.00118419f $X=1.089 $Y=0.167 $X2=0.862
+ $Y2=0.2295
cc_234 N_11_c_415_n N_Q_M33_d 3.87022e-19 $X=1.269 $Y=0.136 $X2=0 $Y2=0
cc_235 N_11_c_415_n N_Q_c_461_n 8.43851e-19 $X=1.269 $Y=0.136 $X2=0.783
+ $Y2=0.105
cc_236 N_11_M15_g N_Q_c_462_n 3.57913e-19 $X=1.215 $Y=0.0675 $X2=0.783 $Y2=0.105
cc_237 N_11_M16_g N_Q_c_462_n 4.61823e-19 $X=1.269 $Y=0.0675 $X2=0.783 $Y2=0.105
cc_238 N_11_c_415_n N_Q_c_464_n 7.60428e-19 $X=1.269 $Y=0.136 $X2=0.936
+ $Y2=0.036
cc_239 N_11_M14_g N_Q_c_465_n 4.31409e-19 $X=1.161 $Y=0.0675 $X2=0.792 $Y2=0.036
cc_240 N_11_c_415_n N_Q_c_465_n 0.00142439f $X=1.269 $Y=0.136 $X2=0.792
+ $Y2=0.036
cc_241 N_11_c_440_p N_Q_c_465_n 5.02824e-19 $X=1.161 $Y=0.136 $X2=0.792
+ $Y2=0.036
cc_242 N_11_M15_g N_Q_c_468_n 3.53956e-19 $X=1.215 $Y=0.0675 $X2=0.864 $Y2=0.036
cc_243 N_11_M16_g N_Q_c_468_n 4.56718e-19 $X=1.269 $Y=0.0675 $X2=0.864 $Y2=0.036
cc_244 N_11_M14_g N_Q_c_470_n 3.94108e-19 $X=1.161 $Y=0.0675 $X2=0.9 $Y2=0.036
cc_245 N_11_c_415_n N_Q_c_470_n 0.00145408f $X=1.269 $Y=0.136 $X2=0.9 $Y2=0.036
cc_246 N_11_c_411_n N_Q_c_470_n 0.0013429f $X=1.08 $Y=0.234 $X2=0.9 $Y2=0.036
cc_247 N_11_c_440_p N_Q_c_470_n 5.18971e-19 $X=1.161 $Y=0.136 $X2=0.9 $Y2=0.036
cc_248 N_11_c_415_n N_Q_c_474_n 4.1631e-19 $X=1.269 $Y=0.136 $X2=0.918 $Y2=0.234
cc_249 N_11_c_410_n N_Q_c_475_n 0.00134363f $X=1.08 $Y=0.036 $X2=0.945 $Y2=0.117
cc_250 N_11_c_449_p N_Q_c_476_n 2.95672e-19 $X=1.143 $Y=0.136 $X2=0.945
+ $Y2=0.171
cc_251 N_11_c_450_p N_Q_c_477_n 0.00134363f $X=1.089 $Y=0.069 $X2=0 $Y2=0
cc_252 N_11_c_451_p N_Q_c_478_n 0.0013429f $X=1.089 $Y=0.225 $X2=0 $Y2=0
cc_253 N_11_c_449_p N_Q_c_478_n 3.06781e-19 $X=1.143 $Y=0.136 $X2=0 $Y2=0

* END of "./DFFHQx4_ASAP7_75t_SRAM.pex.sp.DFFHQX4_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DFFLQNx1_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:25:38 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DFFLQNx1_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DFFLQNx1_ASAP7_75t_SRAM.pex.sp.pex"
* File: DFFLQNx1_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:25:38 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%CLK 2 5 7 12 14 17 VSS
c18 17 VSS 1.44512e-20 $X=0.081 $Y=0.1305
c19 14 VSS 0.00705007f $X=0.081 $Y=0.135
c20 12 VSS 0.00709305f $X=0.082 $Y=0.119
c21 5 VSS 0.00184374f $X=0.081 $Y=0.135
c22 2 VSS 0.0629f $X=0.081 $Y=0.054
r23 16 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r24 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r25 12 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.126
r26 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%4 2 5 7 10 13 16 22 25 28 31 36 43 47 50 52 58
+ 59 60 64 67 74 79 84 88 89 92 96 99 100 101 103 111 124 132 148 VSS
c102 148 VSS 4.19842e-19 $X=0.18 $Y=0.189
c103 147 VSS 1.53928e-19 $X=0.189 $Y=0.189
c104 141 VSS 7.0154e-20 $X=0.03 $Y=0.189
c105 140 VSS 5.9624e-19 $X=0.027 $Y=0.189
c106 124 VSS 6.81413e-19 $X=0.513 $Y=0.18
c107 111 VSS 4.0846e-19 $X=0.351 $Y=0.135
c108 103 VSS 0.00656068f $X=0.513 $Y=0.189
c109 101 VSS 0.00251877f $X=0.29 $Y=0.189
c110 100 VSS 0.00602789f $X=0.229 $Y=0.189
c111 99 VSS 7.60117e-19 $X=0.351 $Y=0.189
c112 96 VSS 4.13996e-19 $X=0.159 $Y=0.189
c113 92 VSS 4.95554e-19 $X=0.033 $Y=0.189
c114 89 VSS 7.37649e-20 $X=0.189 $Y=0.172
c115 88 VSS 5.63427e-19 $X=0.189 $Y=0.164
c116 87 VSS 1.04741e-19 $X=0.189 $Y=0.18
c117 85 VSS 9.32637e-20 $X=0.148 $Y=0.135
c118 84 VSS 9.68735e-19 $X=0.145 $Y=0.135
c119 79 VSS 0.00149077f $X=0.18 $Y=0.135
c120 77 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c121 76 VSS 0.00169428f $X=0.047 $Y=0.234
c122 74 VSS 0.00250477f $X=0.054 $Y=0.234
c123 72 VSS 0.00306385f $X=0.027 $Y=0.234
c124 70 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c125 69 VSS 0.00205521f $X=0.047 $Y=0.036
c126 67 VSS 0.00250477f $X=0.054 $Y=0.036
c127 65 VSS 0.00305101f $X=0.027 $Y=0.036
c128 64 VSS 4.99402e-19 $X=0.018 $Y=0.2125
c129 63 VSS 1.14289e-19 $X=0.018 $Y=0.2
c130 62 VSS 4.86272e-19 $X=0.018 $Y=0.225
c131 60 VSS 0.00271341f $X=0.018 $Y=0.125
c132 59 VSS 9.57865e-19 $X=0.018 $Y=0.07
c133 58 VSS 0.00235012f $X=0.018 $Y=0.18
c134 55 VSS 0.00530434f $X=0.056 $Y=0.216
c135 52 VSS 2.98509e-19 $X=0.071 $Y=0.216
c136 50 VSS 0.00492487f $X=0.056 $Y=0.054
c137 47 VSS 2.98509e-19 $X=0.071 $Y=0.054
c138 43 VSS 0.0585267f $X=0.725 $Y=0.178
c139 36 VSS 0.00123999f $X=0.464 $Y=0.178
c140 28 VSS 0.0616846f $X=0.729 $Y=0.178
c141 25 VSS 1.44609e-19 $X=0.621 $Y=0.178
c142 22 VSS 0.0600171f $X=0.621 $Y=0.0405
c143 16 VSS 0.0602253f $X=0.459 $Y=0.0405
c144 10 VSS 0.0608611f $X=0.351 $Y=0.135
c145 5 VSS 0.00277501f $X=0.135 $Y=0.135
c146 2 VSS 0.0623856f $X=0.135 $Y=0.054
r147 148 149 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.189 $X2=0.1845 $Y2=0.189
r148 147 149 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.189 $X2=0.1845 $Y2=0.189
r149 140 141 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.03 $Y2=0.189
r150 137 140 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.027 $Y2=0.189
r151 131 132 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.351 $Y=0.167 $X2=0.351 $Y2=0.178
r152 123 124 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r153 111 131 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.167
r154 103 124 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r155 100 101 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.189 $X2=0.29 $Y2=0.189
r156 99 132 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.178
r157 98 103 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.513 $Y2=0.189
r158 98 101 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.29 $Y2=0.189
r159 98 99 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.189 $X2=0.351
+ $Y2=0.189
r160 96 148 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.159
+ $Y=0.189 $X2=0.18 $Y2=0.189
r161 95 100 4.75309 $w=1.8e-08 $l=7e-08 $layer=M2 $thickness=3.6e-08 $X=0.159
+ $Y=0.189 $X2=0.229 $Y2=0.189
r162 95 96 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.159 $Y=0.189 $X2=0.159
+ $Y2=0.189
r163 92 141 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.03 $Y2=0.189
r164 91 95 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.159 $Y2=0.189
r165 91 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.189 $X2=0.033
+ $Y2=0.189
r166 88 89 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.172
r167 87 147 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.189
r168 87 89 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.172
r169 86 88 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.164
r170 84 85 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.145
+ $Y=0.135 $X2=0.148 $Y2=0.135
r171 81 84 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.145 $Y2=0.135
r172 79 86 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r173 79 85 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.148 $Y2=0.135
r174 76 77 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r175 74 77 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r176 72 76 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r177 69 70 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r178 67 70 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r179 65 69 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r180 63 64 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r181 62 72 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r182 62 64 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r183 61 137 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.189
r184 61 63 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.2
r185 59 60 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.125
r186 58 137 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.189
r187 58 60 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.125
r188 57 65 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r189 57 59 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r190 55 74 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r191 52 55 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r192 50 67 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r193 47 50 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r194 36 123 39.0385 $w=2.6e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.178 $X2=0.513 $Y2=0.178
r195 28 43 3.07692 $w=2.6e-08 $l=4e-09 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.178 $X2=0.725 $Y2=0.178
r196 28 31 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.178 $X2=0.729 $Y2=0.2295
r197 25 43 82.8571 $w=2.6e-08 $l=1.04e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.725 $Y2=0.178
r198 25 123 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.513 $Y2=0.178
r199 22 25 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0405 $X2=0.621 $Y2=0.178
r200 19 36 3.84615 $w=2.6e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.178 $X2=0.464 $Y2=0.178
r201 16 19 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.178
r202 10 111 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135
+ $X2=0.351 $Y2=0.135
r203 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r204 5 81 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r205 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r206 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%D 2 5 7 12 14 17 VSS
c21 17 VSS 2.32756e-19 $X=0.297 $Y=0.126
c22 14 VSS 0.0072156f $X=0.297 $Y=0.135
c23 12 VSS 0.00703905f $X=0.298 $Y=0.082
c24 5 VSS 0.00200686f $X=0.297 $Y=0.135
c25 2 VSS 0.061556f $X=0.297 $Y=0.0675
r26 16 17 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.126
r27 14 17 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.126
r28 12 16 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.082 $X2=0.297 $Y2=0.106
r29 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r30 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r31 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%6 2 5 7 10 13 15 17 22 25 27 32 34 39 40 42 45
+ 51 53 54 58 63 73 74 76 VSS
c70 76 VSS 7.89434e-19 $X=0.243 $Y=0.2115
c71 74 VSS 9.16337e-19 $X=0.243 $Y=0.126
c72 73 VSS 0.00233088f $X=0.243 $Y=0.106
c73 63 VSS 0.00103743f $X=0.675 $Y=0.135
c74 58 VSS 9.14968e-19 $X=0.405 $Y=0.135
c75 54 VSS 0.00260015f $X=0.601 $Y=0.153
c76 53 VSS 0.00786313f $X=0.527 $Y=0.153
c77 51 VSS 0.00404346f $X=0.675 $Y=0.153
c78 45 VSS 0.00167753f $X=0.243 $Y=0.153
c79 42 VSS 5.5218e-19 $X=0.243 $Y=0.225
c80 40 VSS 0.00181981f $X=0.216 $Y=0.234
c81 39 VSS 0.00525711f $X=0.198 $Y=0.234
c82 34 VSS 0.00482554f $X=0.234 $Y=0.234
c83 33 VSS 0.00200074f $X=0.216 $Y=0.036
c84 32 VSS 0.00545403f $X=0.198 $Y=0.036
c85 27 VSS 0.00500597f $X=0.234 $Y=0.036
c86 25 VSS 0.00648533f $X=0.16 $Y=0.216
c87 20 VSS 0.00602272f $X=0.16 $Y=0.054
c88 13 VSS 0.0021498f $X=0.675 $Y=0.135
c89 10 VSS 0.0585656f $X=0.675 $Y=0.0405
c90 5 VSS 0.00163668f $X=0.405 $Y=0.135
c91 2 VSS 0.058827f $X=0.405 $Y=0.0675
r92 75 76 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.198 $X2=0.243 $Y2=0.2115
r93 73 74 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.106 $X2=0.243 $Y2=0.126
r94 53 54 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.601 $Y2=0.153
r95 51 54 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.675
+ $Y=0.153 $X2=0.601 $Y2=0.153
r96 51 63 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.675 $Y=0.153 $X2=0.675
+ $Y2=0.153
r97 48 53 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.527 $Y2=0.153
r98 48 58 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r99 45 75 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.198
r100 45 74 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.126
r101 44 48 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.405 $Y2=0.153
r102 44 45 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.153 $X2=0.243
+ $Y2=0.153
r103 42 76 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.2115
r104 41 73 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.106
r105 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.216 $Y2=0.234
r106 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.198 $Y2=0.234
r107 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r108 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r109 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.216 $Y2=0.036
r110 29 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r111 27 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r112 27 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r113 25 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r114 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r115 20 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r116 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r117 13 63 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.135 $X2=0.675
+ $Y2=0.135
r118 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2295
r119 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.135
r120 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r121 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2295
r122 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%7 2 5 7 9 10 13 14 17 19 22 29 30 31 33 40 47 48
+ 49 50 51 52 54 55 VSS
c45 56 VSS 3.57489e-19 $X=0.612 $Y=0.09
c46 55 VSS 1.84136e-19 $X=0.603 $Y=0.09
c47 54 VSS 5.96246e-19 $X=0.621 $Y=0.09
c48 52 VSS 4.34894e-19 $X=0.621 $Y=0.214
c49 51 VSS 4.90038e-19 $X=0.621 $Y=0.203
c50 50 VSS 1.59683e-19 $X=0.621 $Y=0.167
c51 49 VSS 2.90654e-19 $X=0.621 $Y=0.165
c52 48 VSS 3.07094e-19 $X=0.621 $Y=0.14
c53 47 VSS 3.66508e-19 $X=0.621 $Y=0.122
c54 46 VSS 3.22511e-19 $X=0.621 $Y=0.225
c55 40 VSS 0.00154565f $X=0.594 $Y=0.054
c56 33 VSS 0.00268134f $X=0.594 $Y=0.234
c57 31 VSS 0.00427376f $X=0.612 $Y=0.234
c58 30 VSS 1.96699e-19 $X=0.583 $Y=0.09
c59 29 VSS 0.00266746f $X=0.581 $Y=0.09
c60 24 VSS 5.17345e-20 $X=0.585 $Y=0.09
c61 22 VSS 0.0179398f $X=0.65 $Y=0.2295
c62 19 VSS 3.14771e-19 $X=0.665 $Y=0.2295
c63 17 VSS 2.5391e-19 $X=0.592 $Y=0.2295
c64 13 VSS 0.0281519f $X=0.594 $Y=0.0405
c65 9 VSS 6.29543e-19 $X=0.611 $Y=0.0405
c66 5 VSS 0.00233073f $X=0.513 $Y=0.09
c67 2 VSS 0.0584396f $X=0.513 $Y=0.0405
r68 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.603
+ $Y=0.09 $X2=0.612 $Y2=0.09
r69 54 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.612 $Y2=0.09
r70 53 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.09 $X2=0.603 $Y2=0.09
r71 51 52 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.214
r72 50 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.203
r73 49 50 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.167
r74 48 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r75 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r76 46 52 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.214
r77 45 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.09
r78 45 47 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.122
r79 38 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.09
r80 38 40 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.054
r81 31 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r82 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r83 29 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.581
+ $Y=0.09 $X2=0.583 $Y2=0.09
r84 26 29 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.09 $X2=0.581 $Y2=0.09
r85 24 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.594 $Y2=0.09
r86 24 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.583 $Y2=0.09
r87 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2295 $X2=0.65 $Y2=0.2295
r88 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.592
+ $Y=0.2295 $X2=0.65 $Y2=0.2295
r89 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r90 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r91 13 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.054 $X2=0.594
+ $Y2=0.054
r92 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.594 $Y2=0.0405
r93 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0405 $X2=0.594 $Y2=0.0405
r94 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.09 $X2=0.513
+ $Y2=0.09
r95 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.09 $X2=0.513 $Y2=0.2295
r96 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.09
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%8 2 5 7 9 14 17 21 22 25 30 31 33 35 36 37 38 39
+ 41 42 43 44 48 50 51 52 53 58 60 61 VSS
c55 64 VSS 2.84134e-19 $X=0.459 $Y=0.131
c56 61 VSS 0.00334468f $X=0.45 $Y=0.036
c57 60 VSS 0.00243127f $X=0.459 $Y=0.036
c58 58 VSS 0.00276391f $X=0.432 $Y=0.036
c59 53 VSS 4.23521e-19 $X=0.5445 $Y=0.131
c60 52 VSS 3.49205e-20 $X=0.522 $Y=0.131
c61 51 VSS 2.00095e-19 $X=0.504 $Y=0.131
c62 50 VSS 0.00133241f $X=0.496 $Y=0.131
c63 48 VSS 5.65734e-19 $X=0.567 $Y=0.131
c64 45 VSS 4.53296e-19 $X=0.459 $Y=0.214
c65 44 VSS 2.01779e-19 $X=0.459 $Y=0.203
c66 43 VSS 6.09344e-21 $X=0.459 $Y=0.167
c67 42 VSS 1.60693e-19 $X=0.459 $Y=0.165
c68 41 VSS 3.22878e-19 $X=0.459 $Y=0.225
c69 39 VSS 2.48018e-19 $X=0.459 $Y=0.114
c70 38 VSS 2.26591e-19 $X=0.459 $Y=0.106
c71 37 VSS 9.45429e-20 $X=0.459 $Y=0.099
c72 36 VSS 8.12259e-19 $X=0.459 $Y=0.081
c73 35 VSS 2.08428e-19 $X=0.459 $Y=0.122
c74 33 VSS 0.00142907f $X=0.434 $Y=0.234
c75 32 VSS 3.66528e-19 $X=0.418 $Y=0.234
c76 31 VSS 0.00146362f $X=0.414 $Y=0.234
c77 30 VSS 0.00368178f $X=0.396 $Y=0.234
c78 25 VSS 0.00389542f $X=0.45 $Y=0.234
c79 24 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c80 21 VSS 0.00348256f $X=0.378 $Y=0.2025
c81 16 VSS 5.70081e-19 $X=0.432 $Y=0.0405
c82 5 VSS 0.00195718f $X=0.567 $Y=0.1305
c83 2 VSS 0.0591962f $X=0.567 $Y=0.0405
r84 61 62 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r85 60 62 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r86 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r87 57 58 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r88 52 53 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r89 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r90 50 51 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.496
+ $Y=0.131 $X2=0.504 $Y2=0.131
r91 48 53 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r92 46 64 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r93 46 50 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.496 $Y2=0.131
r94 44 45 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.203 $X2=0.459 $Y2=0.214
r95 43 44 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.167 $X2=0.459 $Y2=0.203
r96 42 43 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.167
r97 41 45 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r98 40 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r99 40 42 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.165
r100 38 39 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.106 $X2=0.459 $Y2=0.114
r101 37 38 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.099 $X2=0.459 $Y2=0.106
r102 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.099
r103 35 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r104 35 39 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.114
r105 34 60 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r106 34 36 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.081
r107 32 33 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.234 $X2=0.434 $Y2=0.234
r108 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.418 $Y2=0.234
r109 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r110 27 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r111 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r112 25 33 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.434 $Y2=0.234
r113 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r114 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r115 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r116 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r117 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r118 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r119 13 58 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r120 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r121 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r122 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r123 5 48 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.131 $X2=0.567
+ $Y2=0.131
r124 5 7 370.904 $w=2e-08 $l=9.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1305 $X2=0.567 $Y2=0.2295
r125 2 5 337.185 $w=2e-08 $l=9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.1305
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%9 2 5 7 9 14 21 25 26 30 31 32 33 34 39 40 42 43
+ 44 45 46 VSS
c26 46 VSS 1.15795e-19 $X=0.945 $Y=0.171
c27 45 VSS 9.68363e-19 $X=0.945 $Y=0.167
c28 44 VSS 8.8218e-19 $X=0.945 $Y=0.117
c29 43 VSS 0.00183078f $X=0.945 $Y=0.09
c30 42 VSS 0.00237212f $X=0.945 $Y=0.225
c31 40 VSS 0.0018377f $X=0.918 $Y=0.234
c32 39 VSS 0.0056872f $X=0.9 $Y=0.234
c33 34 VSS 0.00462933f $X=0.936 $Y=0.234
c34 33 VSS 0.00189638f $X=0.9 $Y=0.036
c35 32 VSS 0.00352438f $X=0.882 $Y=0.036
c36 31 VSS 0.00146362f $X=0.846 $Y=0.036
c37 30 VSS 0.00508235f $X=0.828 $Y=0.036
c38 26 VSS 0.00226308f $X=0.792 $Y=0.036
c39 25 VSS 0.00657446f $X=0.936 $Y=0.036
c40 21 VSS 0.00122443f $X=0.783 $Y=0.105
c41 17 VSS 0.0048151f $X=0.862 $Y=0.2295
c42 12 VSS 0.00513464f $X=0.862 $Y=0.0405
c43 5 VSS 0.00277722f $X=0.783 $Y=0.1055
c44 2 VSS 0.0590816f $X=0.783 $Y=0.0405
r45 45 46 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.167 $X2=0.945 $Y2=0.171
r46 44 45 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.117 $X2=0.945 $Y2=0.167
r47 43 44 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.09 $X2=0.945 $Y2=0.117
r48 42 46 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.171
r49 41 43 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.09
r50 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.234 $X2=0.918 $Y2=0.234
r51 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.9 $Y2=0.234
r52 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r53 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.918 $Y2=0.234
r54 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r55 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.846 $Y2=0.036
r56 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r57 28 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.846 $Y2=0.036
r58 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.036 $X2=0.828 $Y2=0.036
r59 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r60 25 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.9 $Y2=0.036
r61 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.783 $Y=0.045 $X2=0.792 $Y2=0.036
r62 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.105
r63 17 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234 $X2=0.864
+ $Y2=0.234
r64 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2295 $X2=0.862 $Y2=0.2295
r65 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036 $X2=0.864
+ $Y2=0.036
r66 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.862 $Y2=0.0405
r67 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.105 $X2=0.783
+ $Y2=0.105
r68 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.1055 $X2=0.783 $Y2=0.2295
r69 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.1055
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%10 2 7 10 15 17 18 21 22 23 26 27 32 33 35 37 38
+ 39 40 41 43 44 46 47 50 57 58 66 69 73 76 84 VSS
c59 84 VSS 0.00206151f $X=0.999 $Y=0.135
c60 76 VSS 0.00771499f $X=0.999 $Y=0.153
c61 73 VSS 0.00150008f $X=0.891 $Y=0.153
c62 70 VSS 4.17512e-19 $X=0.837 $Y=0.162
c63 69 VSS 1.52743e-19 $X=0.729 $Y=0.162
c64 66 VSS 0.00370746f $X=0.72 $Y=0.234
c65 65 VSS 0.00266816f $X=0.729 $Y=0.234
c66 58 VSS 4.30636e-19 $X=0.866 $Y=0.162
c67 57 VSS 1.48695e-19 $X=0.85 $Y=0.162
c68 55 VSS 2.75449e-19 $X=0.882 $Y=0.162
c69 50 VSS 3.94906e-19 $X=0.837 $Y=0.135
c70 47 VSS 3.26354e-19 $X=0.792 $Y=0.162
c71 46 VSS 0.00206921f $X=0.774 $Y=0.162
c72 44 VSS 0.00192346f $X=0.828 $Y=0.162
c73 43 VSS 0.00136716f $X=0.729 $Y=0.225
c74 41 VSS 1.52884e-19 $X=0.729 $Y=0.136
c75 40 VSS 9.59255e-20 $X=0.729 $Y=0.119
c76 39 VSS 1.29374e-19 $X=0.729 $Y=0.099
c77 38 VSS 3.52175e-19 $X=0.729 $Y=0.081
c78 37 VSS 2.74133e-19 $X=0.729 $Y=0.153
c79 35 VSS 0.00166816f $X=0.704 $Y=0.036
c80 34 VSS 4.57836e-19 $X=0.688 $Y=0.036
c81 33 VSS 0.00146362f $X=0.684 $Y=0.036
c82 32 VSS 0.00370471f $X=0.666 $Y=0.036
c83 27 VSS 0.00409787f $X=0.72 $Y=0.036
c84 26 VSS 0.00276615f $X=0.702 $Y=0.2295
c85 22 VSS 5.63046e-19 $X=0.719 $Y=0.2295
c86 21 VSS 0.0349304f $X=0.648 $Y=0.0405
c87 17 VSS 5.63046e-19 $X=0.665 $Y=0.0405
c88 13 VSS 0.00246634f $X=0.999 $Y=0.135
c89 10 VSS 0.0656618f $X=0.999 $Y=0.0675
c90 5 VSS 0.00189441f $X=0.837 $Y=0.135
c91 2 VSS 0.0618222f $X=0.837 $Y=0.0405
r92 76 84 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.999 $Y=0.153 $X2=0.999
+ $Y2=0.153
r93 72 76 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.999 $Y2=0.153
r94 72 73 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r95 66 67 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.234 $X2=0.7245 $Y2=0.234
r96 65 67 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.234 $X2=0.7245 $Y2=0.234
r97 62 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.234 $X2=0.72 $Y2=0.234
r98 57 58 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.85
+ $Y=0.162 $X2=0.866 $Y2=0.162
r99 56 70 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.837 $Y2=0.162
r100 56 57 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.85 $Y2=0.162
r101 55 73 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.891 $Y2=0.162
r102 55 58 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.866 $Y2=0.162
r103 48 70 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.162
r104 48 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.135
r105 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.162 $X2=0.792 $Y2=0.162
r106 45 69 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.729 $Y2=0.162
r107 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.774 $Y2=0.162
r108 44 70 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.837 $Y2=0.162
r109 44 47 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.792 $Y2=0.162
r110 43 65 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.225 $X2=0.729 $Y2=0.234
r111 42 69 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.162
r112 42 43 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.225
r113 40 41 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.119 $X2=0.729 $Y2=0.136
r114 39 40 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.099 $X2=0.729 $Y2=0.119
r115 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.081 $X2=0.729 $Y2=0.099
r116 37 69 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.162
r117 37 41 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.136
r118 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.045 $X2=0.729 $Y2=0.081
r119 34 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.036 $X2=0.704 $Y2=0.036
r120 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.688 $Y2=0.036
r121 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.684 $Y2=0.036
r122 29 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.666 $Y2=0.036
r123 27 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.036 $X2=0.729 $Y2=0.045
r124 27 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.704 $Y2=0.036
r125 26 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.234
+ $X2=0.702 $Y2=0.234
r126 23 26 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2295 $X2=0.702 $Y2=0.2295
r127 22 26 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2295 $X2=0.702 $Y2=0.2295
r128 21 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r129 18 21 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0405 $X2=0.648 $Y2=0.0405
r130 17 21 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r131 13 84 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.135 $X2=0.999
+ $Y2=0.135
r132 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.135 $X2=0.999 $Y2=0.2025
r133 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.135
r134 5 50 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.135 $X2=0.837
+ $Y2=0.135
r135 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.2295
r136 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.0405 $X2=0.837 $Y2=0.135
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%QN 1 6 12 14 15 16 19 22 30 VSS
c7 30 VSS 0.00418221f $X=1.044 $Y=0.234
c8 29 VSS 0.00278493f $X=1.053 $Y=0.234
c9 22 VSS 0.00418221f $X=1.044 $Y=0.036
c10 21 VSS 0.00278493f $X=1.053 $Y=0.036
c11 19 VSS 0.00646415f $X=1.026 $Y=0.036
c12 16 VSS 0.00348183f $X=1.053 $Y=0.167
c13 15 VSS 0.00213993f $X=1.053 $Y=0.09
c14 12 VSS 0.00270985f $X=1.053 $Y=0.225
c15 9 VSS 0.00688271f $X=1.024 $Y=0.2025
c16 4 VSS 3.02808e-19 $X=1.024 $Y=0.0675
r17 30 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.234 $X2=1.0485 $Y2=0.234
r18 29 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.234 $X2=1.0485 $Y2=0.234
r19 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.234 $X2=1.044 $Y2=0.234
r20 22 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=1.0485 $Y2=0.036
r21 21 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.036 $X2=1.0485 $Y2=0.036
r22 18 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.036 $X2=1.044 $Y2=0.036
r23 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.036 $X2=1.026
+ $Y2=0.036
r24 15 16 5.22839 $w=1.8e-08 $l=7.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.09 $X2=1.053 $Y2=0.167
r25 14 16 3.80247 $w=1.8e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.223 $X2=1.053 $Y2=0.167
r26 12 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.225 $X2=1.053 $Y2=0.234
r27 12 14 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.225 $X2=1.053 $Y2=0.223
r28 11 21 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.045 $X2=1.053 $Y2=0.036
r29 11 15 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.045 $X2=1.053 $Y2=0.09
r30 9 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.234 $X2=1.026
+ $Y2=0.234
r31 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=1.009
+ $Y=0.2025 $X2=1.024 $Y2=0.2025
r32 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.026
+ $Y=0.0675 $X2=1.026 $Y2=0.036
r33 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.009
+ $Y=0.0675 $X2=1.024 $Y2=0.0675
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%12 1 6 9 VSS
c6 9 VSS 0.0266112f $X=0.38 $Y=0.0675
c7 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c8 4 VSS 3.22674e-19 $X=0.322 $Y=0.0675
r9 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r10 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%13 1 6 9 VSS
c10 9 VSS 0.0209308f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.69239e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%14 1 6 9 VSS
c8 9 VSS 0.0191793f $X=0.758 $Y=0.0405
c9 6 VSS 3.14771e-19 $X=0.773 $Y=0.0405
c10 4 VSS 2.61968e-19 $X=0.7 $Y=0.0405
r11 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r12 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.7
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r13 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.685
+ $Y=0.0405 $X2=0.7 $Y2=0.0405
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%15 1 2 VSS
c0 1 VSS 0.00225696f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%16 1 2 VSS
c1 1 VSS 0.00201018f $X=0.341 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends

.subckt PM_DFFLQNX1_ASAP7_75T_SRAM%17 1 2 VSS
c0 1 VSS 0.00219822f $X=0.773 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2295 $X2=0.739 $Y2=0.2295
.ends


* END of "./DFFLQNx1_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DFFLQNx1_ASAP7_75t_SRAM  VSS VDD CLK D QN
* 
* QN	QN
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_12_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_6_M3_g N_12_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_15_M4_d N_4_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_15_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_10_M7_d N_4_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.611
+ $Y=0.027
M8 N_14_M8_d N_6_M8_g N_10_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M9 VSS N_9_M9_g N_14_M9_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_9_M10_d N_10_M10_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.027
M11 N_QN_M11_d N_10_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M12 VDD N_CLK_M12_g N_4_M12_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M13 N_6_M13_d N_4_M13_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M14 N_16_M14_d N_D_M14_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M15 N_8_M15_d N_4_M15_g N_16_M15_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M16 N_13_M16_d N_6_M16_g N_8_M16_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M17 VDD N_7_M17_g N_13_M17_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M18 N_7_M18_d N_8_M18_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M19 N_10_M19_d N_6_M19_g N_7_M19_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.665 $Y=0.216
M20 N_17_M20_d N_4_M20_g N_10_M20_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.719 $Y=0.216
M21 VDD N_9_M21_g N_17_M21_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M22 N_9_M22_d N_10_M22_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.216
M23 N_QN_M23_d N_10_M23_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
*
* 
* .include "DFFLQNx1_ASAP7_75t_SRAM.pex.sp.DFFLQNX1_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DFFLQNx1_ASAP7_75t_SRAM.pex.sp.DFFLQNX1_ASAP7_75T_SRAM.pxi"
* File: DFFLQNx1_ASAP7_75t_SRAM.pex.sp.DFFLQNX1_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:25:38 2017
* 
x_PM_DFFLQNX1_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M12_g CLK N_CLK_c_4_p
+ N_CLK_c_10_p VSS PM_DFFLQNX1_ASAP7_75T_SRAM%CLK
x_PM_DFFLQNX1_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_20_n N_4_M13_g N_4_c_34_p N_4_M15_g
+ N_4_M4_g N_4_M7_g N_4_c_77_p N_4_c_43_p N_4_M20_g N_4_c_89_p N_4_c_44_p
+ N_4_M0_s N_4_c_21_n N_4_M12_s N_4_c_22_n N_4_c_23_n N_4_c_24_n N_4_c_25_n
+ N_4_c_26_n N_4_c_27_n N_4_c_47_p N_4_c_28_n N_4_c_29_n N_4_c_30_n N_4_c_31_n
+ N_4_c_32_n N_4_c_58_p N_4_c_33_n N_4_c_36_p N_4_c_37_p N_4_c_38_p N_4_c_61_p
+ N_4_c_94_p N_4_c_46_p VSS PM_DFFLQNX1_ASAP7_75T_SRAM%4
x_PM_DFFLQNX1_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_122_n N_D_M14_g D N_D_c_123_n
+ N_D_c_133_p VSS PM_DFFLQNX1_ASAP7_75T_SRAM%D
x_PM_DFFLQNX1_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_147_n N_6_M16_g N_6_M8_g N_6_c_151_n
+ N_6_M19_g N_6_M1_d N_6_M13_d N_6_c_152_n N_6_c_172_n N_6_c_142_n N_6_c_154_n
+ N_6_c_143_n N_6_c_158_n N_6_c_174_n N_6_c_159_n N_6_c_161_n N_6_c_162_n
+ N_6_c_183_p N_6_c_168_n N_6_c_170_n N_6_c_144_n N_6_c_180_n N_6_c_181_n VSS
+ PM_DFFLQNX1_ASAP7_75T_SRAM%6
x_PM_DFFLQNX1_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_237_p N_7_M17_g N_7_M7_s N_7_M6_d
+ N_7_c_216_n N_7_M18_d N_7_c_217_n N_7_M19_s N_7_c_219_n N_7_c_235_p
+ N_7_c_228_n N_7_c_255_p N_7_c_229_n N_7_c_236_p N_7_c_221_n N_7_c_240_p
+ N_7_c_222_n N_7_c_223_n N_7_c_224_n N_7_c_253_p N_7_c_226_n N_7_c_233_n VSS
+ PM_DFFLQNX1_ASAP7_75T_SRAM%7
x_PM_DFFLQNX1_ASAP7_75T_SRAM%8 N_8_M6_g N_8_c_280_n N_8_M18_g N_8_M3_d N_8_M4_s
+ N_8_M15_d N_8_c_260_n N_8_M16_s N_8_c_308_p N_8_c_262_n N_8_c_283_n
+ N_8_c_309_p N_8_c_285_n N_8_c_263_n N_8_c_264_n N_8_c_298_n N_8_c_286_n
+ N_8_c_310_p N_8_c_265_n N_8_c_266_n N_8_c_268_n N_8_c_299_n N_8_c_272_n
+ N_8_c_300_n N_8_c_273_n N_8_c_275_n N_8_c_291_n N_8_c_303_n N_8_c_278_n VSS
+ PM_DFFLQNX1_ASAP7_75T_SRAM%8
x_PM_DFFLQNX1_ASAP7_75T_SRAM%9 N_9_M9_g N_9_c_318_p N_9_M21_g N_9_M10_d N_9_M22_d
+ N_9_c_317_p N_9_c_329_p N_9_c_316_p N_9_c_321_p N_9_c_315_p N_9_c_325_p
+ N_9_c_327_p N_9_c_336_p N_9_c_326_p N_9_c_330_p N_9_c_320_p N_9_c_334_p
+ N_9_c_332_p N_9_c_328_p N_9_c_333_p VSS PM_DFFLQNX1_ASAP7_75T_SRAM%9
x_PM_DFFLQNX1_ASAP7_75T_SRAM%10 N_10_M10_g N_10_M22_g N_10_M11_g N_10_M23_g
+ N_10_M8_s N_10_M7_d N_10_c_339_n N_10_M20_s N_10_M19_d N_10_c_341_n
+ N_10_c_372_n N_10_c_352_n N_10_c_353_n N_10_c_394_p N_10_c_355_n N_10_c_364_n
+ N_10_c_342_n N_10_c_343_n N_10_c_344_n N_10_c_345_n N_10_c_377_n N_10_c_347_n
+ N_10_c_378_n N_10_c_380_n N_10_c_381_n N_10_c_382_n N_10_c_348_n N_10_c_349_n
+ N_10_c_383_n N_10_c_357_n N_10_c_388_n VSS PM_DFFLQNX1_ASAP7_75T_SRAM%10
x_PM_DFFLQNX1_ASAP7_75T_SRAM%QN N_QN_M11_d N_QN_M23_d N_QN_c_397_n QN N_QN_c_398_n
+ N_QN_c_401_n N_QN_c_403_n N_QN_c_399_n N_QN_c_400_n VSS
+ PM_DFFLQNX1_ASAP7_75T_SRAM%QN
x_PM_DFFLQNX1_ASAP7_75T_SRAM%12 N_12_M2_d N_12_M3_s N_12_c_404_n VSS
+ PM_DFFLQNX1_ASAP7_75T_SRAM%12
x_PM_DFFLQNX1_ASAP7_75T_SRAM%13 N_13_M16_d N_13_M17_s N_13_c_411_n VSS
+ PM_DFFLQNX1_ASAP7_75T_SRAM%13
x_PM_DFFLQNX1_ASAP7_75T_SRAM%14 N_14_M8_d N_14_M9_s N_14_c_420_n VSS
+ PM_DFFLQNX1_ASAP7_75T_SRAM%14
x_PM_DFFLQNX1_ASAP7_75T_SRAM%15 N_15_M5_s N_15_M4_d VSS PM_DFFLQNX1_ASAP7_75T_SRAM%15
x_PM_DFFLQNX1_ASAP7_75T_SRAM%16 N_16_M15_s N_16_M14_d VSS
+ PM_DFFLQNX1_ASAP7_75T_SRAM%16
x_PM_DFFLQNX1_ASAP7_75T_SRAM%17 N_17_M21_s N_17_M20_d VSS
+ PM_DFFLQNX1_ASAP7_75T_SRAM%17
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_CLK_c_2_p N_4_c_20_n 0.00124017f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 CLK N_4_c_21_n 3.57152e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_4 N_CLK_c_4_p N_4_c_22_n 0.00206543f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.18
cc_5 CLK N_4_c_23_n 2.75361e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.07
cc_6 CLK N_4_c_24_n 0.00206543f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.125
cc_7 N_CLK_c_4_p N_4_c_25_n 2.75361e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2125
cc_8 CLK N_4_c_26_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_4_p N_4_c_27_n 5.03453e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_10_p N_4_c_28_n 8.76278e-19 $X=0.081 $Y=0.1305 $X2=0.145 $Y2=0.135
cc_11 N_CLK_c_4_p N_4_c_29_n 3.53816e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.164
cc_12 N_CLK_c_4_p N_4_c_30_n 6.15177e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.172
cc_13 N_CLK_c_4_p N_4_c_31_n 0.00138527f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.189
cc_14 N_CLK_c_4_p N_4_c_32_n 9.65218e-19 $X=0.081 $Y=0.135 $X2=0.159 $Y2=0.189
cc_15 N_CLK_c_4_p N_4_c_33_n 0.00167589f $X=0.081 $Y=0.135 $X2=0.229 $Y2=0.189
cc_16 CLK N_6_c_142_n 6.45949e-19 $X=0.082 $Y=0.119 $X2=0 $Y2=0
cc_17 N_CLK_c_4_p N_6_c_143_n 6.54444e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_18 CLK N_6_c_144_n 6.20748e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.234
cc_19 N_4_c_34_p N_D_M2_g 0.00341068f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.054
cc_20 N_4_c_34_p N_D_c_122_n 0.0010364f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 N_4_c_36_p N_D_c_123_n 2.29805e-19 $X=0.29 $Y=0.189 $X2=0.081 $Y2=0.135
cc_22 N_4_c_37_p N_D_c_123_n 0.00102387f $X=0.513 $Y=0.189 $X2=0.081 $Y2=0.135
cc_23 N_4_c_38_p N_D_c_123_n 0.00337064f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_4_c_34_p N_6_M3_g 0.00355599f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.054
cc_25 N_4_M4_g N_6_M3_g 0.00355599f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_26 N_4_c_34_p N_6_c_147_n 0.00103664f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_27 N_4_M7_g N_6_M8_g 0.00355599f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_28 N_4_c_43_p N_6_M8_g 0.00355599f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_29 N_4_c_44_p N_6_M8_g 0.00250257f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_30 N_4_c_44_p N_6_c_151_n 0.00180656f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_31 N_4_c_46_p N_6_c_152_n 0.00135022f $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_32 N_4_c_47_p N_6_c_142_n 0.0010851f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_33 N_4_c_36_p N_6_c_154_n 4.24027e-19 $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_34 N_4_c_32_n N_6_c_143_n 0.00285029f $X=0.159 $Y=0.189 $X2=0 $Y2=0
cc_35 N_4_c_33_n N_6_c_143_n 6.46981e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_36 N_4_c_46_p N_6_c_143_n 2.904e-19 $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_37 N_4_c_33_n N_6_c_158_n 4.24027e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_38 N_4_c_47_p N_6_c_159_n 0.00351854f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_39 N_4_c_36_p N_6_c_159_n 0.00102595f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_40 N_4_c_44_p N_6_c_161_n 6.40799e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_41 N_4_c_44_p N_6_c_162_n 0.00187197f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_42 N_4_c_29_n N_6_c_162_n 3.52457e-19 $X=0.189 $Y=0.164 $X2=0 $Y2=0
cc_43 N_4_c_58_p N_6_c_162_n 2.46239e-19 $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_44 N_4_c_36_p N_6_c_162_n 0.0253778f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_45 N_4_c_38_p N_6_c_162_n 0.00115493f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_61_p N_6_c_162_n 2.81476e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_47 N_4_c_37_p N_6_c_168_n 2.98936e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_48 N_4_c_38_p N_6_c_168_n 0.00170246f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_49 N_4_c_44_p N_6_c_170_n 0.00124003f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_50 N_4_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_51 N_4_M7_g N_7_M5_g 2.13359e-19 $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_52 N_4_c_44_p N_7_M5_g 0.00205997f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_53 N_4_c_61_p N_7_M5_g 3.15189e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_54 N_4_c_44_p N_7_c_216_n 5.49754e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_55 N_4_c_44_p N_7_c_217_n 2.12581e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.1305
cc_56 N_4_c_44_p N_7_M19_s 2.50995e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_57 N_4_M7_g N_7_c_219_n 0.00200065f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_58 N_4_c_44_p N_7_c_219_n 0.00322783f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_59 N_4_M7_g N_7_c_221_n 3.04073e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_60 N_4_M7_g N_7_c_222_n 2.22997e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_61 N_4_c_61_p N_7_c_223_n 5.74745e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_62 N_4_c_77_p N_7_c_224_n 0.00193027f $X=0.621 $Y=0.178 $X2=0 $Y2=0
cc_63 N_4_c_44_p N_7_c_224_n 0.00189849f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_64 N_4_M7_g N_7_c_226_n 3.8308e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_65 N_4_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_66 N_4_M7_g N_8_M6_g 0.00341068f $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_67 N_4_c_44_p N_8_M6_g 0.00302156f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_68 N_4_c_37_p N_8_c_260_n 3.15319e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_69 N_4_c_38_p N_8_c_260_n 0.00136448f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_70 N_4_c_37_p N_8_c_262_n 0.00161272f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_71 N_4_M4_g N_8_c_263_n 3.80535e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_72 N_4_M4_g N_8_c_264_n 2.08362e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_73 N_4_M4_g N_8_c_265_n 2.27303e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_74 N_4_c_89_p N_8_c_266_n 4.73369e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_75 N_4_c_61_p N_8_c_266_n 0.00174159f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_76 N_4_c_89_p N_8_c_268_n 0.0017128f $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_77 N_4_c_44_p N_8_c_268_n 5.88593e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_78 N_4_c_37_p N_8_c_268_n 0.00102123f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_79 N_4_c_94_p N_8_c_268_n 3.42482e-19 $X=0.351 $Y=0.178 $X2=0 $Y2=0
cc_80 N_4_c_44_p N_8_c_272_n 8.16411e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_81 N_4_c_44_p N_8_c_273_n 3.32592e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_82 N_4_c_61_p N_8_c_273_n 8.9822e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_83 N_4_c_44_p N_8_c_275_n 5.02733e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_84 N_4_c_43_p N_9_M9_g 0.00341068f $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_85 N_4_c_43_p N_10_M10_g 2.13359e-19 $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_86 N_4_c_44_p N_10_c_339_n 8.27829e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_87 N_4_c_44_p N_10_M20_s 3.37661e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_88 N_4_c_44_p N_10_c_341_n 0.00145657f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_89 N_4_c_43_p N_10_c_342_n 2.71526e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_90 N_4_c_43_p N_10_c_343_n 2.11119e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_91 N_4_c_43_p N_10_c_344_n 2.58771e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_92 N_4_c_43_p N_10_c_345_n 0.00229157f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_93 N_4_c_44_p N_10_c_345_n 7.89371e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_94 N_4_c_43_p N_10_c_347_n 4.55487e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_95 N_4_c_44_p N_10_c_348_n 4.45535e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_96 N_4_c_43_p N_10_c_349_n 5.68093e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_97 N_4_c_44_p N_10_c_349_n 2.2968e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_98 N_4_c_34_p N_12_c_404_n 0.00526068f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_99 N_4_c_44_p N_13_M17_s 2.36286e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.216
cc_100 N_4_M4_g N_13_c_411_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_101 N_4_c_89_p N_13_c_411_n 5.41258e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_102 N_4_c_44_p N_13_c_411_n 0.00230928f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_103 N_4_c_37_p N_13_c_411_n 7.09553e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_104 N_4_c_43_p N_14_c_420_n 0.00198387f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_105 N_4_c_44_p N_14_c_420_n 4.51352e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_106 N_D_M2_g N_6_M3_g 2.82885e-19 $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_107 D N_6_c_172_n 0.00115224f $X=0.298 $Y=0.082 $X2=0.729 $Y2=0.178
cc_108 N_D_c_123_n N_6_c_154_n 0.00115224f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_109 N_D_c_123_n N_6_c_174_n 0.00115224f $X=0.297 $Y=0.135 $X2=0.725 $Y2=0.178
cc_110 N_D_c_123_n N_6_c_159_n 0.00124565f $X=0.297 $Y=0.135 $X2=0.729 $Y2=0.178
cc_111 D N_6_c_162_n 2.27807e-19 $X=0.298 $Y=0.082 $X2=0.056 $Y2=0.216
cc_112 N_D_c_123_n N_6_c_162_n 9.62099e-19 $X=0.297 $Y=0.135 $X2=0.056 $Y2=0.216
cc_113 N_D_c_133_p N_6_c_168_n 4.3159e-19 $X=0.297 $Y=0.126 $X2=0.018 $Y2=0.18
cc_114 D N_6_c_144_n 0.00115224f $X=0.298 $Y=0.082 $X2=0.054 $Y2=0.234
cc_115 N_D_c_133_p N_6_c_180_n 0.00115224f $X=0.297 $Y=0.126 $X2=0.054 $Y2=0.234
cc_116 N_D_c_123_n N_6_c_181_n 0.00115224f $X=0.297 $Y=0.135 $X2=0.047 $Y2=0.234
cc_117 N_D_c_123_n N_8_c_260_n 3.88702e-19 $X=0.297 $Y=0.135 $X2=0.621
+ $Y2=0.0405
cc_118 N_D_c_123_n N_8_c_262_n 8.77202e-19 $X=0.297 $Y=0.135 $X2=0.729
+ $Y2=0.2295
cc_119 D N_8_c_278_n 2.04306e-19 $X=0.298 $Y=0.082 $X2=0.018 $Y2=0.198
cc_120 D N_12_c_404_n 0.00430488f $X=0.298 $Y=0.082 $X2=0.351 $Y2=0.135
cc_121 N_D_c_123_n N_16_M15_s 3.05674e-19 $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_122 N_6_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_123 N_6_c_183_p N_7_c_228_n 2.96121e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_124 N_6_c_161_n N_7_c_229_n 2.61213e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_125 N_6_c_183_p N_7_c_229_n 2.61213e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_126 N_6_c_170_n N_7_c_221_n 0.00327797f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_127 N_6_c_161_n N_7_c_222_n 0.00115177f $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_128 N_6_c_161_n N_7_c_233_n 2.96121e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_129 N_6_M8_g N_8_M6_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_130 N_6_c_151_n N_8_c_280_n 4.12331e-19 $X=0.675 $Y=0.135 $X2=0.081 $Y2=0.135
cc_131 N_6_c_183_p N_8_c_280_n 2.64012e-19 $X=0.601 $Y=0.153 $X2=0.081 $Y2=0.135
cc_132 N_6_c_168_n N_8_c_260_n 2.25088e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_133 N_6_M3_g N_8_c_283_n 3.49806e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_134 N_6_c_168_n N_8_c_283_n 3.83282e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_135 N_6_c_168_n N_8_c_285_n 9.70699e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_136 N_6_c_168_n N_8_c_286_n 9.70699e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_137 N_6_c_162_n N_8_c_265_n 0.00118282f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_138 N_6_c_168_n N_8_c_265_n 0.00106411f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_139 N_6_c_162_n N_8_c_272_n 0.00138951f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_140 N_6_c_183_p N_8_c_275_n 0.00138951f $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_141 N_6_c_162_n N_8_c_291_n 2.54113e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_142 N_6_c_162_n N_8_c_278_n 3.92135e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_143 N_6_M8_g N_9_M9_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_144 N_6_c_161_n N_10_c_339_n 2.24654e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_145 N_6_c_161_n N_10_c_352_n 5.06919e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_146 N_6_M8_g N_10_c_353_n 3.43727e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_147 N_6_c_170_n N_10_c_353_n 5.96743e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_148 N_6_c_161_n N_10_c_355_n 2.34004e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_149 N_6_c_170_n N_10_c_343_n 0.00329725f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_150 N_6_c_161_n N_10_c_357_n 2.83245e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_151 N_6_c_162_n N_12_c_404_n 8.35084e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_152 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_153 N_7_c_235_p N_8_M6_g 3.91159e-19 $X=0.581 $Y=0.09 $X2=0.135 $Y2=0.054
cc_154 N_7_c_236_p N_8_c_263_n 2.10569e-19 $X=0.594 $Y=0.054 $X2=0.464 $Y2=0.178
cc_155 N_7_c_237_p N_8_c_264_n 3.19692e-19 $X=0.513 $Y=0.09 $X2=0 $Y2=0
cc_156 N_7_c_235_p N_8_c_264_n 0.00107929f $X=0.581 $Y=0.09 $X2=0 $Y2=0
cc_157 N_7_c_221_n N_8_c_298_n 2.4251e-19 $X=0.621 $Y=0.122 $X2=0 $Y2=0
cc_158 N_7_c_240_p N_8_c_299_n 9.84729e-19 $X=0.621 $Y=0.14 $X2=0.056 $Y2=0.054
cc_159 N_7_c_235_p N_8_c_300_n 0.00507595f $X=0.581 $Y=0.09 $X2=0 $Y2=0
cc_160 N_7_M5_g N_8_c_273_n 3.12986e-19 $X=0.513 $Y=0.0405 $X2=0.071 $Y2=0.216
cc_161 N_7_c_237_p N_8_c_291_n 5.2508e-19 $X=0.513 $Y=0.09 $X2=0.018 $Y2=0.18
cc_162 N_7_c_236_p N_8_c_303_n 2.10569e-19 $X=0.594 $Y=0.054 $X2=0.018 $Y2=0.125
cc_163 N_7_c_216_n N_10_c_339_n 0.00328169f $X=0.594 $Y=0.0405 $X2=0.621
+ $Y2=0.0405
cc_164 N_7_c_236_p N_10_c_339_n 3.00222e-19 $X=0.594 $Y=0.054 $X2=0.621
+ $Y2=0.0405
cc_165 N_7_c_226_n N_10_c_339_n 2.70684e-19 $X=0.621 $Y=0.09 $X2=0.621
+ $Y2=0.0405
cc_166 N_7_c_219_n N_10_c_341_n 0.00222825f $X=0.65 $Y=0.2295 $X2=0 $Y2=0
cc_167 N_7_c_216_n N_10_c_352_n 3.50513e-19 $X=0.594 $Y=0.0405 $X2=0 $Y2=0
cc_168 N_7_c_236_p N_10_c_352_n 5.0339e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_169 N_7_c_236_p N_10_c_364_n 2.21141e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_170 N_7_c_226_n N_10_c_342_n 4.36168e-19 $X=0.621 $Y=0.09 $X2=0 $Y2=0
cc_171 N_7_c_253_p N_10_c_345_n 4.36168e-19 $X=0.621 $Y=0.214 $X2=0.725
+ $Y2=0.178
cc_172 N_7_c_219_n N_10_c_348_n 3.64454e-19 $X=0.65 $Y=0.2295 $X2=0.054
+ $Y2=0.036
cc_173 N_7_c_255_p N_10_c_348_n 4.86017e-19 $X=0.612 $Y=0.234 $X2=0.054
+ $Y2=0.036
cc_174 N_7_c_224_n N_10_c_349_n 4.36168e-19 $X=0.621 $Y=0.203 $X2=0.047
+ $Y2=0.036
cc_175 N_8_c_260_n N_12_c_404_n 0.00119636f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.135
cc_176 N_8_c_291_n N_12_c_404_n 0.00390673f $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_177 N_8_c_278_n N_12_c_404_n 4.41747e-19 $X=0.45 $Y=0.036 $X2=0.351 $Y2=0.135
cc_178 N_8_c_260_n N_13_c_411_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.135
cc_179 N_8_c_308_p N_13_c_411_n 0.00209454f $X=0.45 $Y=0.234 $X2=0.351 $Y2=0.135
cc_180 N_8_c_309_p N_13_c_411_n 0.0013184f $X=0.434 $Y=0.234 $X2=0.351 $Y2=0.135
cc_181 N_8_c_310_p N_13_c_411_n 0.00116187f $X=0.459 $Y=0.225 $X2=0.351
+ $Y2=0.135
cc_182 N_8_c_291_n N_13_c_411_n 5.72158e-19 $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_183 N_9_M9_g N_10_M10_g 0.00268443f $X=0.783 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_184 N_9_c_315_p N_10_M10_g 3.74489e-19 $X=0.846 $Y=0.036 $X2=0.135 $Y2=0.054
cc_185 N_9_c_316_p N_10_c_372_n 0.00141609f $X=0.792 $Y=0.036 $X2=0.729
+ $Y2=0.178
cc_186 N_9_c_317_p N_10_c_364_n 0.00141609f $X=0.783 $Y=0.105 $X2=0 $Y2=0
cc_187 N_9_c_318_p N_10_c_342_n 3.34766e-19 $X=0.783 $Y=0.1055 $X2=0 $Y2=0
cc_188 N_9_c_317_p N_10_c_342_n 0.00141609f $X=0.783 $Y=0.105 $X2=0 $Y2=0
cc_189 N_9_c_320_p N_10_c_345_n 2.41112e-19 $X=0.945 $Y=0.225 $X2=0.725
+ $Y2=0.178
cc_190 N_9_c_321_p N_10_c_377_n 2.65946e-19 $X=0.828 $Y=0.036 $X2=0 $Y2=0
cc_191 N_9_M9_g N_10_c_378_n 6.3699e-19 $X=0.783 $Y=0.0405 $X2=0.071 $Y2=0.054
cc_192 N_9_c_317_p N_10_c_378_n 9.10342e-19 $X=0.783 $Y=0.105 $X2=0.071
+ $Y2=0.054
cc_193 N_9_c_315_p N_10_c_380_n 4.40983e-19 $X=0.846 $Y=0.036 $X2=0.056
+ $Y2=0.054
cc_194 N_9_c_325_p N_10_c_381_n 5.181e-19 $X=0.882 $Y=0.036 $X2=0.018 $Y2=0.045
cc_195 N_9_c_326_p N_10_c_382_n 0.00149072f $X=0.9 $Y=0.234 $X2=0.018 $Y2=0.18
cc_196 N_9_c_327_p N_10_c_383_n 4.52584e-19 $X=0.9 $Y=0.036 $X2=0.054 $Y2=0.234
cc_197 N_9_c_328_p N_10_c_383_n 0.00299476f $X=0.945 $Y=0.167 $X2=0.054
+ $Y2=0.234
cc_198 N_9_c_329_p N_10_c_357_n 2.40515e-19 $X=0.936 $Y=0.036 $X2=0.047
+ $Y2=0.234
cc_199 N_9_c_330_p N_10_c_357_n 7.44774e-19 $X=0.918 $Y=0.234 $X2=0.047
+ $Y2=0.234
cc_200 N_9_c_328_p N_10_c_357_n 9.28741e-19 $X=0.945 $Y=0.167 $X2=0.047
+ $Y2=0.234
cc_201 N_9_c_332_p N_10_c_388_n 0.00323003f $X=0.945 $Y=0.117 $X2=0.145
+ $Y2=0.135
cc_202 N_9_c_333_p N_QN_c_397_n 3.5495e-19 $X=0.945 $Y=0.171 $X2=0.351
+ $Y2=0.2025
cc_203 N_9_c_334_p N_QN_c_398_n 3.5495e-19 $X=0.945 $Y=0.09 $X2=0.459 $Y2=0.0405
cc_204 N_9_c_329_p N_QN_c_399_n 4.40179e-19 $X=0.936 $Y=0.036 $X2=0.621
+ $Y2=0.0405
cc_205 N_9_c_336_p N_QN_c_400_n 4.34861e-19 $X=0.936 $Y=0.234 $X2=0.729
+ $Y2=0.2295
cc_206 N_9_c_316_p N_14_c_420_n 7.33799e-19 $X=0.792 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_207 N_10_c_357_n N_QN_c_401_n 2.28166e-19 $X=0.999 $Y=0.153 $X2=0.459
+ $Y2=0.0405
cc_208 N_10_c_388_n N_QN_c_401_n 0.0033202f $X=0.999 $Y=0.135 $X2=0.459
+ $Y2=0.0405
cc_209 N_10_c_388_n N_QN_c_403_n 5.42522e-19 $X=0.999 $Y=0.135 $X2=0.459
+ $Y2=0.178
cc_210 N_10_c_339_n N_14_c_420_n 0.00182708f $X=0.648 $Y=0.0405 $X2=0.351
+ $Y2=0.135
cc_211 N_10_c_372_n N_14_c_420_n 0.00205226f $X=0.72 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_212 N_10_c_394_p N_14_c_420_n 0.0013184f $X=0.704 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_213 N_10_c_364_n N_14_c_420_n 0.00103589f $X=0.729 $Y=0.081 $X2=0.351
+ $Y2=0.135
cc_214 N_10_c_347_n N_14_c_420_n 4.02739e-19 $X=0.774 $Y=0.162 $X2=0.351
+ $Y2=0.135

* END of "./DFFLQNx1_ASAP7_75t_SRAM.pex.sp.DFFLQNX1_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DFFLQNx2_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:26:01 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DFFLQNx2_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DFFLQNx2_ASAP7_75t_SRAM.pex.sp.pex"
* File: DFFLQNx2_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:26:01 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%CLK 2 5 7 12 14 17 VSS
c18 17 VSS 1.44512e-20 $X=0.081 $Y=0.1305
c19 14 VSS 0.00705007f $X=0.081 $Y=0.135
c20 12 VSS 0.00709305f $X=0.082 $Y=0.119
c21 5 VSS 0.00184374f $X=0.081 $Y=0.135
c22 2 VSS 0.0629f $X=0.081 $Y=0.054
r23 16 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r24 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r25 12 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.126
r26 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%4 2 5 7 10 13 16 22 25 28 31 36 43 47 50 52 58
+ 59 60 64 67 74 79 84 88 89 92 96 99 100 101 103 111 124 132 148 VSS
c102 148 VSS 4.19842e-19 $X=0.18 $Y=0.189
c103 147 VSS 1.53928e-19 $X=0.189 $Y=0.189
c104 141 VSS 7.0154e-20 $X=0.03 $Y=0.189
c105 140 VSS 5.9624e-19 $X=0.027 $Y=0.189
c106 124 VSS 6.81413e-19 $X=0.513 $Y=0.18
c107 111 VSS 4.0846e-19 $X=0.351 $Y=0.135
c108 103 VSS 0.00656068f $X=0.513 $Y=0.189
c109 101 VSS 0.00251877f $X=0.29 $Y=0.189
c110 100 VSS 0.00602789f $X=0.229 $Y=0.189
c111 99 VSS 7.60117e-19 $X=0.351 $Y=0.189
c112 96 VSS 4.13996e-19 $X=0.159 $Y=0.189
c113 92 VSS 4.95554e-19 $X=0.033 $Y=0.189
c114 89 VSS 7.37649e-20 $X=0.189 $Y=0.172
c115 88 VSS 5.63427e-19 $X=0.189 $Y=0.164
c116 87 VSS 1.04741e-19 $X=0.189 $Y=0.18
c117 85 VSS 9.32637e-20 $X=0.148 $Y=0.135
c118 84 VSS 9.68735e-19 $X=0.145 $Y=0.135
c119 79 VSS 0.00149077f $X=0.18 $Y=0.135
c120 77 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c121 76 VSS 0.00169428f $X=0.047 $Y=0.234
c122 74 VSS 0.00250477f $X=0.054 $Y=0.234
c123 72 VSS 0.00306385f $X=0.027 $Y=0.234
c124 70 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c125 69 VSS 0.00205521f $X=0.047 $Y=0.036
c126 67 VSS 0.00250477f $X=0.054 $Y=0.036
c127 65 VSS 0.00305101f $X=0.027 $Y=0.036
c128 64 VSS 4.99402e-19 $X=0.018 $Y=0.2125
c129 63 VSS 1.14289e-19 $X=0.018 $Y=0.2
c130 62 VSS 4.86272e-19 $X=0.018 $Y=0.225
c131 60 VSS 0.00271341f $X=0.018 $Y=0.125
c132 59 VSS 9.57865e-19 $X=0.018 $Y=0.07
c133 58 VSS 0.00235012f $X=0.018 $Y=0.18
c134 55 VSS 0.00530434f $X=0.056 $Y=0.216
c135 52 VSS 2.98509e-19 $X=0.071 $Y=0.216
c136 50 VSS 0.00492487f $X=0.056 $Y=0.054
c137 47 VSS 2.98509e-19 $X=0.071 $Y=0.054
c138 43 VSS 0.0585267f $X=0.725 $Y=0.178
c139 36 VSS 0.00123999f $X=0.464 $Y=0.178
c140 28 VSS 0.0616846f $X=0.729 $Y=0.178
c141 25 VSS 1.44609e-19 $X=0.621 $Y=0.178
c142 22 VSS 0.0600171f $X=0.621 $Y=0.0405
c143 16 VSS 0.0602253f $X=0.459 $Y=0.0405
c144 10 VSS 0.0608611f $X=0.351 $Y=0.135
c145 5 VSS 0.00277501f $X=0.135 $Y=0.135
c146 2 VSS 0.0623856f $X=0.135 $Y=0.054
r147 148 149 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.189 $X2=0.1845 $Y2=0.189
r148 147 149 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.189 $X2=0.1845 $Y2=0.189
r149 140 141 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.03 $Y2=0.189
r150 137 140 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.027 $Y2=0.189
r151 131 132 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.351 $Y=0.167 $X2=0.351 $Y2=0.178
r152 123 124 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r153 111 131 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.167
r154 103 124 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r155 100 101 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.189 $X2=0.29 $Y2=0.189
r156 99 132 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.178
r157 98 103 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.513 $Y2=0.189
r158 98 101 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.29 $Y2=0.189
r159 98 99 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.189 $X2=0.351
+ $Y2=0.189
r160 96 148 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.159
+ $Y=0.189 $X2=0.18 $Y2=0.189
r161 95 100 4.75309 $w=1.8e-08 $l=7e-08 $layer=M2 $thickness=3.6e-08 $X=0.159
+ $Y=0.189 $X2=0.229 $Y2=0.189
r162 95 96 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.159 $Y=0.189 $X2=0.159
+ $Y2=0.189
r163 92 141 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.03 $Y2=0.189
r164 91 95 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.159 $Y2=0.189
r165 91 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.189 $X2=0.033
+ $Y2=0.189
r166 88 89 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.172
r167 87 147 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.189
r168 87 89 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.172
r169 86 88 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.164
r170 84 85 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.145
+ $Y=0.135 $X2=0.148 $Y2=0.135
r171 81 84 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.145 $Y2=0.135
r172 79 86 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r173 79 85 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.148 $Y2=0.135
r174 76 77 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r175 74 77 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r176 72 76 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r177 69 70 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r178 67 70 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r179 65 69 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r180 63 64 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r181 62 72 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r182 62 64 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r183 61 137 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.189
r184 61 63 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.2
r185 59 60 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.125
r186 58 137 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.189
r187 58 60 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.125
r188 57 65 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r189 57 59 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r190 55 74 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r191 52 55 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r192 50 67 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r193 47 50 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r194 36 123 39.0385 $w=2.6e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.178 $X2=0.513 $Y2=0.178
r195 28 43 3.07692 $w=2.6e-08 $l=4e-09 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.178 $X2=0.725 $Y2=0.178
r196 28 31 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.178 $X2=0.729 $Y2=0.2295
r197 25 43 82.8571 $w=2.6e-08 $l=1.04e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.725 $Y2=0.178
r198 25 123 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.513 $Y2=0.178
r199 22 25 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0405 $X2=0.621 $Y2=0.178
r200 19 36 3.84615 $w=2.6e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.178 $X2=0.464 $Y2=0.178
r201 16 19 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.178
r202 10 111 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135
+ $X2=0.351 $Y2=0.135
r203 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r204 5 81 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r205 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r206 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%D 2 5 7 12 14 17 VSS
c21 17 VSS 2.32756e-19 $X=0.297 $Y=0.126
c22 14 VSS 0.0072156f $X=0.297 $Y=0.135
c23 12 VSS 0.00703905f $X=0.298 $Y=0.082
c24 5 VSS 0.00200686f $X=0.297 $Y=0.135
c25 2 VSS 0.061556f $X=0.297 $Y=0.0675
r26 16 17 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.126
r27 14 17 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.126
r28 12 16 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.082 $X2=0.297 $Y2=0.106
r29 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r30 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r31 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%6 2 5 7 10 13 15 17 22 25 27 32 34 39 40 42 45
+ 51 53 54 58 63 73 74 76 VSS
c70 76 VSS 7.89434e-19 $X=0.243 $Y=0.2115
c71 74 VSS 9.16337e-19 $X=0.243 $Y=0.126
c72 73 VSS 0.00233088f $X=0.243 $Y=0.106
c73 63 VSS 0.00103743f $X=0.675 $Y=0.135
c74 58 VSS 9.14968e-19 $X=0.405 $Y=0.135
c75 54 VSS 0.00260015f $X=0.601 $Y=0.153
c76 53 VSS 0.00786313f $X=0.527 $Y=0.153
c77 51 VSS 0.00404346f $X=0.675 $Y=0.153
c78 45 VSS 0.00167753f $X=0.243 $Y=0.153
c79 42 VSS 5.5218e-19 $X=0.243 $Y=0.225
c80 40 VSS 0.00181981f $X=0.216 $Y=0.234
c81 39 VSS 0.00525711f $X=0.198 $Y=0.234
c82 34 VSS 0.00482554f $X=0.234 $Y=0.234
c83 33 VSS 0.00200074f $X=0.216 $Y=0.036
c84 32 VSS 0.00545403f $X=0.198 $Y=0.036
c85 27 VSS 0.00500597f $X=0.234 $Y=0.036
c86 25 VSS 0.00648533f $X=0.16 $Y=0.216
c87 20 VSS 0.00602272f $X=0.16 $Y=0.054
c88 13 VSS 0.0021498f $X=0.675 $Y=0.135
c89 10 VSS 0.0585656f $X=0.675 $Y=0.0405
c90 5 VSS 0.00163668f $X=0.405 $Y=0.135
c91 2 VSS 0.058827f $X=0.405 $Y=0.0675
r92 75 76 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.198 $X2=0.243 $Y2=0.2115
r93 73 74 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.106 $X2=0.243 $Y2=0.126
r94 53 54 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.601 $Y2=0.153
r95 51 54 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.675
+ $Y=0.153 $X2=0.601 $Y2=0.153
r96 51 63 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.675 $Y=0.153 $X2=0.675
+ $Y2=0.153
r97 48 53 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.527 $Y2=0.153
r98 48 58 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r99 45 75 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.198
r100 45 74 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.126
r101 44 48 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.405 $Y2=0.153
r102 44 45 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.153 $X2=0.243
+ $Y2=0.153
r103 42 76 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.2115
r104 41 73 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.106
r105 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.216 $Y2=0.234
r106 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.198 $Y2=0.234
r107 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r108 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r109 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.216 $Y2=0.036
r110 29 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r111 27 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r112 27 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r113 25 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r114 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r115 20 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r116 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r117 13 63 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.135 $X2=0.675
+ $Y2=0.135
r118 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2295
r119 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.135
r120 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r121 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2295
r122 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%7 2 5 7 9 10 13 14 17 19 22 29 30 31 33 40 47 48
+ 49 50 51 52 54 55 VSS
c45 56 VSS 3.57489e-19 $X=0.612 $Y=0.09
c46 55 VSS 1.84136e-19 $X=0.603 $Y=0.09
c47 54 VSS 5.96246e-19 $X=0.621 $Y=0.09
c48 52 VSS 4.34894e-19 $X=0.621 $Y=0.214
c49 51 VSS 4.90038e-19 $X=0.621 $Y=0.203
c50 50 VSS 1.59683e-19 $X=0.621 $Y=0.167
c51 49 VSS 2.90654e-19 $X=0.621 $Y=0.165
c52 48 VSS 3.07094e-19 $X=0.621 $Y=0.14
c53 47 VSS 3.66508e-19 $X=0.621 $Y=0.122
c54 46 VSS 3.22511e-19 $X=0.621 $Y=0.225
c55 40 VSS 0.00154565f $X=0.594 $Y=0.054
c56 33 VSS 0.00268134f $X=0.594 $Y=0.234
c57 31 VSS 0.00427376f $X=0.612 $Y=0.234
c58 30 VSS 1.96699e-19 $X=0.583 $Y=0.09
c59 29 VSS 0.00266746f $X=0.581 $Y=0.09
c60 24 VSS 5.17345e-20 $X=0.585 $Y=0.09
c61 22 VSS 0.0179398f $X=0.65 $Y=0.2295
c62 19 VSS 3.14771e-19 $X=0.665 $Y=0.2295
c63 17 VSS 2.5391e-19 $X=0.592 $Y=0.2295
c64 13 VSS 0.0281519f $X=0.594 $Y=0.0405
c65 9 VSS 6.29543e-19 $X=0.611 $Y=0.0405
c66 5 VSS 0.00233073f $X=0.513 $Y=0.09
c67 2 VSS 0.0584396f $X=0.513 $Y=0.0405
r68 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.603
+ $Y=0.09 $X2=0.612 $Y2=0.09
r69 54 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.612 $Y2=0.09
r70 53 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.09 $X2=0.603 $Y2=0.09
r71 51 52 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.214
r72 50 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.203
r73 49 50 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.167
r74 48 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r75 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r76 46 52 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.214
r77 45 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.09
r78 45 47 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.122
r79 38 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.09
r80 38 40 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.054
r81 31 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r82 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r83 29 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.581
+ $Y=0.09 $X2=0.583 $Y2=0.09
r84 26 29 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.09 $X2=0.581 $Y2=0.09
r85 24 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.594 $Y2=0.09
r86 24 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.583 $Y2=0.09
r87 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2295 $X2=0.65 $Y2=0.2295
r88 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.592
+ $Y=0.2295 $X2=0.65 $Y2=0.2295
r89 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r90 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r91 13 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.054 $X2=0.594
+ $Y2=0.054
r92 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.594 $Y2=0.0405
r93 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0405 $X2=0.594 $Y2=0.0405
r94 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.09 $X2=0.513
+ $Y2=0.09
r95 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.09 $X2=0.513 $Y2=0.2295
r96 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.09
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%8 2 5 7 9 14 17 21 22 25 30 31 33 35 36 37 38 39
+ 41 42 43 44 48 50 51 52 53 58 60 61 VSS
c55 64 VSS 2.84134e-19 $X=0.459 $Y=0.131
c56 61 VSS 0.00334468f $X=0.45 $Y=0.036
c57 60 VSS 0.00243127f $X=0.459 $Y=0.036
c58 58 VSS 0.00276391f $X=0.432 $Y=0.036
c59 53 VSS 4.23521e-19 $X=0.5445 $Y=0.131
c60 52 VSS 3.49205e-20 $X=0.522 $Y=0.131
c61 51 VSS 2.00095e-19 $X=0.504 $Y=0.131
c62 50 VSS 0.00133241f $X=0.496 $Y=0.131
c63 48 VSS 5.65734e-19 $X=0.567 $Y=0.131
c64 45 VSS 4.53296e-19 $X=0.459 $Y=0.214
c65 44 VSS 2.01779e-19 $X=0.459 $Y=0.203
c66 43 VSS 6.09344e-21 $X=0.459 $Y=0.167
c67 42 VSS 1.60693e-19 $X=0.459 $Y=0.165
c68 41 VSS 3.22878e-19 $X=0.459 $Y=0.225
c69 39 VSS 2.48018e-19 $X=0.459 $Y=0.114
c70 38 VSS 2.26591e-19 $X=0.459 $Y=0.106
c71 37 VSS 9.45429e-20 $X=0.459 $Y=0.099
c72 36 VSS 8.12259e-19 $X=0.459 $Y=0.081
c73 35 VSS 2.08428e-19 $X=0.459 $Y=0.122
c74 33 VSS 0.00142907f $X=0.434 $Y=0.234
c75 32 VSS 3.66528e-19 $X=0.418 $Y=0.234
c76 31 VSS 0.00146362f $X=0.414 $Y=0.234
c77 30 VSS 0.00368178f $X=0.396 $Y=0.234
c78 25 VSS 0.00389542f $X=0.45 $Y=0.234
c79 24 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c80 21 VSS 0.00348256f $X=0.378 $Y=0.2025
c81 16 VSS 5.70081e-19 $X=0.432 $Y=0.0405
c82 5 VSS 0.00195718f $X=0.567 $Y=0.1305
c83 2 VSS 0.0591962f $X=0.567 $Y=0.0405
r84 61 62 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r85 60 62 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r86 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r87 57 58 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r88 52 53 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r89 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r90 50 51 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.496
+ $Y=0.131 $X2=0.504 $Y2=0.131
r91 48 53 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r92 46 64 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r93 46 50 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.496 $Y2=0.131
r94 44 45 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.203 $X2=0.459 $Y2=0.214
r95 43 44 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.167 $X2=0.459 $Y2=0.203
r96 42 43 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.167
r97 41 45 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r98 40 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r99 40 42 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.165
r100 38 39 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.106 $X2=0.459 $Y2=0.114
r101 37 38 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.099 $X2=0.459 $Y2=0.106
r102 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.099
r103 35 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r104 35 39 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.114
r105 34 60 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r106 34 36 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.081
r107 32 33 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.234 $X2=0.434 $Y2=0.234
r108 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.418 $Y2=0.234
r109 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r110 27 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r111 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r112 25 33 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.434 $Y2=0.234
r113 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r114 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r115 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r116 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r117 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r118 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r119 13 58 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r120 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r121 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r122 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r123 5 48 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.131 $X2=0.567
+ $Y2=0.131
r124 5 7 370.904 $w=2e-08 $l=9.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1305 $X2=0.567 $Y2=0.2295
r125 2 5 337.185 $w=2e-08 $l=9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.1305
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%9 2 5 7 9 14 21 25 26 30 31 32 33 34 39 40 42 44
+ 45 VSS
c24 46 VSS 1.99706e-19 $X=0.945 $Y=0.171
c25 45 VSS 0.00100047f $X=0.945 $Y=0.167
c26 44 VSS 8.83619e-19 $X=0.945 $Y=0.117
c27 43 VSS 0.00226287f $X=0.945 $Y=0.09
c28 42 VSS 0.00286673f $X=0.945 $Y=0.225
c29 40 VSS 0.0018377f $X=0.918 $Y=0.234
c30 39 VSS 0.0056872f $X=0.9 $Y=0.234
c31 34 VSS 0.00462933f $X=0.936 $Y=0.234
c32 33 VSS 0.00189638f $X=0.9 $Y=0.036
c33 32 VSS 0.00352438f $X=0.882 $Y=0.036
c34 31 VSS 0.00146362f $X=0.846 $Y=0.036
c35 30 VSS 0.00508235f $X=0.828 $Y=0.036
c36 26 VSS 0.00226308f $X=0.792 $Y=0.036
c37 25 VSS 0.00657446f $X=0.936 $Y=0.036
c38 21 VSS 0.00122443f $X=0.783 $Y=0.105
c39 17 VSS 0.0048151f $X=0.862 $Y=0.2295
c40 12 VSS 0.00513464f $X=0.862 $Y=0.0405
c41 5 VSS 0.00277722f $X=0.783 $Y=0.1055
c42 2 VSS 0.0590816f $X=0.783 $Y=0.0405
r43 45 46 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.167 $X2=0.945 $Y2=0.171
r44 44 45 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.117 $X2=0.945 $Y2=0.167
r45 43 44 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.09 $X2=0.945 $Y2=0.117
r46 42 46 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.171
r47 41 43 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.09
r48 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.234 $X2=0.918 $Y2=0.234
r49 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.9 $Y2=0.234
r50 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r51 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.918 $Y2=0.234
r52 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r53 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.846 $Y2=0.036
r54 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r55 28 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.846 $Y2=0.036
r56 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.036 $X2=0.828 $Y2=0.036
r57 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r58 25 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.9 $Y2=0.036
r59 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.783 $Y=0.045 $X2=0.792 $Y2=0.036
r60 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.105
r61 17 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234 $X2=0.864
+ $Y2=0.234
r62 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2295 $X2=0.862 $Y2=0.2295
r63 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036 $X2=0.864
+ $Y2=0.036
r64 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.862 $Y2=0.0405
r65 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.105 $X2=0.783
+ $Y2=0.105
r66 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.1055 $X2=0.783 $Y2=0.2295
r67 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.1055
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%10 2 7 10 15 18 21 23 25 26 29 30 31 34 35 40 41
+ 43 45 46 47 48 49 51 52 54 55 58 65 66 74 77 81 84 92 VSS
c67 92 VSS 0.00216926f $X=0.999 $Y=0.135
c68 84 VSS 0.00793307f $X=0.999 $Y=0.153
c69 81 VSS 0.00150008f $X=0.891 $Y=0.153
c70 78 VSS 4.17512e-19 $X=0.837 $Y=0.162
c71 77 VSS 1.52743e-19 $X=0.729 $Y=0.162
c72 74 VSS 0.00370746f $X=0.72 $Y=0.234
c73 73 VSS 0.00266816f $X=0.729 $Y=0.234
c74 66 VSS 4.30636e-19 $X=0.866 $Y=0.162
c75 65 VSS 1.48695e-19 $X=0.85 $Y=0.162
c76 63 VSS 2.75449e-19 $X=0.882 $Y=0.162
c77 58 VSS 3.94906e-19 $X=0.837 $Y=0.135
c78 55 VSS 3.26354e-19 $X=0.792 $Y=0.162
c79 54 VSS 0.00206921f $X=0.774 $Y=0.162
c80 52 VSS 0.00192346f $X=0.828 $Y=0.162
c81 51 VSS 0.00136716f $X=0.729 $Y=0.225
c82 49 VSS 1.52884e-19 $X=0.729 $Y=0.136
c83 48 VSS 9.59255e-20 $X=0.729 $Y=0.119
c84 47 VSS 1.29374e-19 $X=0.729 $Y=0.099
c85 46 VSS 3.52175e-19 $X=0.729 $Y=0.081
c86 45 VSS 2.74133e-19 $X=0.729 $Y=0.153
c87 43 VSS 0.00166816f $X=0.704 $Y=0.036
c88 42 VSS 4.57836e-19 $X=0.688 $Y=0.036
c89 41 VSS 0.00146362f $X=0.684 $Y=0.036
c90 40 VSS 0.00370471f $X=0.666 $Y=0.036
c91 35 VSS 0.00409787f $X=0.72 $Y=0.036
c92 34 VSS 0.00276615f $X=0.702 $Y=0.2295
c93 30 VSS 5.63046e-19 $X=0.719 $Y=0.2295
c94 29 VSS 0.0349304f $X=0.648 $Y=0.0405
c95 25 VSS 5.63046e-19 $X=0.665 $Y=0.0405
c96 21 VSS 0.00476599f $X=1.053 $Y=0.135
c97 18 VSS 0.0616937f $X=1.053 $Y=0.0675
c98 10 VSS 0.0612321f $X=0.999 $Y=0.0675
c99 5 VSS 0.00189441f $X=0.837 $Y=0.135
c100 2 VSS 0.0618222f $X=0.837 $Y=0.0405
r101 84 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.999 $Y=0.153 $X2=0.999
+ $Y2=0.153
r102 80 84 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.999 $Y2=0.153
r103 80 81 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r104 74 75 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.234 $X2=0.7245 $Y2=0.234
r105 73 75 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.234 $X2=0.7245 $Y2=0.234
r106 70 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.234 $X2=0.72 $Y2=0.234
r107 65 66 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.85
+ $Y=0.162 $X2=0.866 $Y2=0.162
r108 64 78 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.837 $Y2=0.162
r109 64 65 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.85 $Y2=0.162
r110 63 81 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.891 $Y2=0.162
r111 63 66 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.866 $Y2=0.162
r112 56 78 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.162
r113 56 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.135
r114 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.162 $X2=0.792 $Y2=0.162
r115 53 77 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.729 $Y2=0.162
r116 53 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.774 $Y2=0.162
r117 52 78 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.837 $Y2=0.162
r118 52 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.792 $Y2=0.162
r119 51 73 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.225 $X2=0.729 $Y2=0.234
r120 50 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.162
r121 50 51 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.225
r122 48 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.119 $X2=0.729 $Y2=0.136
r123 47 48 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.099 $X2=0.729 $Y2=0.119
r124 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.081 $X2=0.729 $Y2=0.099
r125 45 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.162
r126 45 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.136
r127 44 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.045 $X2=0.729 $Y2=0.081
r128 42 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.036 $X2=0.704 $Y2=0.036
r129 41 42 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.688 $Y2=0.036
r130 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.684 $Y2=0.036
r131 37 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.666 $Y2=0.036
r132 35 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.036 $X2=0.729 $Y2=0.045
r133 35 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.704 $Y2=0.036
r134 34 70 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.234
+ $X2=0.702 $Y2=0.234
r135 31 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2295 $X2=0.702 $Y2=0.2295
r136 30 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2295 $X2=0.702 $Y2=0.2295
r137 29 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r138 26 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0405 $X2=0.648 $Y2=0.0405
r139 25 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r140 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.135 $X2=1.053 $Y2=0.2025
r141 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.0675 $X2=1.053 $Y2=0.135
r142 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.999
+ $Y=0.135 $X2=1.053 $Y2=0.135
r143 13 92 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.135 $X2=0.999
+ $Y2=0.135
r144 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.135 $X2=0.999 $Y2=0.2025
r145 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.135
r146 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.135 $X2=0.837
+ $Y2=0.135
r147 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.2295
r148 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.0405 $X2=0.837 $Y2=0.135
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%QN 1 2 6 7 10 11 14 16 24 26 VSS
c13 28 VSS 0.00180641f $X=1.106 $Y=0.196
c14 26 VSS 0.00147086f $X=1.106 $Y=0.1155
c15 25 VSS 0.00247539f $X=1.106 $Y=0.09
c16 24 VSS 0.00279276f $X=1.103 $Y=0.141
c17 22 VSS 0.00150428f $X=1.106 $Y=0.225
c18 16 VSS 0.014442f $X=1.097 $Y=0.234
c19 14 VSS 0.00966022f $X=1.026 $Y=0.036
c20 11 VSS 0.014442f $X=1.097 $Y=0.036
c21 10 VSS 0.00941949f $X=1.026 $Y=0.2025
c22 6 VSS 5.72268e-19 $X=1.043 $Y=0.2025
c23 1 VSS 5.72268e-19 $X=1.043 $Y=0.0675
r24 27 28 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.106
+ $Y=0.167 $X2=1.106 $Y2=0.196
r25 25 26 1.73148 $w=1.8e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=1.106
+ $Y=0.09 $X2=1.106 $Y2=0.1155
r26 24 27 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.106
+ $Y=0.141 $X2=1.106 $Y2=0.167
r27 24 26 1.73148 $w=1.8e-08 $l=2.55e-08 $layer=M1 $thickness=3.6e-08 $X=1.106
+ $Y=0.141 $X2=1.106 $Y2=0.1155
r28 22 28 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.106
+ $Y=0.225 $X2=1.106 $Y2=0.196
r29 21 25 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.106
+ $Y=0.045 $X2=1.106 $Y2=0.09
r30 16 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.097 $Y=0.234 $X2=1.106 $Y2=0.225
r31 16 18 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.097
+ $Y=0.234 $X2=1.026 $Y2=0.234
r32 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.036 $X2=1.026
+ $Y2=0.036
r33 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.097 $Y=0.036 $X2=1.106 $Y2=0.045
r34 11 13 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.097
+ $Y=0.036 $X2=1.026 $Y2=0.036
r35 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.234 $X2=1.026
+ $Y2=0.234
r36 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.2025 $X2=1.026 $Y2=0.2025
r37 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.043 $Y=0.2025 $X2=1.026 $Y2=0.2025
r38 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.026
+ $Y=0.0675 $X2=1.026 $Y2=0.036
r39 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.009
+ $Y=0.0675 $X2=1.026 $Y2=0.0675
r40 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.043
+ $Y=0.0675 $X2=1.026 $Y2=0.0675
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%12 1 6 9 VSS
c6 9 VSS 0.0266112f $X=0.38 $Y=0.0675
c7 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c8 4 VSS 3.22674e-19 $X=0.322 $Y=0.0675
r9 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r10 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%13 1 6 9 VSS
c10 9 VSS 0.0209308f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.69239e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%14 1 6 9 VSS
c8 9 VSS 0.0191793f $X=0.758 $Y=0.0405
c9 6 VSS 3.14771e-19 $X=0.773 $Y=0.0405
c10 4 VSS 2.61968e-19 $X=0.7 $Y=0.0405
r11 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r12 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.7
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r13 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.685
+ $Y=0.0405 $X2=0.7 $Y2=0.0405
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%15 1 2 VSS
c0 1 VSS 0.00225696f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%16 1 2 VSS
c1 1 VSS 0.00201018f $X=0.341 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends

.subckt PM_DFFLQNX2_ASAP7_75T_SRAM%17 1 2 VSS
c0 1 VSS 0.00219822f $X=0.773 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2295 $X2=0.739 $Y2=0.2295
.ends


* END of "./DFFLQNx2_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DFFLQNx2_ASAP7_75t_SRAM  VSS VDD CLK D QN
* 
* QN	QN
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_12_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_6_M3_g N_12_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_15_M4_d N_4_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_15_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_10_M7_d N_4_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.611
+ $Y=0.027
M8 N_14_M8_d N_6_M8_g N_10_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M9 VSS N_9_M9_g N_14_M9_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_9_M10_d N_10_M10_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.027
M11 N_QN_M11_d N_10_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M12 N_QN_M12_d N_10_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.027
M13 VDD N_CLK_M13_g N_4_M13_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M14 N_6_M14_d N_4_M14_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M15 N_16_M15_d N_D_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M16 N_8_M16_d N_4_M16_g N_16_M16_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M17 N_13_M17_d N_6_M17_g N_8_M17_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M18 VDD N_7_M18_g N_13_M18_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M19 N_7_M19_d N_8_M19_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M20 N_10_M20_d N_6_M20_g N_7_M20_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.665 $Y=0.216
M21 N_17_M21_d N_4_M21_g N_10_M21_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.719 $Y=0.216
M22 VDD N_9_M22_g N_17_M22_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M23 N_9_M23_d N_10_M23_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.216
M24 N_QN_M24_d N_10_M24_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
M25 N_QN_M25_d N_10_M25_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.162
*
* 
* .include "DFFLQNx2_ASAP7_75t_SRAM.pex.sp.DFFLQNX2_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DFFLQNx2_ASAP7_75t_SRAM.pex.sp.DFFLQNX2_ASAP7_75T_SRAM.pxi"
* File: DFFLQNx2_ASAP7_75t_SRAM.pex.sp.DFFLQNX2_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:26:01 2017
* 
x_PM_DFFLQNX2_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M13_g CLK N_CLK_c_4_p
+ N_CLK_c_10_p VSS PM_DFFLQNX2_ASAP7_75T_SRAM%CLK
x_PM_DFFLQNX2_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_20_n N_4_M14_g N_4_c_34_p N_4_M16_g
+ N_4_M4_g N_4_M7_g N_4_c_77_p N_4_c_43_p N_4_M21_g N_4_c_89_p N_4_c_44_p
+ N_4_M0_s N_4_c_21_n N_4_M13_s N_4_c_22_n N_4_c_23_n N_4_c_24_n N_4_c_25_n
+ N_4_c_26_n N_4_c_27_n N_4_c_47_p N_4_c_28_n N_4_c_29_n N_4_c_30_n N_4_c_31_n
+ N_4_c_32_n N_4_c_58_p N_4_c_33_n N_4_c_36_p N_4_c_37_p N_4_c_38_p N_4_c_61_p
+ N_4_c_94_p N_4_c_46_p VSS PM_DFFLQNX2_ASAP7_75T_SRAM%4
x_PM_DFFLQNX2_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_122_n N_D_M15_g D N_D_c_123_n
+ N_D_c_133_p VSS PM_DFFLQNX2_ASAP7_75T_SRAM%D
x_PM_DFFLQNX2_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_147_n N_6_M17_g N_6_M8_g N_6_c_151_n
+ N_6_M20_g N_6_M1_d N_6_M14_d N_6_c_152_n N_6_c_172_n N_6_c_142_n N_6_c_154_n
+ N_6_c_143_n N_6_c_158_n N_6_c_174_n N_6_c_159_n N_6_c_161_n N_6_c_162_n
+ N_6_c_183_p N_6_c_168_n N_6_c_170_n N_6_c_144_n N_6_c_180_n N_6_c_181_n VSS
+ PM_DFFLQNX2_ASAP7_75T_SRAM%6
x_PM_DFFLQNX2_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_237_p N_7_M18_g N_7_M7_s N_7_M6_d
+ N_7_c_216_n N_7_M19_d N_7_c_217_n N_7_M20_s N_7_c_219_n N_7_c_235_p
+ N_7_c_228_n N_7_c_255_p N_7_c_229_n N_7_c_236_p N_7_c_221_n N_7_c_240_p
+ N_7_c_222_n N_7_c_223_n N_7_c_224_n N_7_c_253_p N_7_c_226_n N_7_c_233_n VSS
+ PM_DFFLQNX2_ASAP7_75T_SRAM%7
x_PM_DFFLQNX2_ASAP7_75T_SRAM%8 N_8_M6_g N_8_c_280_n N_8_M19_g N_8_M3_d N_8_M4_s
+ N_8_M16_d N_8_c_260_n N_8_M17_s N_8_c_308_p N_8_c_262_n N_8_c_283_n
+ N_8_c_309_p N_8_c_285_n N_8_c_263_n N_8_c_264_n N_8_c_298_n N_8_c_286_n
+ N_8_c_310_p N_8_c_265_n N_8_c_266_n N_8_c_268_n N_8_c_299_n N_8_c_272_n
+ N_8_c_300_n N_8_c_273_n N_8_c_275_n N_8_c_291_n N_8_c_303_n N_8_c_278_n VSS
+ PM_DFFLQNX2_ASAP7_75T_SRAM%8
x_PM_DFFLQNX2_ASAP7_75T_SRAM%9 N_9_M9_g N_9_c_318_p N_9_M22_g N_9_M10_d N_9_M23_d
+ N_9_c_317_p N_9_c_329_p N_9_c_316_p N_9_c_321_p N_9_c_315_p N_9_c_325_p
+ N_9_c_327_p N_9_c_334_p N_9_c_326_p N_9_c_330_p N_9_c_320_p N_9_c_332_p
+ N_9_c_328_p VSS PM_DFFLQNX2_ASAP7_75T_SRAM%9
x_PM_DFFLQNX2_ASAP7_75T_SRAM%10 N_10_M10_g N_10_M23_g N_10_M11_g N_10_M24_g
+ N_10_M12_g N_10_c_387_p N_10_M25_g N_10_M8_s N_10_M7_d N_10_c_337_n N_10_M21_s
+ N_10_M20_d N_10_c_339_n N_10_c_370_n N_10_c_350_n N_10_c_351_n N_10_c_400_p
+ N_10_c_353_n N_10_c_362_n N_10_c_340_n N_10_c_341_n N_10_c_342_n N_10_c_343_n
+ N_10_c_375_n N_10_c_345_n N_10_c_376_n N_10_c_378_n N_10_c_379_n N_10_c_380_n
+ N_10_c_346_n N_10_c_347_n N_10_c_381_n N_10_c_355_n N_10_c_386_n VSS
+ PM_DFFLQNX2_ASAP7_75T_SRAM%10
x_PM_DFFLQNX2_ASAP7_75T_SRAM%QN N_QN_M12_d N_QN_M11_d N_QN_M25_d N_QN_M24_d
+ N_QN_c_407_n N_QN_c_403_n N_QN_c_410_n N_QN_c_404_n QN N_QN_c_415_n VSS
+ PM_DFFLQNX2_ASAP7_75T_SRAM%QN
x_PM_DFFLQNX2_ASAP7_75T_SRAM%12 N_12_M2_d N_12_M3_s N_12_c_416_n VSS
+ PM_DFFLQNX2_ASAP7_75T_SRAM%12
x_PM_DFFLQNX2_ASAP7_75T_SRAM%13 N_13_M17_d N_13_M18_s N_13_c_423_n VSS
+ PM_DFFLQNX2_ASAP7_75T_SRAM%13
x_PM_DFFLQNX2_ASAP7_75T_SRAM%14 N_14_M8_d N_14_M9_s N_14_c_432_n VSS
+ PM_DFFLQNX2_ASAP7_75T_SRAM%14
x_PM_DFFLQNX2_ASAP7_75T_SRAM%15 N_15_M5_s N_15_M4_d VSS PM_DFFLQNX2_ASAP7_75T_SRAM%15
x_PM_DFFLQNX2_ASAP7_75T_SRAM%16 N_16_M16_s N_16_M15_d VSS
+ PM_DFFLQNX2_ASAP7_75T_SRAM%16
x_PM_DFFLQNX2_ASAP7_75T_SRAM%17 N_17_M22_s N_17_M21_d VSS
+ PM_DFFLQNX2_ASAP7_75T_SRAM%17
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_CLK_c_2_p N_4_c_20_n 0.00124017f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 CLK N_4_c_21_n 3.57152e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_4 N_CLK_c_4_p N_4_c_22_n 0.00206543f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.18
cc_5 CLK N_4_c_23_n 2.75361e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.07
cc_6 CLK N_4_c_24_n 0.00206543f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.125
cc_7 N_CLK_c_4_p N_4_c_25_n 2.75361e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2125
cc_8 CLK N_4_c_26_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_4_p N_4_c_27_n 5.03453e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_10_p N_4_c_28_n 8.76278e-19 $X=0.081 $Y=0.1305 $X2=0.145 $Y2=0.135
cc_11 N_CLK_c_4_p N_4_c_29_n 3.53816e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.164
cc_12 N_CLK_c_4_p N_4_c_30_n 6.15177e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.172
cc_13 N_CLK_c_4_p N_4_c_31_n 0.00138527f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.189
cc_14 N_CLK_c_4_p N_4_c_32_n 9.65218e-19 $X=0.081 $Y=0.135 $X2=0.159 $Y2=0.189
cc_15 N_CLK_c_4_p N_4_c_33_n 0.00167589f $X=0.081 $Y=0.135 $X2=0.229 $Y2=0.189
cc_16 CLK N_6_c_142_n 6.45949e-19 $X=0.082 $Y=0.119 $X2=0 $Y2=0
cc_17 N_CLK_c_4_p N_6_c_143_n 6.54444e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_18 CLK N_6_c_144_n 6.20748e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.234
cc_19 N_4_c_34_p N_D_M2_g 0.00341068f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.054
cc_20 N_4_c_34_p N_D_c_122_n 0.0010364f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 N_4_c_36_p N_D_c_123_n 2.29805e-19 $X=0.29 $Y=0.189 $X2=0.081 $Y2=0.135
cc_22 N_4_c_37_p N_D_c_123_n 0.00102387f $X=0.513 $Y=0.189 $X2=0.081 $Y2=0.135
cc_23 N_4_c_38_p N_D_c_123_n 0.00337064f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_4_c_34_p N_6_M3_g 0.00355599f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.054
cc_25 N_4_M4_g N_6_M3_g 0.00355599f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_26 N_4_c_34_p N_6_c_147_n 0.00103664f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_27 N_4_M7_g N_6_M8_g 0.00355599f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_28 N_4_c_43_p N_6_M8_g 0.00355599f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_29 N_4_c_44_p N_6_M8_g 0.00250257f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_30 N_4_c_44_p N_6_c_151_n 0.00180656f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_31 N_4_c_46_p N_6_c_152_n 0.00135022f $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_32 N_4_c_47_p N_6_c_142_n 0.0010851f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_33 N_4_c_36_p N_6_c_154_n 4.24027e-19 $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_34 N_4_c_32_n N_6_c_143_n 0.00285029f $X=0.159 $Y=0.189 $X2=0 $Y2=0
cc_35 N_4_c_33_n N_6_c_143_n 6.46981e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_36 N_4_c_46_p N_6_c_143_n 2.904e-19 $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_37 N_4_c_33_n N_6_c_158_n 4.24027e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_38 N_4_c_47_p N_6_c_159_n 0.00351854f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_39 N_4_c_36_p N_6_c_159_n 0.00102595f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_40 N_4_c_44_p N_6_c_161_n 6.40799e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_41 N_4_c_44_p N_6_c_162_n 0.00187197f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_42 N_4_c_29_n N_6_c_162_n 3.52457e-19 $X=0.189 $Y=0.164 $X2=0 $Y2=0
cc_43 N_4_c_58_p N_6_c_162_n 2.46239e-19 $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_44 N_4_c_36_p N_6_c_162_n 0.0253778f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_45 N_4_c_38_p N_6_c_162_n 0.00115493f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_61_p N_6_c_162_n 2.81476e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_47 N_4_c_37_p N_6_c_168_n 2.98936e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_48 N_4_c_38_p N_6_c_168_n 0.00170246f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_49 N_4_c_44_p N_6_c_170_n 0.00124003f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_50 N_4_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_51 N_4_M7_g N_7_M5_g 2.13359e-19 $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_52 N_4_c_44_p N_7_M5_g 0.00205997f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_53 N_4_c_61_p N_7_M5_g 3.15189e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_54 N_4_c_44_p N_7_c_216_n 5.49754e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_55 N_4_c_44_p N_7_c_217_n 2.12581e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.1305
cc_56 N_4_c_44_p N_7_M20_s 2.50995e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_57 N_4_M7_g N_7_c_219_n 0.00200065f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_58 N_4_c_44_p N_7_c_219_n 0.00322783f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_59 N_4_M7_g N_7_c_221_n 3.04073e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_60 N_4_M7_g N_7_c_222_n 2.22997e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_61 N_4_c_61_p N_7_c_223_n 5.74745e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_62 N_4_c_77_p N_7_c_224_n 0.00193027f $X=0.621 $Y=0.178 $X2=0 $Y2=0
cc_63 N_4_c_44_p N_7_c_224_n 0.00189849f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_64 N_4_M7_g N_7_c_226_n 3.8308e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_65 N_4_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_66 N_4_M7_g N_8_M6_g 0.00341068f $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_67 N_4_c_44_p N_8_M6_g 0.00302156f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_68 N_4_c_37_p N_8_c_260_n 3.15319e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_69 N_4_c_38_p N_8_c_260_n 0.00136448f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_70 N_4_c_37_p N_8_c_262_n 0.00161272f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_71 N_4_M4_g N_8_c_263_n 3.80535e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_72 N_4_M4_g N_8_c_264_n 2.08362e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_73 N_4_M4_g N_8_c_265_n 2.27303e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_74 N_4_c_89_p N_8_c_266_n 4.73369e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_75 N_4_c_61_p N_8_c_266_n 0.00174159f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_76 N_4_c_89_p N_8_c_268_n 0.0017128f $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_77 N_4_c_44_p N_8_c_268_n 5.88593e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_78 N_4_c_37_p N_8_c_268_n 0.00102123f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_79 N_4_c_94_p N_8_c_268_n 3.42482e-19 $X=0.351 $Y=0.178 $X2=0 $Y2=0
cc_80 N_4_c_44_p N_8_c_272_n 8.16411e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_81 N_4_c_44_p N_8_c_273_n 3.32592e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_82 N_4_c_61_p N_8_c_273_n 8.9822e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_83 N_4_c_44_p N_8_c_275_n 5.02733e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_84 N_4_c_43_p N_9_M9_g 0.00341068f $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_85 N_4_c_43_p N_10_M10_g 2.13359e-19 $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_86 N_4_c_44_p N_10_c_337_n 8.27829e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_87 N_4_c_44_p N_10_M21_s 3.37661e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_88 N_4_c_44_p N_10_c_339_n 0.00145657f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_89 N_4_c_43_p N_10_c_340_n 2.71526e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_90 N_4_c_43_p N_10_c_341_n 2.11119e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_91 N_4_c_43_p N_10_c_342_n 2.58771e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_92 N_4_c_43_p N_10_c_343_n 0.00229157f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_93 N_4_c_44_p N_10_c_343_n 7.89371e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_94 N_4_c_43_p N_10_c_345_n 4.55487e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_95 N_4_c_44_p N_10_c_346_n 4.45535e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_96 N_4_c_43_p N_10_c_347_n 5.68093e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_97 N_4_c_44_p N_10_c_347_n 2.2968e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_98 N_4_c_34_p N_12_c_416_n 0.00526068f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_99 N_4_c_44_p N_13_M18_s 2.36286e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.216
cc_100 N_4_M4_g N_13_c_423_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_101 N_4_c_89_p N_13_c_423_n 5.41258e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_102 N_4_c_44_p N_13_c_423_n 0.00230928f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_103 N_4_c_37_p N_13_c_423_n 7.09553e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_104 N_4_c_43_p N_14_c_432_n 0.00198387f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_105 N_4_c_44_p N_14_c_432_n 4.51352e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_106 N_D_M2_g N_6_M3_g 2.82885e-19 $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_107 D N_6_c_172_n 0.00115224f $X=0.298 $Y=0.082 $X2=0.729 $Y2=0.178
cc_108 N_D_c_123_n N_6_c_154_n 0.00115224f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_109 N_D_c_123_n N_6_c_174_n 0.00115224f $X=0.297 $Y=0.135 $X2=0.725 $Y2=0.178
cc_110 N_D_c_123_n N_6_c_159_n 0.00124565f $X=0.297 $Y=0.135 $X2=0.729 $Y2=0.178
cc_111 D N_6_c_162_n 2.27807e-19 $X=0.298 $Y=0.082 $X2=0.056 $Y2=0.216
cc_112 N_D_c_123_n N_6_c_162_n 9.62099e-19 $X=0.297 $Y=0.135 $X2=0.056 $Y2=0.216
cc_113 N_D_c_133_p N_6_c_168_n 4.3159e-19 $X=0.297 $Y=0.126 $X2=0.018 $Y2=0.18
cc_114 D N_6_c_144_n 0.00115224f $X=0.298 $Y=0.082 $X2=0.054 $Y2=0.234
cc_115 N_D_c_133_p N_6_c_180_n 0.00115224f $X=0.297 $Y=0.126 $X2=0.054 $Y2=0.234
cc_116 N_D_c_123_n N_6_c_181_n 0.00115224f $X=0.297 $Y=0.135 $X2=0.047 $Y2=0.234
cc_117 N_D_c_123_n N_8_c_260_n 3.88702e-19 $X=0.297 $Y=0.135 $X2=0.621
+ $Y2=0.0405
cc_118 N_D_c_123_n N_8_c_262_n 8.77202e-19 $X=0.297 $Y=0.135 $X2=0.729
+ $Y2=0.2295
cc_119 D N_8_c_278_n 2.04306e-19 $X=0.298 $Y=0.082 $X2=0.018 $Y2=0.198
cc_120 D N_12_c_416_n 0.00430488f $X=0.298 $Y=0.082 $X2=0.351 $Y2=0.135
cc_121 N_D_c_123_n N_16_M16_s 3.05674e-19 $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_122 N_6_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_123 N_6_c_183_p N_7_c_228_n 2.96121e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_124 N_6_c_161_n N_7_c_229_n 2.61213e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_125 N_6_c_183_p N_7_c_229_n 2.61213e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_126 N_6_c_170_n N_7_c_221_n 0.00327797f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_127 N_6_c_161_n N_7_c_222_n 0.00115177f $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_128 N_6_c_161_n N_7_c_233_n 2.96121e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_129 N_6_M8_g N_8_M6_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_130 N_6_c_151_n N_8_c_280_n 4.12331e-19 $X=0.675 $Y=0.135 $X2=0.081 $Y2=0.135
cc_131 N_6_c_183_p N_8_c_280_n 2.64012e-19 $X=0.601 $Y=0.153 $X2=0.081 $Y2=0.135
cc_132 N_6_c_168_n N_8_c_260_n 2.25088e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_133 N_6_M3_g N_8_c_283_n 3.49806e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_134 N_6_c_168_n N_8_c_283_n 3.83282e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_135 N_6_c_168_n N_8_c_285_n 9.70699e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_136 N_6_c_168_n N_8_c_286_n 9.70699e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_137 N_6_c_162_n N_8_c_265_n 0.00118282f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_138 N_6_c_168_n N_8_c_265_n 0.00106411f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_139 N_6_c_162_n N_8_c_272_n 0.00138951f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_140 N_6_c_183_p N_8_c_275_n 0.00138951f $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_141 N_6_c_162_n N_8_c_291_n 2.54113e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_142 N_6_c_162_n N_8_c_278_n 3.92135e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_143 N_6_M8_g N_9_M9_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_144 N_6_c_161_n N_10_c_337_n 2.24654e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_145 N_6_c_161_n N_10_c_350_n 5.06919e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_146 N_6_M8_g N_10_c_351_n 3.43727e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_147 N_6_c_170_n N_10_c_351_n 5.96743e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_148 N_6_c_161_n N_10_c_353_n 2.34004e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_149 N_6_c_170_n N_10_c_341_n 0.00329725f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_150 N_6_c_161_n N_10_c_355_n 2.83245e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_151 N_6_c_162_n N_12_c_416_n 8.35084e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_152 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_153 N_7_c_235_p N_8_M6_g 3.91159e-19 $X=0.581 $Y=0.09 $X2=0.135 $Y2=0.054
cc_154 N_7_c_236_p N_8_c_263_n 2.10569e-19 $X=0.594 $Y=0.054 $X2=0.464 $Y2=0.178
cc_155 N_7_c_237_p N_8_c_264_n 3.19692e-19 $X=0.513 $Y=0.09 $X2=0 $Y2=0
cc_156 N_7_c_235_p N_8_c_264_n 0.00107929f $X=0.581 $Y=0.09 $X2=0 $Y2=0
cc_157 N_7_c_221_n N_8_c_298_n 2.4251e-19 $X=0.621 $Y=0.122 $X2=0 $Y2=0
cc_158 N_7_c_240_p N_8_c_299_n 9.84729e-19 $X=0.621 $Y=0.14 $X2=0.056 $Y2=0.054
cc_159 N_7_c_235_p N_8_c_300_n 0.00507595f $X=0.581 $Y=0.09 $X2=0 $Y2=0
cc_160 N_7_M5_g N_8_c_273_n 3.12986e-19 $X=0.513 $Y=0.0405 $X2=0.071 $Y2=0.216
cc_161 N_7_c_237_p N_8_c_291_n 5.2508e-19 $X=0.513 $Y=0.09 $X2=0.018 $Y2=0.18
cc_162 N_7_c_236_p N_8_c_303_n 2.10569e-19 $X=0.594 $Y=0.054 $X2=0.018 $Y2=0.125
cc_163 N_7_c_216_n N_10_c_337_n 0.00328169f $X=0.594 $Y=0.0405 $X2=0 $Y2=0
cc_164 N_7_c_236_p N_10_c_337_n 3.00222e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_165 N_7_c_226_n N_10_c_337_n 2.70684e-19 $X=0.621 $Y=0.09 $X2=0 $Y2=0
cc_166 N_7_c_219_n N_10_c_339_n 0.00222825f $X=0.65 $Y=0.2295 $X2=0 $Y2=0
cc_167 N_7_c_216_n N_10_c_350_n 3.50513e-19 $X=0.594 $Y=0.0405 $X2=0 $Y2=0
cc_168 N_7_c_236_p N_10_c_350_n 5.0339e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_169 N_7_c_236_p N_10_c_362_n 2.21141e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_170 N_7_c_226_n N_10_c_340_n 4.36168e-19 $X=0.621 $Y=0.09 $X2=0.071 $Y2=0.054
cc_171 N_7_c_253_p N_10_c_343_n 4.36168e-19 $X=0.621 $Y=0.214 $X2=0 $Y2=0
cc_172 N_7_c_219_n N_10_c_346_n 3.64454e-19 $X=0.65 $Y=0.2295 $X2=0.054
+ $Y2=0.234
cc_173 N_7_c_255_p N_10_c_346_n 4.86017e-19 $X=0.612 $Y=0.234 $X2=0.054
+ $Y2=0.234
cc_174 N_7_c_224_n N_10_c_347_n 4.36168e-19 $X=0.621 $Y=0.203 $X2=0.0505
+ $Y2=0.234
cc_175 N_8_c_260_n N_12_c_416_n 0.00119636f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.135
cc_176 N_8_c_291_n N_12_c_416_n 0.00390673f $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_177 N_8_c_278_n N_12_c_416_n 4.41747e-19 $X=0.45 $Y=0.036 $X2=0.351 $Y2=0.135
cc_178 N_8_c_260_n N_13_c_423_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.135
cc_179 N_8_c_308_p N_13_c_423_n 0.00209454f $X=0.45 $Y=0.234 $X2=0.351 $Y2=0.135
cc_180 N_8_c_309_p N_13_c_423_n 0.0013184f $X=0.434 $Y=0.234 $X2=0.351 $Y2=0.135
cc_181 N_8_c_310_p N_13_c_423_n 0.00116187f $X=0.459 $Y=0.225 $X2=0.351
+ $Y2=0.135
cc_182 N_8_c_291_n N_13_c_423_n 5.72158e-19 $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_183 N_9_M9_g N_10_M10_g 0.00268443f $X=0.783 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_184 N_9_c_315_p N_10_M10_g 3.74489e-19 $X=0.846 $Y=0.036 $X2=0.135 $Y2=0.054
cc_185 N_9_c_316_p N_10_c_370_n 0.00141609f $X=0.792 $Y=0.036 $X2=0.464
+ $Y2=0.178
cc_186 N_9_c_317_p N_10_c_362_n 0.00141609f $X=0.783 $Y=0.105 $X2=0 $Y2=0
cc_187 N_9_c_318_p N_10_c_340_n 3.34766e-19 $X=0.783 $Y=0.1055 $X2=0.071
+ $Y2=0.054
cc_188 N_9_c_317_p N_10_c_340_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.071
+ $Y2=0.054
cc_189 N_9_c_320_p N_10_c_343_n 2.41112e-19 $X=0.945 $Y=0.225 $X2=0 $Y2=0
cc_190 N_9_c_321_p N_10_c_375_n 2.65946e-19 $X=0.828 $Y=0.036 $X2=0.071
+ $Y2=0.216
cc_191 N_9_M9_g N_10_c_376_n 6.3699e-19 $X=0.783 $Y=0.0405 $X2=0.056 $Y2=0.216
cc_192 N_9_c_317_p N_10_c_376_n 9.10342e-19 $X=0.783 $Y=0.105 $X2=0.056
+ $Y2=0.216
cc_193 N_9_c_315_p N_10_c_378_n 4.40983e-19 $X=0.846 $Y=0.036 $X2=0.018 $Y2=0.18
cc_194 N_9_c_325_p N_10_c_379_n 5.181e-19 $X=0.882 $Y=0.036 $X2=0.027 $Y2=0.036
cc_195 N_9_c_326_p N_10_c_380_n 0.00149072f $X=0.9 $Y=0.234 $X2=0.054 $Y2=0.036
cc_196 N_9_c_327_p N_10_c_381_n 4.52584e-19 $X=0.9 $Y=0.036 $X2=0.135 $Y2=0.135
cc_197 N_9_c_328_p N_10_c_381_n 0.00299476f $X=0.945 $Y=0.167 $X2=0.135
+ $Y2=0.135
cc_198 N_9_c_329_p N_10_c_355_n 2.40515e-19 $X=0.936 $Y=0.036 $X2=0.145
+ $Y2=0.135
cc_199 N_9_c_330_p N_10_c_355_n 7.44774e-19 $X=0.918 $Y=0.234 $X2=0.145
+ $Y2=0.135
cc_200 N_9_c_328_p N_10_c_355_n 9.28741e-19 $X=0.945 $Y=0.167 $X2=0.145
+ $Y2=0.135
cc_201 N_9_c_332_p N_10_c_386_n 0.0032313f $X=0.945 $Y=0.117 $X2=0.033 $Y2=0.189
cc_202 N_9_c_329_p N_QN_c_403_n 4.62613e-19 $X=0.936 $Y=0.036 $X2=0 $Y2=0
cc_203 N_9_c_334_p N_QN_c_404_n 4.53762e-19 $X=0.936 $Y=0.234 $X2=0.459
+ $Y2=0.0405
cc_204 N_9_c_316_p N_14_c_432_n 7.33799e-19 $X=0.792 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_205 N_10_c_387_p N_QN_M12_d 3.80663e-19 $X=1.053 $Y=0.135 $X2=0.135 $Y2=0.054
cc_206 N_10_c_387_p N_QN_M25_d 3.78829e-19 $X=1.053 $Y=0.135 $X2=0.135 $Y2=0.216
cc_207 N_10_c_387_p N_QN_c_407_n 8.00061e-19 $X=1.053 $Y=0.135 $X2=0.351
+ $Y2=0.135
cc_208 N_10_M12_g N_QN_c_403_n 4.59284e-19 $X=1.053 $Y=0.0675 $X2=0 $Y2=0
cc_209 N_10_c_387_p N_QN_c_403_n 5.51214e-19 $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_210 N_10_c_387_p N_QN_c_410_n 8.00061e-19 $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_211 N_10_c_386_n N_QN_c_410_n 6.27102e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_212 N_10_M12_g N_QN_c_404_n 4.59284e-19 $X=1.053 $Y=0.0675 $X2=0.459
+ $Y2=0.0405
cc_213 N_10_c_387_p N_QN_c_404_n 5.49974e-19 $X=1.053 $Y=0.135 $X2=0.459
+ $Y2=0.0405
cc_214 N_10_c_387_p QN 3.92396e-19 $X=1.053 $Y=0.135 $X2=0.621 $Y2=0.178
cc_215 N_10_c_386_n N_QN_c_415_n 9.94215e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_216 N_10_c_337_n N_14_c_432_n 0.00182708f $X=0.648 $Y=0.0405 $X2=0.351
+ $Y2=0.135
cc_217 N_10_c_370_n N_14_c_432_n 0.00205226f $X=0.72 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_218 N_10_c_400_p N_14_c_432_n 0.0013184f $X=0.704 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_219 N_10_c_362_n N_14_c_432_n 0.00103589f $X=0.729 $Y=0.081 $X2=0.351
+ $Y2=0.135
cc_220 N_10_c_345_n N_14_c_432_n 4.02739e-19 $X=0.774 $Y=0.162 $X2=0.351
+ $Y2=0.135

* END of "./DFFLQNx2_ASAP7_75t_SRAM.pex.sp.DFFLQNX2_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DFFLQNx3_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:26:23 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DFFLQNx3_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DFFLQNx3_ASAP7_75t_SRAM.pex.sp.pex"
* File: DFFLQNx3_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:26:23 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%CLK 2 5 7 12 14 17 VSS
c18 17 VSS 1.44512e-20 $X=0.081 $Y=0.1305
c19 14 VSS 0.00705007f $X=0.081 $Y=0.135
c20 12 VSS 0.00709305f $X=0.082 $Y=0.119
c21 5 VSS 0.00184374f $X=0.081 $Y=0.135
c22 2 VSS 0.0629f $X=0.081 $Y=0.054
r23 16 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r24 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r25 12 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.126
r26 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%4 2 5 7 10 13 16 22 25 28 31 36 43 47 50 52 58
+ 59 60 64 67 74 79 84 88 89 92 96 99 100 101 103 111 124 132 148 VSS
c102 148 VSS 4.19842e-19 $X=0.18 $Y=0.189
c103 147 VSS 1.53928e-19 $X=0.189 $Y=0.189
c104 141 VSS 7.0154e-20 $X=0.03 $Y=0.189
c105 140 VSS 5.9624e-19 $X=0.027 $Y=0.189
c106 124 VSS 6.81413e-19 $X=0.513 $Y=0.18
c107 111 VSS 4.0846e-19 $X=0.351 $Y=0.135
c108 103 VSS 0.00656068f $X=0.513 $Y=0.189
c109 101 VSS 0.00251877f $X=0.29 $Y=0.189
c110 100 VSS 0.00602789f $X=0.229 $Y=0.189
c111 99 VSS 7.60117e-19 $X=0.351 $Y=0.189
c112 96 VSS 4.13996e-19 $X=0.159 $Y=0.189
c113 92 VSS 4.95554e-19 $X=0.033 $Y=0.189
c114 89 VSS 7.37649e-20 $X=0.189 $Y=0.172
c115 88 VSS 5.63427e-19 $X=0.189 $Y=0.164
c116 87 VSS 1.04741e-19 $X=0.189 $Y=0.18
c117 85 VSS 9.32637e-20 $X=0.148 $Y=0.135
c118 84 VSS 9.68735e-19 $X=0.145 $Y=0.135
c119 79 VSS 0.00149077f $X=0.18 $Y=0.135
c120 77 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c121 76 VSS 0.00169428f $X=0.047 $Y=0.234
c122 74 VSS 0.00250477f $X=0.054 $Y=0.234
c123 72 VSS 0.00306385f $X=0.027 $Y=0.234
c124 70 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c125 69 VSS 0.00205521f $X=0.047 $Y=0.036
c126 67 VSS 0.00250477f $X=0.054 $Y=0.036
c127 65 VSS 0.00305101f $X=0.027 $Y=0.036
c128 64 VSS 4.99402e-19 $X=0.018 $Y=0.2125
c129 63 VSS 1.14289e-19 $X=0.018 $Y=0.2
c130 62 VSS 4.86272e-19 $X=0.018 $Y=0.225
c131 60 VSS 0.00271341f $X=0.018 $Y=0.125
c132 59 VSS 9.57865e-19 $X=0.018 $Y=0.07
c133 58 VSS 0.00235012f $X=0.018 $Y=0.18
c134 55 VSS 0.00530434f $X=0.056 $Y=0.216
c135 52 VSS 2.98509e-19 $X=0.071 $Y=0.216
c136 50 VSS 0.00492487f $X=0.056 $Y=0.054
c137 47 VSS 2.98509e-19 $X=0.071 $Y=0.054
c138 43 VSS 0.0585267f $X=0.725 $Y=0.178
c139 36 VSS 0.00123999f $X=0.464 $Y=0.178
c140 28 VSS 0.0616846f $X=0.729 $Y=0.178
c141 25 VSS 1.44609e-19 $X=0.621 $Y=0.178
c142 22 VSS 0.0600171f $X=0.621 $Y=0.0405
c143 16 VSS 0.0602253f $X=0.459 $Y=0.0405
c144 10 VSS 0.0608611f $X=0.351 $Y=0.135
c145 5 VSS 0.00277501f $X=0.135 $Y=0.135
c146 2 VSS 0.0623856f $X=0.135 $Y=0.054
r147 148 149 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.189 $X2=0.1845 $Y2=0.189
r148 147 149 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.189 $X2=0.1845 $Y2=0.189
r149 140 141 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.03 $Y2=0.189
r150 137 140 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.027 $Y2=0.189
r151 131 132 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.351 $Y=0.167 $X2=0.351 $Y2=0.178
r152 123 124 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r153 111 131 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.167
r154 103 124 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r155 100 101 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.189 $X2=0.29 $Y2=0.189
r156 99 132 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.178
r157 98 103 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.513 $Y2=0.189
r158 98 101 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.29 $Y2=0.189
r159 98 99 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.189 $X2=0.351
+ $Y2=0.189
r160 96 148 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.159
+ $Y=0.189 $X2=0.18 $Y2=0.189
r161 95 100 4.75309 $w=1.8e-08 $l=7e-08 $layer=M2 $thickness=3.6e-08 $X=0.159
+ $Y=0.189 $X2=0.229 $Y2=0.189
r162 95 96 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.159 $Y=0.189 $X2=0.159
+ $Y2=0.189
r163 92 141 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.03 $Y2=0.189
r164 91 95 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.159 $Y2=0.189
r165 91 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.189 $X2=0.033
+ $Y2=0.189
r166 88 89 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.172
r167 87 147 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.189
r168 87 89 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.172
r169 86 88 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.164
r170 84 85 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.145
+ $Y=0.135 $X2=0.148 $Y2=0.135
r171 81 84 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.145 $Y2=0.135
r172 79 86 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r173 79 85 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.148 $Y2=0.135
r174 76 77 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r175 74 77 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r176 72 76 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r177 69 70 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r178 67 70 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r179 65 69 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r180 63 64 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r181 62 72 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r182 62 64 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r183 61 137 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.189
r184 61 63 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.2
r185 59 60 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.125
r186 58 137 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.189
r187 58 60 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.125
r188 57 65 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r189 57 59 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r190 55 74 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r191 52 55 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r192 50 67 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r193 47 50 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r194 36 123 39.0385 $w=2.6e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.178 $X2=0.513 $Y2=0.178
r195 28 43 3.07692 $w=2.6e-08 $l=4e-09 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.178 $X2=0.725 $Y2=0.178
r196 28 31 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.178 $X2=0.729 $Y2=0.2295
r197 25 43 82.8571 $w=2.6e-08 $l=1.04e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.725 $Y2=0.178
r198 25 123 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.513 $Y2=0.178
r199 22 25 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0405 $X2=0.621 $Y2=0.178
r200 19 36 3.84615 $w=2.6e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.178 $X2=0.464 $Y2=0.178
r201 16 19 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.178
r202 10 111 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135
+ $X2=0.351 $Y2=0.135
r203 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r204 5 81 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r205 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r206 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%D 2 5 7 12 14 17 VSS
c21 17 VSS 2.32756e-19 $X=0.297 $Y=0.126
c22 14 VSS 0.0072156f $X=0.297 $Y=0.135
c23 12 VSS 0.00703905f $X=0.298 $Y=0.082
c24 5 VSS 0.00200686f $X=0.297 $Y=0.135
c25 2 VSS 0.061556f $X=0.297 $Y=0.0675
r26 16 17 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.126
r27 14 17 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.126
r28 12 16 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.082 $X2=0.297 $Y2=0.106
r29 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r30 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r31 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%6 2 5 7 10 13 15 17 22 25 27 32 34 39 40 42 45
+ 51 53 54 58 63 73 74 76 VSS
c70 76 VSS 7.89434e-19 $X=0.243 $Y=0.2115
c71 74 VSS 9.16337e-19 $X=0.243 $Y=0.126
c72 73 VSS 0.00233088f $X=0.243 $Y=0.106
c73 63 VSS 0.00103743f $X=0.675 $Y=0.135
c74 58 VSS 9.14968e-19 $X=0.405 $Y=0.135
c75 54 VSS 0.00260015f $X=0.601 $Y=0.153
c76 53 VSS 0.00786313f $X=0.527 $Y=0.153
c77 51 VSS 0.00404346f $X=0.675 $Y=0.153
c78 45 VSS 0.00167753f $X=0.243 $Y=0.153
c79 42 VSS 5.5218e-19 $X=0.243 $Y=0.225
c80 40 VSS 0.00181981f $X=0.216 $Y=0.234
c81 39 VSS 0.00525711f $X=0.198 $Y=0.234
c82 34 VSS 0.00482554f $X=0.234 $Y=0.234
c83 33 VSS 0.00200074f $X=0.216 $Y=0.036
c84 32 VSS 0.00545403f $X=0.198 $Y=0.036
c85 27 VSS 0.00500597f $X=0.234 $Y=0.036
c86 25 VSS 0.00648533f $X=0.16 $Y=0.216
c87 20 VSS 0.00602272f $X=0.16 $Y=0.054
c88 13 VSS 0.0021498f $X=0.675 $Y=0.135
c89 10 VSS 0.0585656f $X=0.675 $Y=0.0405
c90 5 VSS 0.00163668f $X=0.405 $Y=0.135
c91 2 VSS 0.058827f $X=0.405 $Y=0.0675
r92 75 76 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.198 $X2=0.243 $Y2=0.2115
r93 73 74 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.106 $X2=0.243 $Y2=0.126
r94 53 54 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.601 $Y2=0.153
r95 51 54 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.675
+ $Y=0.153 $X2=0.601 $Y2=0.153
r96 51 63 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.675 $Y=0.153 $X2=0.675
+ $Y2=0.153
r97 48 53 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.527 $Y2=0.153
r98 48 58 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r99 45 75 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.198
r100 45 74 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.126
r101 44 48 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.405 $Y2=0.153
r102 44 45 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.153 $X2=0.243
+ $Y2=0.153
r103 42 76 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.2115
r104 41 73 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.106
r105 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.216 $Y2=0.234
r106 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.198 $Y2=0.234
r107 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r108 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r109 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.216 $Y2=0.036
r110 29 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r111 27 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r112 27 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r113 25 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r114 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r115 20 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r116 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r117 13 63 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.135 $X2=0.675
+ $Y2=0.135
r118 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2295
r119 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.135
r120 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r121 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2295
r122 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%7 2 5 7 9 10 13 14 17 19 22 29 30 31 33 40 47 48
+ 49 50 51 52 54 55 VSS
c45 56 VSS 3.57489e-19 $X=0.612 $Y=0.09
c46 55 VSS 1.84136e-19 $X=0.603 $Y=0.09
c47 54 VSS 5.96246e-19 $X=0.621 $Y=0.09
c48 52 VSS 4.34894e-19 $X=0.621 $Y=0.214
c49 51 VSS 4.90038e-19 $X=0.621 $Y=0.203
c50 50 VSS 1.59683e-19 $X=0.621 $Y=0.167
c51 49 VSS 2.90654e-19 $X=0.621 $Y=0.165
c52 48 VSS 3.07094e-19 $X=0.621 $Y=0.14
c53 47 VSS 3.66508e-19 $X=0.621 $Y=0.122
c54 46 VSS 3.22511e-19 $X=0.621 $Y=0.225
c55 40 VSS 0.00154565f $X=0.594 $Y=0.054
c56 33 VSS 0.00268134f $X=0.594 $Y=0.234
c57 31 VSS 0.00427376f $X=0.612 $Y=0.234
c58 30 VSS 1.96699e-19 $X=0.583 $Y=0.09
c59 29 VSS 0.00266746f $X=0.581 $Y=0.09
c60 24 VSS 5.17345e-20 $X=0.585 $Y=0.09
c61 22 VSS 0.0179398f $X=0.65 $Y=0.2295
c62 19 VSS 3.14771e-19 $X=0.665 $Y=0.2295
c63 17 VSS 2.5391e-19 $X=0.592 $Y=0.2295
c64 13 VSS 0.0281519f $X=0.594 $Y=0.0405
c65 9 VSS 6.29543e-19 $X=0.611 $Y=0.0405
c66 5 VSS 0.00233073f $X=0.513 $Y=0.09
c67 2 VSS 0.0584396f $X=0.513 $Y=0.0405
r68 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.603
+ $Y=0.09 $X2=0.612 $Y2=0.09
r69 54 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.612 $Y2=0.09
r70 53 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.09 $X2=0.603 $Y2=0.09
r71 51 52 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.214
r72 50 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.203
r73 49 50 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.167
r74 48 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r75 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r76 46 52 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.214
r77 45 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.09
r78 45 47 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.122
r79 38 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.09
r80 38 40 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.054
r81 31 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r82 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r83 29 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.581
+ $Y=0.09 $X2=0.583 $Y2=0.09
r84 26 29 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.09 $X2=0.581 $Y2=0.09
r85 24 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.594 $Y2=0.09
r86 24 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.583 $Y2=0.09
r87 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2295 $X2=0.65 $Y2=0.2295
r88 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.592
+ $Y=0.2295 $X2=0.65 $Y2=0.2295
r89 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r90 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r91 13 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.054 $X2=0.594
+ $Y2=0.054
r92 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.594 $Y2=0.0405
r93 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0405 $X2=0.594 $Y2=0.0405
r94 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.09 $X2=0.513
+ $Y2=0.09
r95 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.09 $X2=0.513 $Y2=0.2295
r96 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.09
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%8 2 5 7 9 14 17 21 22 25 30 31 33 35 36 37 38 39
+ 41 42 43 44 48 50 51 52 53 58 60 61 VSS
c55 64 VSS 2.84134e-19 $X=0.459 $Y=0.131
c56 61 VSS 0.00334468f $X=0.45 $Y=0.036
c57 60 VSS 0.00243127f $X=0.459 $Y=0.036
c58 58 VSS 0.00276391f $X=0.432 $Y=0.036
c59 53 VSS 4.23521e-19 $X=0.5445 $Y=0.131
c60 52 VSS 3.49205e-20 $X=0.522 $Y=0.131
c61 51 VSS 2.00095e-19 $X=0.504 $Y=0.131
c62 50 VSS 0.00133241f $X=0.496 $Y=0.131
c63 48 VSS 5.65734e-19 $X=0.567 $Y=0.131
c64 45 VSS 4.53296e-19 $X=0.459 $Y=0.214
c65 44 VSS 2.01779e-19 $X=0.459 $Y=0.203
c66 43 VSS 6.09344e-21 $X=0.459 $Y=0.167
c67 42 VSS 1.60693e-19 $X=0.459 $Y=0.165
c68 41 VSS 3.22878e-19 $X=0.459 $Y=0.225
c69 39 VSS 2.48018e-19 $X=0.459 $Y=0.114
c70 38 VSS 2.26591e-19 $X=0.459 $Y=0.106
c71 37 VSS 9.45429e-20 $X=0.459 $Y=0.099
c72 36 VSS 8.12259e-19 $X=0.459 $Y=0.081
c73 35 VSS 2.08428e-19 $X=0.459 $Y=0.122
c74 33 VSS 0.00142907f $X=0.434 $Y=0.234
c75 32 VSS 3.66528e-19 $X=0.418 $Y=0.234
c76 31 VSS 0.00146362f $X=0.414 $Y=0.234
c77 30 VSS 0.00368178f $X=0.396 $Y=0.234
c78 25 VSS 0.00389542f $X=0.45 $Y=0.234
c79 24 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c80 21 VSS 0.00348256f $X=0.378 $Y=0.2025
c81 16 VSS 5.70081e-19 $X=0.432 $Y=0.0405
c82 5 VSS 0.00195718f $X=0.567 $Y=0.1305
c83 2 VSS 0.0591962f $X=0.567 $Y=0.0405
r84 61 62 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r85 60 62 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r86 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r87 57 58 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r88 52 53 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r89 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r90 50 51 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.496
+ $Y=0.131 $X2=0.504 $Y2=0.131
r91 48 53 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r92 46 64 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r93 46 50 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.496 $Y2=0.131
r94 44 45 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.203 $X2=0.459 $Y2=0.214
r95 43 44 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.167 $X2=0.459 $Y2=0.203
r96 42 43 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.167
r97 41 45 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r98 40 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r99 40 42 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.165
r100 38 39 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.106 $X2=0.459 $Y2=0.114
r101 37 38 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.099 $X2=0.459 $Y2=0.106
r102 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.099
r103 35 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r104 35 39 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.114
r105 34 60 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r106 34 36 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.081
r107 32 33 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.234 $X2=0.434 $Y2=0.234
r108 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.418 $Y2=0.234
r109 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r110 27 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r111 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r112 25 33 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.434 $Y2=0.234
r113 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r114 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r115 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r116 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r117 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r118 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r119 13 58 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r120 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r121 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r122 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r123 5 48 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.131 $X2=0.567
+ $Y2=0.131
r124 5 7 370.904 $w=2e-08 $l=9.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1305 $X2=0.567 $Y2=0.2295
r125 2 5 337.185 $w=2e-08 $l=9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.1305
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%9 2 5 7 9 14 21 25 26 30 31 32 33 34 39 40 42 44
+ 45 VSS
c24 46 VSS 1.88981e-19 $X=0.945 $Y=0.171
c25 45 VSS 0.00101091f $X=0.945 $Y=0.167
c26 44 VSS 8.83619e-19 $X=0.945 $Y=0.117
c27 43 VSS 0.00236812f $X=0.945 $Y=0.09
c28 42 VSS 0.00301787f $X=0.945 $Y=0.225
c29 40 VSS 0.0018377f $X=0.918 $Y=0.234
c30 39 VSS 0.0056872f $X=0.9 $Y=0.234
c31 34 VSS 0.00462933f $X=0.936 $Y=0.234
c32 33 VSS 0.00189638f $X=0.9 $Y=0.036
c33 32 VSS 0.00352438f $X=0.882 $Y=0.036
c34 31 VSS 0.00146362f $X=0.846 $Y=0.036
c35 30 VSS 0.00508235f $X=0.828 $Y=0.036
c36 26 VSS 0.00226308f $X=0.792 $Y=0.036
c37 25 VSS 0.00657044f $X=0.936 $Y=0.036
c38 21 VSS 0.00122443f $X=0.783 $Y=0.105
c39 17 VSS 0.0048151f $X=0.862 $Y=0.2295
c40 12 VSS 0.00513461f $X=0.862 $Y=0.0405
c41 5 VSS 0.00277722f $X=0.783 $Y=0.1055
c42 2 VSS 0.0590816f $X=0.783 $Y=0.0405
r43 45 46 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.167 $X2=0.945 $Y2=0.171
r44 44 45 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.117 $X2=0.945 $Y2=0.167
r45 43 44 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.09 $X2=0.945 $Y2=0.117
r46 42 46 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.171
r47 41 43 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.09
r48 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.234 $X2=0.918 $Y2=0.234
r49 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.9 $Y2=0.234
r50 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r51 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.918 $Y2=0.234
r52 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r53 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.846 $Y2=0.036
r54 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r55 28 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.846 $Y2=0.036
r56 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.036 $X2=0.828 $Y2=0.036
r57 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r58 25 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.9 $Y2=0.036
r59 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.783 $Y=0.045 $X2=0.792 $Y2=0.036
r60 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.105
r61 17 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234 $X2=0.864
+ $Y2=0.234
r62 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2295 $X2=0.862 $Y2=0.2295
r63 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036 $X2=0.864
+ $Y2=0.036
r64 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.862 $Y2=0.0405
r65 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.105 $X2=0.783
+ $Y2=0.105
r66 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.1055 $X2=0.783 $Y2=0.2295
r67 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.1055
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%10 2 7 10 15 18 23 26 29 31 33 34 37 38 39 42 43
+ 48 49 51 53 54 55 56 57 59 60 62 63 66 73 74 82 85 89 92 100 VSS
c69 100 VSS 0.00217412f $X=0.999 $Y=0.136
c70 92 VSS 0.00790847f $X=0.999 $Y=0.153
c71 89 VSS 0.00149614f $X=0.891 $Y=0.153
c72 86 VSS 4.17512e-19 $X=0.837 $Y=0.162
c73 85 VSS 1.52743e-19 $X=0.729 $Y=0.162
c74 82 VSS 0.00370746f $X=0.72 $Y=0.234
c75 81 VSS 0.00266816f $X=0.729 $Y=0.234
c76 74 VSS 4.30636e-19 $X=0.866 $Y=0.162
c77 73 VSS 1.48695e-19 $X=0.85 $Y=0.162
c78 71 VSS 2.75449e-19 $X=0.882 $Y=0.162
c79 66 VSS 3.94906e-19 $X=0.837 $Y=0.135
c80 63 VSS 3.26354e-19 $X=0.792 $Y=0.162
c81 62 VSS 0.00206921f $X=0.774 $Y=0.162
c82 60 VSS 0.00192346f $X=0.828 $Y=0.162
c83 59 VSS 0.00136716f $X=0.729 $Y=0.225
c84 57 VSS 1.52884e-19 $X=0.729 $Y=0.136
c85 56 VSS 9.59255e-20 $X=0.729 $Y=0.119
c86 55 VSS 1.29374e-19 $X=0.729 $Y=0.099
c87 54 VSS 3.52175e-19 $X=0.729 $Y=0.081
c88 53 VSS 2.74133e-19 $X=0.729 $Y=0.153
c89 51 VSS 0.00166816f $X=0.704 $Y=0.036
c90 50 VSS 4.57836e-19 $X=0.688 $Y=0.036
c91 49 VSS 0.00146362f $X=0.684 $Y=0.036
c92 48 VSS 0.00370471f $X=0.666 $Y=0.036
c93 43 VSS 0.00409787f $X=0.72 $Y=0.036
c94 42 VSS 0.00276615f $X=0.702 $Y=0.2295
c95 38 VSS 5.63046e-19 $X=0.719 $Y=0.2295
c96 37 VSS 0.0349304f $X=0.648 $Y=0.0405
c97 33 VSS 5.63046e-19 $X=0.665 $Y=0.0405
c98 29 VSS 0.0132556f $X=1.107 $Y=0.136
c99 26 VSS 0.0647964f $X=1.107 $Y=0.0675
c100 18 VSS 0.0617066f $X=1.053 $Y=0.0675
c101 10 VSS 0.0610431f $X=0.999 $Y=0.0675
c102 5 VSS 0.00189441f $X=0.837 $Y=0.135
c103 2 VSS 0.0618222f $X=0.837 $Y=0.0405
r104 92 100 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.999 $Y=0.153 $X2=0.999
+ $Y2=0.153
r105 88 92 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.999 $Y2=0.153
r106 88 89 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r107 82 83 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.234 $X2=0.7245 $Y2=0.234
r108 81 83 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.234 $X2=0.7245 $Y2=0.234
r109 78 82 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.234 $X2=0.72 $Y2=0.234
r110 73 74 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.85
+ $Y=0.162 $X2=0.866 $Y2=0.162
r111 72 86 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.837 $Y2=0.162
r112 72 73 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.85 $Y2=0.162
r113 71 89 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.891 $Y2=0.162
r114 71 74 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.866 $Y2=0.162
r115 64 86 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.162
r116 64 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.135
r117 62 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.162 $X2=0.792 $Y2=0.162
r118 61 85 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.729 $Y2=0.162
r119 61 62 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.774 $Y2=0.162
r120 60 86 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.837 $Y2=0.162
r121 60 63 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.792 $Y2=0.162
r122 59 81 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.225 $X2=0.729 $Y2=0.234
r123 58 85 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.162
r124 58 59 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.225
r125 56 57 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.119 $X2=0.729 $Y2=0.136
r126 55 56 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.099 $X2=0.729 $Y2=0.119
r127 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.081 $X2=0.729 $Y2=0.099
r128 53 85 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.162
r129 53 57 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.136
r130 52 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.045 $X2=0.729 $Y2=0.081
r131 50 51 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.036 $X2=0.704 $Y2=0.036
r132 49 50 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.688 $Y2=0.036
r133 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.684 $Y2=0.036
r134 45 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.666 $Y2=0.036
r135 43 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.036 $X2=0.729 $Y2=0.045
r136 43 51 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.704 $Y2=0.036
r137 42 78 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.234
+ $X2=0.702 $Y2=0.234
r138 39 42 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2295 $X2=0.702 $Y2=0.2295
r139 38 42 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2295 $X2=0.702 $Y2=0.2295
r140 37 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r141 34 37 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0405 $X2=0.648 $Y2=0.0405
r142 33 37 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r143 29 31 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.136 $X2=1.107 $Y2=0.2025
r144 26 29 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.0675 $X2=1.107 $Y2=0.136
r145 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.053
+ $Y=0.136 $X2=1.107 $Y2=0.136
r146 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.136 $X2=1.053 $Y2=0.2025
r147 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.0675 $X2=1.053 $Y2=0.136
r148 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.999
+ $Y=0.136 $X2=1.053 $Y2=0.136
r149 13 100 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.136
+ $X2=0.999 $Y2=0.136
r150 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.136 $X2=0.999 $Y2=0.2025
r151 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.136
r152 5 66 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.135 $X2=0.837
+ $Y2=0.135
r153 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.2295
r154 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.0405 $X2=0.837 $Y2=0.135
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%QN 1 2 6 11 12 15 16 21 23 24 31 42 44 VSS
c15 46 VSS 0.00143312f $X=1.162 $Y=0.196
c16 44 VSS 9.70664e-19 $X=1.162 $Y=0.1095
c17 43 VSS 0.00218124f $X=1.162 $Y=0.09
c18 42 VSS 0.00322575f $X=1.161 $Y=0.129
c19 40 VSS 0.00139892f $X=1.162 $Y=0.225
c20 31 VSS 0.0196976f $X=1.153 $Y=0.234
c21 30 VSS 0.00635401f $X=1.134 $Y=0.036
c22 24 VSS 0.0096322f $X=1.026 $Y=0.036
c23 23 VSS 0.00148748f $X=1.026 $Y=0.036
c24 21 VSS 0.0182937f $X=1.153 $Y=0.036
c25 19 VSS 0.00670088f $X=1.132 $Y=0.2025
c26 15 VSS 0.00940513f $X=1.026 $Y=0.2025
c27 11 VSS 5.72268e-19 $X=1.043 $Y=0.2025
c28 9 VSS 3.44349e-19 $X=1.132 $Y=0.0675
c29 1 VSS 5.4768e-19 $X=1.043 $Y=0.0675
r30 45 46 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.167 $X2=1.162 $Y2=0.196
r31 43 44 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.09 $X2=1.162 $Y2=0.1095
r32 42 45 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.129 $X2=1.162 $Y2=0.167
r33 42 44 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.129 $X2=1.162 $Y2=0.1095
r34 40 46 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.225 $X2=1.162 $Y2=0.196
r35 39 43 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.162
+ $Y=0.045 $X2=1.162 $Y2=0.09
r36 33 37 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.234 $X2=1.134 $Y2=0.234
r37 31 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.153 $Y=0.234 $X2=1.162 $Y2=0.225
r38 31 37 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.153
+ $Y=0.234 $X2=1.134 $Y2=0.234
r39 29 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.134 $Y=0.036 $X2=1.134
+ $Y2=0.036
r40 23 29 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.036 $X2=1.134 $Y2=0.036
r41 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.036 $X2=1.026
+ $Y2=0.036
r42 21 39 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.153 $Y=0.036 $X2=1.162 $Y2=0.045
r43 21 29 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.153
+ $Y=0.036 $X2=1.134 $Y2=0.036
r44 19 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.134 $Y=0.234 $X2=1.134
+ $Y2=0.234
r45 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.117 $Y=0.2025 $X2=1.132 $Y2=0.2025
r46 15 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.234 $X2=1.026
+ $Y2=0.234
r47 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.2025 $X2=1.026 $Y2=0.2025
r48 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.043 $Y=0.2025 $X2=1.026 $Y2=0.2025
r49 9 30 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.134
+ $Y=0.0675 $X2=1.134 $Y2=0.036
r50 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.117
+ $Y=0.0675 $X2=1.132 $Y2=0.0675
r51 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.026
+ $Y=0.0675 $X2=1.026 $Y2=0.036
r52 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.009
+ $Y=0.0675 $X2=1.026 $Y2=0.0675
r53 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.043
+ $Y=0.0675 $X2=1.026 $Y2=0.0675
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%12 1 6 9 VSS
c6 9 VSS 0.0266112f $X=0.38 $Y=0.0675
c7 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c8 4 VSS 3.22674e-19 $X=0.322 $Y=0.0675
r9 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r10 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%13 1 6 9 VSS
c10 9 VSS 0.0209308f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.69239e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%14 1 6 9 VSS
c8 9 VSS 0.0191793f $X=0.758 $Y=0.0405
c9 6 VSS 3.14771e-19 $X=0.773 $Y=0.0405
c10 4 VSS 2.61968e-19 $X=0.7 $Y=0.0405
r11 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r12 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.7
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r13 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.685
+ $Y=0.0405 $X2=0.7 $Y2=0.0405
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%15 1 2 VSS
c0 1 VSS 0.00225696f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%16 1 2 VSS
c1 1 VSS 0.00201018f $X=0.341 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends

.subckt PM_DFFLQNX3_ASAP7_75T_SRAM%17 1 2 VSS
c0 1 VSS 0.00219822f $X=0.773 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2295 $X2=0.739 $Y2=0.2295
.ends


* END of "./DFFLQNx3_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DFFLQNx3_ASAP7_75t_SRAM  VSS VDD CLK D QN
* 
* QN	QN
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_12_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_6_M3_g N_12_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_15_M4_d N_4_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_15_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_10_M7_d N_4_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.611
+ $Y=0.027
M8 N_14_M8_d N_6_M8_g N_10_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M9 VSS N_9_M9_g N_14_M9_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_9_M10_d N_10_M10_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.027
M11 N_QN_M11_d N_10_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M12 N_QN_M12_d N_10_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.027
M13 N_QN_M13_d N_10_M13_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.027
M14 VDD N_CLK_M14_g N_4_M14_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M15 N_6_M15_d N_4_M15_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M16 N_16_M16_d N_D_M16_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M17 N_8_M17_d N_4_M17_g N_16_M17_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M18 N_13_M18_d N_6_M18_g N_8_M18_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M19 VDD N_7_M19_g N_13_M19_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M20 N_7_M20_d N_8_M20_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M21 N_10_M21_d N_6_M21_g N_7_M21_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.665 $Y=0.216
M22 N_17_M22_d N_4_M22_g N_10_M22_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.719 $Y=0.216
M23 VDD N_9_M23_g N_17_M23_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M24 N_9_M24_d N_10_M24_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.216
M25 N_QN_M25_d N_10_M25_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
M26 N_QN_M26_d N_10_M26_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.162
M27 N_QN_M27_d N_10_M27_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.162
*
* 
* .include "DFFLQNx3_ASAP7_75t_SRAM.pex.sp.DFFLQNX3_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DFFLQNx3_ASAP7_75t_SRAM.pex.sp.DFFLQNX3_ASAP7_75T_SRAM.pxi"
* File: DFFLQNx3_ASAP7_75t_SRAM.pex.sp.DFFLQNX3_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:26:23 2017
* 
x_PM_DFFLQNX3_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M14_g CLK N_CLK_c_4_p
+ N_CLK_c_10_p VSS PM_DFFLQNX3_ASAP7_75T_SRAM%CLK
x_PM_DFFLQNX3_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_20_n N_4_M15_g N_4_c_34_p N_4_M17_g
+ N_4_M4_g N_4_M7_g N_4_c_77_p N_4_c_43_p N_4_M22_g N_4_c_89_p N_4_c_44_p
+ N_4_M0_s N_4_c_21_n N_4_M14_s N_4_c_22_n N_4_c_23_n N_4_c_24_n N_4_c_25_n
+ N_4_c_26_n N_4_c_27_n N_4_c_47_p N_4_c_28_n N_4_c_29_n N_4_c_30_n N_4_c_31_n
+ N_4_c_32_n N_4_c_58_p N_4_c_33_n N_4_c_36_p N_4_c_37_p N_4_c_38_p N_4_c_61_p
+ N_4_c_94_p N_4_c_46_p VSS PM_DFFLQNX3_ASAP7_75T_SRAM%4
x_PM_DFFLQNX3_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_122_n N_D_M16_g D N_D_c_123_n
+ N_D_c_133_p VSS PM_DFFLQNX3_ASAP7_75T_SRAM%D
x_PM_DFFLQNX3_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_147_n N_6_M18_g N_6_M8_g N_6_c_151_n
+ N_6_M21_g N_6_M1_d N_6_M15_d N_6_c_152_n N_6_c_172_n N_6_c_142_n N_6_c_154_n
+ N_6_c_143_n N_6_c_158_n N_6_c_174_n N_6_c_159_n N_6_c_161_n N_6_c_162_n
+ N_6_c_183_p N_6_c_168_n N_6_c_170_n N_6_c_144_n N_6_c_180_n N_6_c_181_n VSS
+ PM_DFFLQNX3_ASAP7_75T_SRAM%6
x_PM_DFFLQNX3_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_237_p N_7_M19_g N_7_M7_s N_7_M6_d
+ N_7_c_216_n N_7_M20_d N_7_c_217_n N_7_M21_s N_7_c_219_n N_7_c_235_p
+ N_7_c_228_n N_7_c_255_p N_7_c_229_n N_7_c_236_p N_7_c_221_n N_7_c_240_p
+ N_7_c_222_n N_7_c_223_n N_7_c_224_n N_7_c_253_p N_7_c_226_n N_7_c_233_n VSS
+ PM_DFFLQNX3_ASAP7_75T_SRAM%7
x_PM_DFFLQNX3_ASAP7_75T_SRAM%8 N_8_M6_g N_8_c_280_n N_8_M20_g N_8_M3_d N_8_M4_s
+ N_8_M17_d N_8_c_260_n N_8_M18_s N_8_c_308_p N_8_c_262_n N_8_c_283_n
+ N_8_c_309_p N_8_c_285_n N_8_c_263_n N_8_c_264_n N_8_c_298_n N_8_c_286_n
+ N_8_c_310_p N_8_c_265_n N_8_c_266_n N_8_c_268_n N_8_c_299_n N_8_c_272_n
+ N_8_c_300_n N_8_c_273_n N_8_c_275_n N_8_c_291_n N_8_c_303_n N_8_c_278_n VSS
+ PM_DFFLQNX3_ASAP7_75T_SRAM%8
x_PM_DFFLQNX3_ASAP7_75T_SRAM%9 N_9_M9_g N_9_c_318_p N_9_M23_g N_9_M10_d N_9_M24_d
+ N_9_c_317_p N_9_c_329_p N_9_c_316_p N_9_c_321_p N_9_c_315_p N_9_c_325_p
+ N_9_c_327_p N_9_c_334_p N_9_c_326_p N_9_c_330_p N_9_c_320_p N_9_c_332_p
+ N_9_c_328_p VSS PM_DFFLQNX3_ASAP7_75T_SRAM%9
x_PM_DFFLQNX3_ASAP7_75T_SRAM%10 N_10_M10_g N_10_M24_g N_10_M11_g N_10_M25_g
+ N_10_M12_g N_10_M26_g N_10_M13_g N_10_c_387_p N_10_M27_g N_10_M8_s N_10_M7_d
+ N_10_c_337_n N_10_M22_s N_10_M21_d N_10_c_339_n N_10_c_370_n N_10_c_350_n
+ N_10_c_351_n N_10_c_402_p N_10_c_353_n N_10_c_362_n N_10_c_340_n N_10_c_341_n
+ N_10_c_342_n N_10_c_343_n N_10_c_375_n N_10_c_345_n N_10_c_376_n N_10_c_378_n
+ N_10_c_379_n N_10_c_380_n N_10_c_346_n N_10_c_347_n N_10_c_381_n N_10_c_355_n
+ N_10_c_386_n VSS PM_DFFLQNX3_ASAP7_75T_SRAM%10
x_PM_DFFLQNX3_ASAP7_75T_SRAM%QN N_QN_M12_d N_QN_M11_d N_QN_M13_d N_QN_M26_d
+ N_QN_M25_d N_QN_c_409_n N_QN_M27_d N_QN_c_410_n N_QN_c_405_n N_QN_c_413_n
+ N_QN_c_406_n QN N_QN_c_419_n VSS PM_DFFLQNX3_ASAP7_75T_SRAM%QN
x_PM_DFFLQNX3_ASAP7_75T_SRAM%12 N_12_M2_d N_12_M3_s N_12_c_420_n VSS
+ PM_DFFLQNX3_ASAP7_75T_SRAM%12
x_PM_DFFLQNX3_ASAP7_75T_SRAM%13 N_13_M18_d N_13_M19_s N_13_c_427_n VSS
+ PM_DFFLQNX3_ASAP7_75T_SRAM%13
x_PM_DFFLQNX3_ASAP7_75T_SRAM%14 N_14_M8_d N_14_M9_s N_14_c_436_n VSS
+ PM_DFFLQNX3_ASAP7_75T_SRAM%14
x_PM_DFFLQNX3_ASAP7_75T_SRAM%15 N_15_M5_s N_15_M4_d VSS PM_DFFLQNX3_ASAP7_75T_SRAM%15
x_PM_DFFLQNX3_ASAP7_75T_SRAM%16 N_16_M17_s N_16_M16_d VSS
+ PM_DFFLQNX3_ASAP7_75T_SRAM%16
x_PM_DFFLQNX3_ASAP7_75T_SRAM%17 N_17_M23_s N_17_M22_d VSS
+ PM_DFFLQNX3_ASAP7_75T_SRAM%17
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_CLK_c_2_p N_4_c_20_n 0.00124017f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 CLK N_4_c_21_n 3.57152e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_4 N_CLK_c_4_p N_4_c_22_n 0.00206543f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.18
cc_5 CLK N_4_c_23_n 2.75361e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.07
cc_6 CLK N_4_c_24_n 0.00206543f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.125
cc_7 N_CLK_c_4_p N_4_c_25_n 2.75361e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2125
cc_8 CLK N_4_c_26_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_4_p N_4_c_27_n 5.03453e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_10_p N_4_c_28_n 8.76278e-19 $X=0.081 $Y=0.1305 $X2=0.145 $Y2=0.135
cc_11 N_CLK_c_4_p N_4_c_29_n 3.53816e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.164
cc_12 N_CLK_c_4_p N_4_c_30_n 6.15177e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.172
cc_13 N_CLK_c_4_p N_4_c_31_n 0.00138527f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.189
cc_14 N_CLK_c_4_p N_4_c_32_n 9.65218e-19 $X=0.081 $Y=0.135 $X2=0.159 $Y2=0.189
cc_15 N_CLK_c_4_p N_4_c_33_n 0.00167589f $X=0.081 $Y=0.135 $X2=0.229 $Y2=0.189
cc_16 CLK N_6_c_142_n 6.45949e-19 $X=0.082 $Y=0.119 $X2=0 $Y2=0
cc_17 N_CLK_c_4_p N_6_c_143_n 6.54444e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_18 CLK N_6_c_144_n 6.20748e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.234
cc_19 N_4_c_34_p N_D_M2_g 0.00341068f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.054
cc_20 N_4_c_34_p N_D_c_122_n 0.0010364f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 N_4_c_36_p N_D_c_123_n 2.29805e-19 $X=0.29 $Y=0.189 $X2=0.081 $Y2=0.135
cc_22 N_4_c_37_p N_D_c_123_n 0.00102387f $X=0.513 $Y=0.189 $X2=0.081 $Y2=0.135
cc_23 N_4_c_38_p N_D_c_123_n 0.00337064f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_4_c_34_p N_6_M3_g 0.00355599f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.054
cc_25 N_4_M4_g N_6_M3_g 0.00355599f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_26 N_4_c_34_p N_6_c_147_n 0.00103664f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_27 N_4_M7_g N_6_M8_g 0.00355599f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_28 N_4_c_43_p N_6_M8_g 0.00355599f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_29 N_4_c_44_p N_6_M8_g 0.00250257f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_30 N_4_c_44_p N_6_c_151_n 0.00180656f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_31 N_4_c_46_p N_6_c_152_n 0.00135022f $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_32 N_4_c_47_p N_6_c_142_n 0.0010851f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_33 N_4_c_36_p N_6_c_154_n 4.24027e-19 $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_34 N_4_c_32_n N_6_c_143_n 0.00285029f $X=0.159 $Y=0.189 $X2=0 $Y2=0
cc_35 N_4_c_33_n N_6_c_143_n 6.46981e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_36 N_4_c_46_p N_6_c_143_n 2.904e-19 $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_37 N_4_c_33_n N_6_c_158_n 4.24027e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_38 N_4_c_47_p N_6_c_159_n 0.00351854f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_39 N_4_c_36_p N_6_c_159_n 0.00102595f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_40 N_4_c_44_p N_6_c_161_n 6.40799e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_41 N_4_c_44_p N_6_c_162_n 0.00187197f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_42 N_4_c_29_n N_6_c_162_n 3.52457e-19 $X=0.189 $Y=0.164 $X2=0 $Y2=0
cc_43 N_4_c_58_p N_6_c_162_n 2.46239e-19 $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_44 N_4_c_36_p N_6_c_162_n 0.0253778f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_45 N_4_c_38_p N_6_c_162_n 0.00115493f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_61_p N_6_c_162_n 2.81476e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_47 N_4_c_37_p N_6_c_168_n 2.98936e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_48 N_4_c_38_p N_6_c_168_n 0.00170246f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_49 N_4_c_44_p N_6_c_170_n 0.00124003f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_50 N_4_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_51 N_4_M7_g N_7_M5_g 2.13359e-19 $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_52 N_4_c_44_p N_7_M5_g 0.00205997f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_53 N_4_c_61_p N_7_M5_g 3.15189e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_54 N_4_c_44_p N_7_c_216_n 5.49754e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_55 N_4_c_44_p N_7_c_217_n 2.12581e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.1305
cc_56 N_4_c_44_p N_7_M21_s 2.50995e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_57 N_4_M7_g N_7_c_219_n 0.00200065f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_58 N_4_c_44_p N_7_c_219_n 0.00322783f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_59 N_4_M7_g N_7_c_221_n 3.04073e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_60 N_4_M7_g N_7_c_222_n 2.22997e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_61 N_4_c_61_p N_7_c_223_n 5.74745e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_62 N_4_c_77_p N_7_c_224_n 0.00193027f $X=0.621 $Y=0.178 $X2=0 $Y2=0
cc_63 N_4_c_44_p N_7_c_224_n 0.00189849f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_64 N_4_M7_g N_7_c_226_n 3.8308e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_65 N_4_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_66 N_4_M7_g N_8_M6_g 0.00341068f $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_67 N_4_c_44_p N_8_M6_g 0.00302156f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_68 N_4_c_37_p N_8_c_260_n 3.15319e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_69 N_4_c_38_p N_8_c_260_n 0.00136448f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_70 N_4_c_37_p N_8_c_262_n 0.00161272f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_71 N_4_M4_g N_8_c_263_n 3.80535e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_72 N_4_M4_g N_8_c_264_n 2.08362e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_73 N_4_M4_g N_8_c_265_n 2.27303e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_74 N_4_c_89_p N_8_c_266_n 4.73369e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_75 N_4_c_61_p N_8_c_266_n 0.00174159f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_76 N_4_c_89_p N_8_c_268_n 0.0017128f $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_77 N_4_c_44_p N_8_c_268_n 5.88593e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_78 N_4_c_37_p N_8_c_268_n 0.00102123f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_79 N_4_c_94_p N_8_c_268_n 3.42482e-19 $X=0.351 $Y=0.178 $X2=0 $Y2=0
cc_80 N_4_c_44_p N_8_c_272_n 8.16411e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_81 N_4_c_44_p N_8_c_273_n 3.32592e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_82 N_4_c_61_p N_8_c_273_n 8.9822e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_83 N_4_c_44_p N_8_c_275_n 5.02733e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_84 N_4_c_43_p N_9_M9_g 0.00341068f $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_85 N_4_c_43_p N_10_M10_g 2.13359e-19 $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_86 N_4_c_44_p N_10_c_337_n 8.27829e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_87 N_4_c_44_p N_10_M22_s 3.37661e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_88 N_4_c_44_p N_10_c_339_n 0.00145657f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_89 N_4_c_43_p N_10_c_340_n 2.71526e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_90 N_4_c_43_p N_10_c_341_n 2.11119e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_91 N_4_c_43_p N_10_c_342_n 2.58771e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_92 N_4_c_43_p N_10_c_343_n 0.00229157f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_93 N_4_c_44_p N_10_c_343_n 7.89371e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_94 N_4_c_43_p N_10_c_345_n 4.55487e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_95 N_4_c_44_p N_10_c_346_n 4.45535e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_96 N_4_c_43_p N_10_c_347_n 5.68093e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_97 N_4_c_44_p N_10_c_347_n 2.2968e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_98 N_4_c_34_p N_12_c_420_n 0.00526068f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_99 N_4_c_44_p N_13_M19_s 2.36286e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.216
cc_100 N_4_M4_g N_13_c_427_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_101 N_4_c_89_p N_13_c_427_n 5.41258e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_102 N_4_c_44_p N_13_c_427_n 0.00230928f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_103 N_4_c_37_p N_13_c_427_n 7.09553e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_104 N_4_c_43_p N_14_c_436_n 0.00198387f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_105 N_4_c_44_p N_14_c_436_n 4.51352e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_106 N_D_M2_g N_6_M3_g 2.82885e-19 $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_107 D N_6_c_172_n 0.00115224f $X=0.298 $Y=0.082 $X2=0.729 $Y2=0.178
cc_108 N_D_c_123_n N_6_c_154_n 0.00115224f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_109 N_D_c_123_n N_6_c_174_n 0.00115224f $X=0.297 $Y=0.135 $X2=0.725 $Y2=0.178
cc_110 N_D_c_123_n N_6_c_159_n 0.00124565f $X=0.297 $Y=0.135 $X2=0.729 $Y2=0.178
cc_111 D N_6_c_162_n 2.27807e-19 $X=0.298 $Y=0.082 $X2=0.056 $Y2=0.216
cc_112 N_D_c_123_n N_6_c_162_n 9.62099e-19 $X=0.297 $Y=0.135 $X2=0.056 $Y2=0.216
cc_113 N_D_c_133_p N_6_c_168_n 4.3159e-19 $X=0.297 $Y=0.126 $X2=0.018 $Y2=0.18
cc_114 D N_6_c_144_n 0.00115224f $X=0.298 $Y=0.082 $X2=0.054 $Y2=0.234
cc_115 N_D_c_133_p N_6_c_180_n 0.00115224f $X=0.297 $Y=0.126 $X2=0.054 $Y2=0.234
cc_116 N_D_c_123_n N_6_c_181_n 0.00115224f $X=0.297 $Y=0.135 $X2=0.047 $Y2=0.234
cc_117 N_D_c_123_n N_8_c_260_n 3.88702e-19 $X=0.297 $Y=0.135 $X2=0.621
+ $Y2=0.0405
cc_118 N_D_c_123_n N_8_c_262_n 8.77202e-19 $X=0.297 $Y=0.135 $X2=0.729
+ $Y2=0.2295
cc_119 D N_8_c_278_n 2.04306e-19 $X=0.298 $Y=0.082 $X2=0.018 $Y2=0.198
cc_120 D N_12_c_420_n 0.00430488f $X=0.298 $Y=0.082 $X2=0.351 $Y2=0.135
cc_121 N_D_c_123_n N_16_M17_s 3.05674e-19 $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_122 N_6_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_123 N_6_c_183_p N_7_c_228_n 2.96121e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_124 N_6_c_161_n N_7_c_229_n 2.61213e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_125 N_6_c_183_p N_7_c_229_n 2.61213e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_126 N_6_c_170_n N_7_c_221_n 0.00327797f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_127 N_6_c_161_n N_7_c_222_n 0.00115177f $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_128 N_6_c_161_n N_7_c_233_n 2.96121e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_129 N_6_M8_g N_8_M6_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_130 N_6_c_151_n N_8_c_280_n 4.12331e-19 $X=0.675 $Y=0.135 $X2=0.081 $Y2=0.135
cc_131 N_6_c_183_p N_8_c_280_n 2.64012e-19 $X=0.601 $Y=0.153 $X2=0.081 $Y2=0.135
cc_132 N_6_c_168_n N_8_c_260_n 2.25088e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_133 N_6_M3_g N_8_c_283_n 3.49806e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_134 N_6_c_168_n N_8_c_283_n 3.83282e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_135 N_6_c_168_n N_8_c_285_n 9.70699e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_136 N_6_c_168_n N_8_c_286_n 9.70699e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_137 N_6_c_162_n N_8_c_265_n 0.00118282f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_138 N_6_c_168_n N_8_c_265_n 0.00106411f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_139 N_6_c_162_n N_8_c_272_n 0.00138951f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_140 N_6_c_183_p N_8_c_275_n 0.00138951f $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_141 N_6_c_162_n N_8_c_291_n 2.54113e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_142 N_6_c_162_n N_8_c_278_n 3.92135e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_143 N_6_M8_g N_9_M9_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_144 N_6_c_161_n N_10_c_337_n 2.24654e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_145 N_6_c_161_n N_10_c_350_n 5.06919e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_146 N_6_M8_g N_10_c_351_n 3.43727e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_147 N_6_c_170_n N_10_c_351_n 5.96743e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_148 N_6_c_161_n N_10_c_353_n 2.34004e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_149 N_6_c_170_n N_10_c_341_n 0.00329725f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_150 N_6_c_161_n N_10_c_355_n 2.83245e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_151 N_6_c_162_n N_12_c_420_n 8.35084e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_152 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_153 N_7_c_235_p N_8_M6_g 3.91159e-19 $X=0.581 $Y=0.09 $X2=0.135 $Y2=0.054
cc_154 N_7_c_236_p N_8_c_263_n 2.10569e-19 $X=0.594 $Y=0.054 $X2=0.464 $Y2=0.178
cc_155 N_7_c_237_p N_8_c_264_n 3.19692e-19 $X=0.513 $Y=0.09 $X2=0 $Y2=0
cc_156 N_7_c_235_p N_8_c_264_n 0.00107929f $X=0.581 $Y=0.09 $X2=0 $Y2=0
cc_157 N_7_c_221_n N_8_c_298_n 2.4251e-19 $X=0.621 $Y=0.122 $X2=0 $Y2=0
cc_158 N_7_c_240_p N_8_c_299_n 9.84729e-19 $X=0.621 $Y=0.14 $X2=0.056 $Y2=0.054
cc_159 N_7_c_235_p N_8_c_300_n 0.00507595f $X=0.581 $Y=0.09 $X2=0 $Y2=0
cc_160 N_7_M5_g N_8_c_273_n 3.12986e-19 $X=0.513 $Y=0.0405 $X2=0.071 $Y2=0.216
cc_161 N_7_c_237_p N_8_c_291_n 5.2508e-19 $X=0.513 $Y=0.09 $X2=0.018 $Y2=0.18
cc_162 N_7_c_236_p N_8_c_303_n 2.10569e-19 $X=0.594 $Y=0.054 $X2=0.018 $Y2=0.125
cc_163 N_7_c_216_n N_10_c_337_n 0.00328169f $X=0.594 $Y=0.0405 $X2=0 $Y2=0
cc_164 N_7_c_236_p N_10_c_337_n 3.00222e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_165 N_7_c_226_n N_10_c_337_n 2.70684e-19 $X=0.621 $Y=0.09 $X2=0 $Y2=0
cc_166 N_7_c_219_n N_10_c_339_n 0.00222825f $X=0.65 $Y=0.2295 $X2=0.725
+ $Y2=0.178
cc_167 N_7_c_216_n N_10_c_350_n 3.50513e-19 $X=0.594 $Y=0.0405 $X2=0.056
+ $Y2=0.054
cc_168 N_7_c_236_p N_10_c_350_n 5.0339e-19 $X=0.594 $Y=0.054 $X2=0.056 $Y2=0.054
cc_169 N_7_c_236_p N_10_c_362_n 2.21141e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_170 N_7_c_226_n N_10_c_340_n 4.36168e-19 $X=0.621 $Y=0.09 $X2=0.056 $Y2=0.216
cc_171 N_7_c_253_p N_10_c_343_n 4.36168e-19 $X=0.621 $Y=0.214 $X2=0.018 $Y2=0.07
cc_172 N_7_c_219_n N_10_c_346_n 3.64454e-19 $X=0.65 $Y=0.2295 $X2=0.135
+ $Y2=0.135
cc_173 N_7_c_255_p N_10_c_346_n 4.86017e-19 $X=0.612 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_174 N_7_c_224_n N_10_c_347_n 4.36168e-19 $X=0.621 $Y=0.203 $X2=0.148
+ $Y2=0.135
cc_175 N_8_c_260_n N_12_c_420_n 0.00119636f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.135
cc_176 N_8_c_291_n N_12_c_420_n 0.00390673f $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_177 N_8_c_278_n N_12_c_420_n 4.41747e-19 $X=0.45 $Y=0.036 $X2=0.351 $Y2=0.135
cc_178 N_8_c_260_n N_13_c_427_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.135
cc_179 N_8_c_308_p N_13_c_427_n 0.00209454f $X=0.45 $Y=0.234 $X2=0.351 $Y2=0.135
cc_180 N_8_c_309_p N_13_c_427_n 0.0013184f $X=0.434 $Y=0.234 $X2=0.351 $Y2=0.135
cc_181 N_8_c_310_p N_13_c_427_n 0.00116187f $X=0.459 $Y=0.225 $X2=0.351
+ $Y2=0.135
cc_182 N_8_c_291_n N_13_c_427_n 5.72158e-19 $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_183 N_9_M9_g N_10_M10_g 0.00268443f $X=0.783 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_184 N_9_c_315_p N_10_M10_g 3.74489e-19 $X=0.846 $Y=0.036 $X2=0.135 $Y2=0.054
cc_185 N_9_c_316_p N_10_c_370_n 0.00141609f $X=0.792 $Y=0.036 $X2=0.725
+ $Y2=0.178
cc_186 N_9_c_317_p N_10_c_362_n 0.00141609f $X=0.783 $Y=0.105 $X2=0 $Y2=0
cc_187 N_9_c_318_p N_10_c_340_n 3.34766e-19 $X=0.783 $Y=0.1055 $X2=0.056
+ $Y2=0.216
cc_188 N_9_c_317_p N_10_c_340_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.056
+ $Y2=0.216
cc_189 N_9_c_320_p N_10_c_343_n 2.41112e-19 $X=0.945 $Y=0.225 $X2=0.018 $Y2=0.07
cc_190 N_9_c_321_p N_10_c_375_n 2.65946e-19 $X=0.828 $Y=0.036 $X2=0.018
+ $Y2=0.125
cc_191 N_9_M9_g N_10_c_376_n 6.3699e-19 $X=0.783 $Y=0.0405 $X2=0.018 $Y2=0.2
cc_192 N_9_c_317_p N_10_c_376_n 9.10342e-19 $X=0.783 $Y=0.105 $X2=0.018 $Y2=0.2
cc_193 N_9_c_315_p N_10_c_378_n 4.40983e-19 $X=0.846 $Y=0.036 $X2=0.054
+ $Y2=0.036
cc_194 N_9_c_325_p N_10_c_379_n 5.181e-19 $X=0.882 $Y=0.036 $X2=0.054 $Y2=0.234
cc_195 N_9_c_326_p N_10_c_380_n 0.00149072f $X=0.9 $Y=0.234 $X2=0.054 $Y2=0.234
cc_196 N_9_c_327_p N_10_c_381_n 4.52584e-19 $X=0.9 $Y=0.036 $X2=0.189 $Y2=0.172
cc_197 N_9_c_328_p N_10_c_381_n 0.00299476f $X=0.945 $Y=0.167 $X2=0.189
+ $Y2=0.172
cc_198 N_9_c_329_p N_10_c_355_n 2.40515e-19 $X=0.936 $Y=0.036 $X2=0.033
+ $Y2=0.189
cc_199 N_9_c_330_p N_10_c_355_n 7.44774e-19 $X=0.918 $Y=0.234 $X2=0.033
+ $Y2=0.189
cc_200 N_9_c_328_p N_10_c_355_n 8.84468e-19 $X=0.945 $Y=0.167 $X2=0.033
+ $Y2=0.189
cc_201 N_9_c_332_p N_10_c_386_n 0.00323217f $X=0.945 $Y=0.117 $X2=0.229
+ $Y2=0.189
cc_202 N_9_c_329_p N_QN_c_405_n 4.8595e-19 $X=0.936 $Y=0.036 $X2=0 $Y2=0
cc_203 N_9_c_334_p N_QN_c_406_n 4.61952e-19 $X=0.936 $Y=0.234 $X2=0.729
+ $Y2=0.2295
cc_204 N_9_c_316_p N_14_c_436_n 7.33799e-19 $X=0.792 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_205 N_10_c_387_p N_QN_M12_d 3.7444e-19 $X=1.107 $Y=0.136 $X2=0.135 $Y2=0.054
cc_206 N_10_c_387_p N_QN_M26_d 3.85232e-19 $X=1.107 $Y=0.136 $X2=0 $Y2=0
cc_207 N_10_c_387_p N_QN_c_409_n 8.43851e-19 $X=1.107 $Y=0.136 $X2=0.459
+ $Y2=0.0405
cc_208 N_10_M12_g N_QN_c_410_n 4.61823e-19 $X=1.053 $Y=0.0675 $X2=0.621
+ $Y2=0.0405
cc_209 N_10_M13_g N_QN_c_410_n 4.61823e-19 $X=1.107 $Y=0.0675 $X2=0.621
+ $Y2=0.0405
cc_210 N_10_c_387_p N_QN_c_405_n 0.00133402f $X=1.107 $Y=0.136 $X2=0 $Y2=0
cc_211 N_10_c_387_p N_QN_c_413_n 7.60428e-19 $X=1.107 $Y=0.136 $X2=0.621
+ $Y2=0.178
cc_212 N_10_c_386_n N_QN_c_413_n 6.32739e-19 $X=0.999 $Y=0.136 $X2=0.621
+ $Y2=0.178
cc_213 N_10_M12_g N_QN_c_406_n 4.56718e-19 $X=1.053 $Y=0.0675 $X2=0.729
+ $Y2=0.2295
cc_214 N_10_M13_g N_QN_c_406_n 4.56718e-19 $X=1.107 $Y=0.0675 $X2=0.729
+ $Y2=0.2295
cc_215 N_10_c_387_p N_QN_c_406_n 0.00135857f $X=1.107 $Y=0.136 $X2=0.729
+ $Y2=0.2295
cc_216 N_10_c_387_p QN 3.65358e-19 $X=1.107 $Y=0.136 $X2=0.725 $Y2=0.178
cc_217 N_10_c_386_n N_QN_c_419_n 4.8083e-19 $X=0.999 $Y=0.136 $X2=0 $Y2=0
cc_218 N_10_c_337_n N_14_c_436_n 0.00182708f $X=0.648 $Y=0.0405 $X2=0.351
+ $Y2=0.135
cc_219 N_10_c_370_n N_14_c_436_n 0.00205226f $X=0.72 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_220 N_10_c_402_p N_14_c_436_n 0.0013184f $X=0.704 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_221 N_10_c_362_n N_14_c_436_n 0.00103589f $X=0.729 $Y=0.081 $X2=0.351
+ $Y2=0.135
cc_222 N_10_c_345_n N_14_c_436_n 4.02739e-19 $X=0.774 $Y=0.162 $X2=0.351
+ $Y2=0.135

* END of "./DFFLQNx3_ASAP7_75t_SRAM.pex.sp.DFFLQNX3_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DFFLQx4_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:26:46 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DFFLQx4_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DFFLQx4_ASAP7_75t_SRAM.pex.sp.pex"
* File: DFFLQx4_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:26:46 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DFFLQX4_ASAP7_75T_SRAM%CLK 2 5 7 12 14 17 VSS
c18 17 VSS 1.44512e-20 $X=0.081 $Y=0.1305
c19 14 VSS 0.00697951f $X=0.081 $Y=0.135
c20 12 VSS 0.00694053f $X=0.082 $Y=0.119
c21 5 VSS 0.00190705f $X=0.081 $Y=0.135
c22 2 VSS 0.0629f $X=0.081 $Y=0.054
r23 16 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r24 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r25 12 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.126
r26 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%4 2 5 7 10 13 16 22 25 28 31 36 43 47 50 52 58 59
+ 60 64 67 74 79 84 88 89 92 96 99 100 101 103 111 124 132 148 VSS
c102 148 VSS 4.19842e-19 $X=0.18 $Y=0.189
c103 147 VSS 1.53928e-19 $X=0.189 $Y=0.189
c104 141 VSS 7.0154e-20 $X=0.03 $Y=0.189
c105 140 VSS 5.9624e-19 $X=0.027 $Y=0.189
c106 124 VSS 6.81413e-19 $X=0.513 $Y=0.18
c107 111 VSS 4.0846e-19 $X=0.351 $Y=0.135
c108 103 VSS 0.00656068f $X=0.513 $Y=0.189
c109 101 VSS 0.0025144f $X=0.29 $Y=0.189
c110 100 VSS 0.00601911f $X=0.229 $Y=0.189
c111 99 VSS 7.60117e-19 $X=0.351 $Y=0.189
c112 96 VSS 4.13928e-19 $X=0.159 $Y=0.189
c113 92 VSS 4.95517e-19 $X=0.033 $Y=0.189
c114 89 VSS 7.37649e-20 $X=0.189 $Y=0.172
c115 88 VSS 5.63427e-19 $X=0.189 $Y=0.164
c116 87 VSS 1.04741e-19 $X=0.189 $Y=0.18
c117 85 VSS 9.32714e-20 $X=0.148 $Y=0.135
c118 84 VSS 9.68697e-19 $X=0.145 $Y=0.135
c119 79 VSS 0.00149077f $X=0.18 $Y=0.135
c120 77 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c121 76 VSS 0.00169428f $X=0.047 $Y=0.234
c122 74 VSS 0.00250477f $X=0.054 $Y=0.234
c123 72 VSS 0.00306385f $X=0.027 $Y=0.234
c124 70 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c125 69 VSS 0.00205521f $X=0.047 $Y=0.036
c126 67 VSS 0.00250477f $X=0.054 $Y=0.036
c127 65 VSS 0.00305101f $X=0.027 $Y=0.036
c128 64 VSS 4.99402e-19 $X=0.018 $Y=0.2125
c129 63 VSS 1.14289e-19 $X=0.018 $Y=0.2
c130 62 VSS 4.86272e-19 $X=0.018 $Y=0.225
c131 60 VSS 0.00271341f $X=0.018 $Y=0.125
c132 59 VSS 9.57865e-19 $X=0.018 $Y=0.07
c133 58 VSS 0.00235012f $X=0.018 $Y=0.18
c134 55 VSS 0.00586466f $X=0.056 $Y=0.216
c135 52 VSS 2.98509e-19 $X=0.071 $Y=0.216
c136 50 VSS 0.00549524f $X=0.056 $Y=0.054
c137 47 VSS 2.98509e-19 $X=0.071 $Y=0.054
c138 43 VSS 0.0592182f $X=0.725 $Y=0.178
c139 36 VSS 0.0013168f $X=0.464 $Y=0.178
c140 28 VSS 0.061209f $X=0.729 $Y=0.178
c141 25 VSS 1.44609e-19 $X=0.621 $Y=0.178
c142 22 VSS 0.0600171f $X=0.621 $Y=0.0405
c143 16 VSS 0.0601675f $X=0.459 $Y=0.0405
c144 10 VSS 0.0609009f $X=0.351 $Y=0.135
c145 5 VSS 0.00210427f $X=0.135 $Y=0.135
c146 2 VSS 0.0623856f $X=0.135 $Y=0.054
r147 148 149 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.189 $X2=0.1845 $Y2=0.189
r148 147 149 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.189 $X2=0.1845 $Y2=0.189
r149 140 141 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.03 $Y2=0.189
r150 137 140 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.027 $Y2=0.189
r151 131 132 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.351 $Y=0.167 $X2=0.351 $Y2=0.178
r152 123 124 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r153 111 131 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.167
r154 103 124 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r155 100 101 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.189 $X2=0.29 $Y2=0.189
r156 99 132 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.178
r157 98 103 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.513 $Y2=0.189
r158 98 101 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.29 $Y2=0.189
r159 98 99 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.189 $X2=0.351
+ $Y2=0.189
r160 96 148 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.159
+ $Y=0.189 $X2=0.18 $Y2=0.189
r161 95 100 4.75309 $w=1.8e-08 $l=7e-08 $layer=M2 $thickness=3.6e-08 $X=0.159
+ $Y=0.189 $X2=0.229 $Y2=0.189
r162 95 96 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.159 $Y=0.189 $X2=0.159
+ $Y2=0.189
r163 92 141 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.03 $Y2=0.189
r164 91 95 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.159 $Y2=0.189
r165 91 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.189 $X2=0.033
+ $Y2=0.189
r166 88 89 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.172
r167 87 147 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.189
r168 87 89 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.172
r169 86 88 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.164
r170 84 85 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.145
+ $Y=0.135 $X2=0.148 $Y2=0.135
r171 81 84 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.145 $Y2=0.135
r172 79 86 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r173 79 85 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.148 $Y2=0.135
r174 76 77 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r175 74 77 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r176 72 76 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r177 69 70 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r178 67 70 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r179 65 69 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r180 63 64 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r181 62 72 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r182 62 64 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r183 61 137 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.189
r184 61 63 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.2
r185 59 60 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.125
r186 58 137 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.189
r187 58 60 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.125
r188 57 65 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r189 57 59 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r190 55 74 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r191 52 55 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r192 50 67 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r193 47 50 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r194 36 123 39.0385 $w=2.6e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.178 $X2=0.513 $Y2=0.178
r195 28 43 3.07692 $w=2.6e-08 $l=4e-09 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.178 $X2=0.725 $Y2=0.178
r196 28 31 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.178 $X2=0.729 $Y2=0.2295
r197 25 43 82.8571 $w=2.6e-08 $l=1.04e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.725 $Y2=0.178
r198 25 123 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.621 $Y=0.178 $X2=0.513 $Y2=0.178
r199 22 25 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0405 $X2=0.621 $Y2=0.178
r200 19 36 3.84615 $w=2.6e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.178 $X2=0.464 $Y2=0.178
r201 16 19 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.178
r202 10 111 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135
+ $X2=0.351 $Y2=0.135
r203 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r204 5 81 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r205 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r206 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%D 2 5 7 12 14 17 VSS
c21 17 VSS 2.32756e-19 $X=0.297 $Y=0.126
c22 14 VSS 0.0072156f $X=0.297 $Y=0.135
c23 12 VSS 0.00703905f $X=0.298 $Y=0.082
c24 5 VSS 0.00213729f $X=0.297 $Y=0.135
c25 2 VSS 0.061556f $X=0.297 $Y=0.0675
r26 16 17 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.126
r27 14 17 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.126
r28 12 16 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.082 $X2=0.297 $Y2=0.106
r29 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r30 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r31 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%6 2 5 7 10 13 15 17 22 25 27 32 34 39 40 42 45 51
+ 53 54 58 63 73 74 76 VSS
c72 76 VSS 7.88952e-19 $X=0.243 $Y=0.2115
c73 74 VSS 8.75359e-19 $X=0.243 $Y=0.126
c74 73 VSS 0.00233088f $X=0.243 $Y=0.106
c75 63 VSS 0.00103743f $X=0.675 $Y=0.135
c76 58 VSS 9.14968e-19 $X=0.405 $Y=0.135
c77 54 VSS 0.00260015f $X=0.601 $Y=0.153
c78 53 VSS 0.00774972f $X=0.527 $Y=0.153
c79 51 VSS 0.00402804f $X=0.675 $Y=0.153
c80 45 VSS 0.00167713f $X=0.243 $Y=0.153
c81 42 VSS 5.5218e-19 $X=0.243 $Y=0.225
c82 40 VSS 0.00181981f $X=0.216 $Y=0.234
c83 39 VSS 0.00525711f $X=0.198 $Y=0.234
c84 34 VSS 0.00482554f $X=0.234 $Y=0.234
c85 33 VSS 0.00200074f $X=0.216 $Y=0.036
c86 32 VSS 0.00545403f $X=0.198 $Y=0.036
c87 27 VSS 0.00500597f $X=0.234 $Y=0.036
c88 25 VSS 0.00714358f $X=0.16 $Y=0.216
c89 20 VSS 0.00667633f $X=0.16 $Y=0.054
c90 13 VSS 0.00207734f $X=0.675 $Y=0.135
c91 10 VSS 0.0585656f $X=0.675 $Y=0.0405
c92 5 VSS 0.00164533f $X=0.405 $Y=0.135
c93 2 VSS 0.058827f $X=0.405 $Y=0.0675
r94 75 76 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.198 $X2=0.243 $Y2=0.2115
r95 73 74 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.106 $X2=0.243 $Y2=0.126
r96 53 54 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.601 $Y2=0.153
r97 51 54 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.675
+ $Y=0.153 $X2=0.601 $Y2=0.153
r98 51 63 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.675 $Y=0.153 $X2=0.675
+ $Y2=0.153
r99 48 53 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.527 $Y2=0.153
r100 48 58 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r101 45 75 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.198
r102 45 74 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.126
r103 44 48 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.405 $Y2=0.153
r104 44 45 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.153 $X2=0.243
+ $Y2=0.153
r105 42 76 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.2115
r106 41 73 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.106
r107 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.216 $Y2=0.234
r108 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.198 $Y2=0.234
r109 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r110 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r111 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.216 $Y2=0.036
r112 29 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r113 27 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r114 27 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r115 25 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r116 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r117 20 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r118 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r119 13 63 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.135 $X2=0.675
+ $Y2=0.135
r120 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2295
r121 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.135
r122 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r123 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2295
r124 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%7 2 5 7 9 10 13 14 17 19 22 29 30 31 33 40 47 48
+ 49 50 51 52 54 55 VSS
c46 56 VSS 3.57489e-19 $X=0.612 $Y=0.09
c47 55 VSS 1.84136e-19 $X=0.603 $Y=0.09
c48 54 VSS 5.96246e-19 $X=0.621 $Y=0.09
c49 52 VSS 4.34097e-19 $X=0.621 $Y=0.214
c50 51 VSS 4.90038e-19 $X=0.621 $Y=0.203
c51 50 VSS 1.59683e-19 $X=0.621 $Y=0.167
c52 49 VSS 2.89857e-19 $X=0.621 $Y=0.165
c53 48 VSS 2.84103e-19 $X=0.621 $Y=0.14
c54 47 VSS 3.66508e-19 $X=0.621 $Y=0.122
c55 46 VSS 3.21714e-19 $X=0.621 $Y=0.225
c56 40 VSS 0.00154565f $X=0.594 $Y=0.054
c57 33 VSS 0.00268134f $X=0.594 $Y=0.234
c58 31 VSS 0.00427376f $X=0.612 $Y=0.234
c59 30 VSS 1.96699e-19 $X=0.583 $Y=0.09
c60 29 VSS 0.00266746f $X=0.581 $Y=0.09
c61 24 VSS 5.17345e-20 $X=0.585 $Y=0.09
c62 22 VSS 0.0185835f $X=0.65 $Y=0.2295
c63 19 VSS 3.14771e-19 $X=0.665 $Y=0.2295
c64 17 VSS 2.5391e-19 $X=0.592 $Y=0.2295
c65 13 VSS 0.00441429f $X=0.594 $Y=0.0405
c66 9 VSS 6.29543e-19 $X=0.611 $Y=0.0405
c67 5 VSS 0.00249952f $X=0.513 $Y=0.09
c68 2 VSS 0.0583002f $X=0.513 $Y=0.0405
r69 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.603
+ $Y=0.09 $X2=0.612 $Y2=0.09
r70 54 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.612 $Y2=0.09
r71 53 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.09 $X2=0.603 $Y2=0.09
r72 51 52 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.214
r73 50 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.203
r74 49 50 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.167
r75 48 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r76 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r77 46 52 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.214
r78 45 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.09
r79 45 47 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.099 $X2=0.621 $Y2=0.122
r80 38 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.09
r81 38 40 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.081 $X2=0.594 $Y2=0.054
r82 31 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r83 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r84 29 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.581
+ $Y=0.09 $X2=0.583 $Y2=0.09
r85 26 29 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.09 $X2=0.581 $Y2=0.09
r86 24 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.594 $Y2=0.09
r87 24 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.09 $X2=0.583 $Y2=0.09
r88 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2295 $X2=0.65 $Y2=0.2295
r89 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.592
+ $Y=0.2295 $X2=0.65 $Y2=0.2295
r90 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r91 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r92 13 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.054 $X2=0.594
+ $Y2=0.054
r93 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.594 $Y2=0.0405
r94 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0405 $X2=0.594 $Y2=0.0405
r95 5 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.09 $X2=0.513
+ $Y2=0.09
r96 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.09 $X2=0.513 $Y2=0.2295
r97 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.09
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%8 2 5 7 9 14 17 21 22 25 30 31 33 35 36 37 38 39
+ 41 42 43 44 48 50 51 52 53 58 60 61 VSS
c57 64 VSS 2.84134e-19 $X=0.459 $Y=0.131
c58 61 VSS 0.0033683f $X=0.45 $Y=0.036
c59 60 VSS 0.00242977f $X=0.459 $Y=0.036
c60 58 VSS 0.00400835f $X=0.432 $Y=0.036
c61 53 VSS 4.23511e-19 $X=0.5445 $Y=0.131
c62 52 VSS 3.49205e-20 $X=0.522 $Y=0.131
c63 51 VSS 2.0008e-19 $X=0.504 $Y=0.131
c64 50 VSS 0.00133205f $X=0.496 $Y=0.131
c65 48 VSS 5.65722e-19 $X=0.567 $Y=0.131
c66 45 VSS 4.52499e-19 $X=0.459 $Y=0.214
c67 44 VSS 2.01779e-19 $X=0.459 $Y=0.203
c68 43 VSS 6.09344e-21 $X=0.459 $Y=0.167
c69 42 VSS 1.59896e-19 $X=0.459 $Y=0.165
c70 41 VSS 3.22081e-19 $X=0.459 $Y=0.225
c71 39 VSS 2.48018e-19 $X=0.459 $Y=0.114
c72 38 VSS 2.28952e-19 $X=0.459 $Y=0.106
c73 37 VSS 9.45429e-20 $X=0.459 $Y=0.099
c74 36 VSS 8.12259e-19 $X=0.459 $Y=0.081
c75 35 VSS 2.08428e-19 $X=0.459 $Y=0.122
c76 33 VSS 0.00142907f $X=0.434 $Y=0.234
c77 32 VSS 3.74355e-19 $X=0.418 $Y=0.234
c78 31 VSS 0.00146362f $X=0.414 $Y=0.234
c79 30 VSS 0.00368961f $X=0.396 $Y=0.234
c80 25 VSS 0.00389542f $X=0.45 $Y=0.234
c81 24 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c82 21 VSS 0.00423578f $X=0.378 $Y=0.2025
c83 16 VSS 5.70081e-19 $X=0.432 $Y=0.0405
c84 5 VSS 0.00175503f $X=0.567 $Y=0.1305
c85 2 VSS 0.0591962f $X=0.567 $Y=0.0405
r86 61 62 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r87 60 62 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r88 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r89 57 58 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r90 52 53 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r91 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r92 50 51 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.496
+ $Y=0.131 $X2=0.504 $Y2=0.131
r93 48 53 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.131 $X2=0.5445 $Y2=0.131
r94 46 64 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r95 46 50 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.496 $Y2=0.131
r96 44 45 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.203 $X2=0.459 $Y2=0.214
r97 43 44 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.167 $X2=0.459 $Y2=0.203
r98 42 43 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.167
r99 41 45 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r100 40 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r101 40 42 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.165
r102 38 39 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.106 $X2=0.459 $Y2=0.114
r103 37 38 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.099 $X2=0.459 $Y2=0.106
r104 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.081 $X2=0.459 $Y2=0.099
r105 35 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r106 35 39 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.114
r107 34 60 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r108 34 36 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.081
r109 32 33 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.234 $X2=0.434 $Y2=0.234
r110 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.418 $Y2=0.234
r111 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r112 27 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r113 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r114 25 33 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.434 $Y2=0.234
r115 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r116 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r117 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r118 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r119 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r120 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r121 13 58 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r122 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r123 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r124 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r125 5 48 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.131 $X2=0.567
+ $Y2=0.131
r126 5 7 370.904 $w=2e-08 $l=9.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1305 $X2=0.567 $Y2=0.2295
r127 2 5 337.185 $w=2e-08 $l=9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.1305
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%9 2 5 7 9 14 21 25 26 30 31 32 33 34 39 40 42 44
+ 45 VSS
c24 46 VSS 2.95823e-19 $X=0.945 $Y=0.171
c25 45 VSS 9.82877e-19 $X=0.945 $Y=0.167
c26 44 VSS 3.06877e-19 $X=0.945 $Y=0.122
c27 43 VSS 0.00344802f $X=0.945 $Y=0.117
c28 42 VSS 0.00284656f $X=0.945 $Y=0.225
c29 40 VSS 0.0018377f $X=0.918 $Y=0.234
c30 39 VSS 0.0056872f $X=0.9 $Y=0.234
c31 34 VSS 0.00462933f $X=0.936 $Y=0.234
c32 33 VSS 0.00189638f $X=0.9 $Y=0.036
c33 32 VSS 0.00352438f $X=0.882 $Y=0.036
c34 31 VSS 0.00146362f $X=0.846 $Y=0.036
c35 30 VSS 0.00478092f $X=0.828 $Y=0.036
c36 26 VSS 0.00226308f $X=0.792 $Y=0.036
c37 25 VSS 0.00657446f $X=0.936 $Y=0.036
c38 21 VSS 0.00135803f $X=0.783 $Y=0.105
c39 17 VSS 0.00535471f $X=0.862 $Y=0.2295
c40 12 VSS 0.00569943f $X=0.862 $Y=0.0405
c41 5 VSS 0.00257499f $X=0.783 $Y=0.1055
c42 2 VSS 0.0589361f $X=0.783 $Y=0.0405
r43 45 46 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.167 $X2=0.945 $Y2=0.171
r44 44 45 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.122 $X2=0.945 $Y2=0.167
r45 43 44 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.117 $X2=0.945 $Y2=0.122
r46 42 46 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.171
r47 41 43 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.117
r48 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.234 $X2=0.918 $Y2=0.234
r49 36 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.9 $Y2=0.234
r50 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r51 34 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.918 $Y2=0.234
r52 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r53 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.846 $Y2=0.036
r54 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r55 28 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.846 $Y2=0.036
r56 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.036 $X2=0.828 $Y2=0.036
r57 25 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r58 25 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.9 $Y2=0.036
r59 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.783 $Y=0.045 $X2=0.792 $Y2=0.036
r60 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.105
r61 17 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234 $X2=0.864
+ $Y2=0.234
r62 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2295 $X2=0.862 $Y2=0.2295
r63 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036 $X2=0.864
+ $Y2=0.036
r64 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.862 $Y2=0.0405
r65 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.105 $X2=0.783
+ $Y2=0.105
r66 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.1055 $X2=0.783 $Y2=0.2295
r67 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.1055
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%10 2 5 7 10 15 18 21 23 25 26 29 30 31 34 35 40
+ 41 43 45 46 47 48 49 51 52 54 55 58 65 66 74 77 81 84 92 VSS
c71 92 VSS 0.00121551f $X=0.999 $Y=0.136
c72 84 VSS 0.00773455f $X=0.999 $Y=0.153
c73 81 VSS 0.00168296f $X=0.891 $Y=0.153
c74 78 VSS 4.17512e-19 $X=0.837 $Y=0.162
c75 77 VSS 1.52743e-19 $X=0.729 $Y=0.162
c76 74 VSS 0.00371016f $X=0.72 $Y=0.234
c77 73 VSS 0.00254161f $X=0.729 $Y=0.234
c78 66 VSS 4.13886e-19 $X=0.866 $Y=0.162
c79 65 VSS 1.34754e-19 $X=0.85 $Y=0.162
c80 63 VSS 2.72392e-19 $X=0.882 $Y=0.162
c81 58 VSS 3.90416e-19 $X=0.837 $Y=0.135
c82 55 VSS 3.26354e-19 $X=0.792 $Y=0.162
c83 54 VSS 0.00200395f $X=0.774 $Y=0.162
c84 52 VSS 0.00182634f $X=0.828 $Y=0.162
c85 51 VSS 0.00130761f $X=0.729 $Y=0.225
c86 49 VSS 1.5228e-19 $X=0.729 $Y=0.136
c87 48 VSS 9.59255e-20 $X=0.729 $Y=0.119
c88 47 VSS 1.29374e-19 $X=0.729 $Y=0.099
c89 46 VSS 3.52175e-19 $X=0.729 $Y=0.081
c90 45 VSS 2.74133e-19 $X=0.729 $Y=0.153
c91 43 VSS 0.00166806f $X=0.704 $Y=0.036
c92 42 VSS 4.59162e-19 $X=0.688 $Y=0.036
c93 41 VSS 0.00146362f $X=0.684 $Y=0.036
c94 40 VSS 0.00370406f $X=0.666 $Y=0.036
c95 35 VSS 0.00402343f $X=0.72 $Y=0.036
c96 34 VSS 0.00352608f $X=0.702 $Y=0.2295
c97 30 VSS 5.63046e-19 $X=0.719 $Y=0.2295
c98 29 VSS 0.0329964f $X=0.648 $Y=0.0405
c99 25 VSS 5.63046e-19 $X=0.665 $Y=0.0405
c100 21 VSS 0.00425996f $X=1.053 $Y=0.136
c101 18 VSS 0.0584171f $X=1.053 $Y=0.0675
c102 10 VSS 0.0615046f $X=0.999 $Y=0.0675
c103 5 VSS 0.0018803f $X=0.837 $Y=0.135
c104 2 VSS 0.0618222f $X=0.837 $Y=0.0405
r105 84 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.999 $Y=0.153 $X2=0.999
+ $Y2=0.153
r106 80 84 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.999 $Y2=0.153
r107 80 81 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r108 74 75 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.234 $X2=0.7245 $Y2=0.234
r109 73 75 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.234 $X2=0.7245 $Y2=0.234
r110 70 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.234 $X2=0.72 $Y2=0.234
r111 65 66 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.85
+ $Y=0.162 $X2=0.866 $Y2=0.162
r112 64 78 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.837 $Y2=0.162
r113 64 65 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.162 $X2=0.85 $Y2=0.162
r114 63 81 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.891 $Y2=0.162
r115 63 66 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.162 $X2=0.866 $Y2=0.162
r116 56 78 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.162
r117 56 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=0.837 $Y2=0.135
r118 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.162 $X2=0.792 $Y2=0.162
r119 53 77 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.729 $Y2=0.162
r120 53 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.162 $X2=0.774 $Y2=0.162
r121 52 78 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.837 $Y2=0.162
r122 52 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.162 $X2=0.792 $Y2=0.162
r123 51 73 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.225 $X2=0.729 $Y2=0.234
r124 50 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.162
r125 50 51 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.171 $X2=0.729 $Y2=0.225
r126 48 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.119 $X2=0.729 $Y2=0.136
r127 47 48 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.099 $X2=0.729 $Y2=0.119
r128 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.081 $X2=0.729 $Y2=0.099
r129 45 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.162
r130 45 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.729 $Y2=0.136
r131 44 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.045 $X2=0.729 $Y2=0.081
r132 42 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.036 $X2=0.704 $Y2=0.036
r133 41 42 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.688 $Y2=0.036
r134 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.684 $Y2=0.036
r135 37 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.666 $Y2=0.036
r136 35 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.036 $X2=0.729 $Y2=0.045
r137 35 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.704 $Y2=0.036
r138 34 70 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.234
+ $X2=0.702 $Y2=0.234
r139 31 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2295 $X2=0.702 $Y2=0.2295
r140 30 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2295 $X2=0.702 $Y2=0.2295
r141 29 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r142 26 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0405 $X2=0.648 $Y2=0.0405
r143 25 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r144 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.136 $X2=1.053 $Y2=0.2025
r145 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.0675 $X2=1.053 $Y2=0.136
r146 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.999
+ $Y=0.136 $X2=1.053 $Y2=0.136
r147 13 92 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.136 $X2=0.999
+ $Y2=0.136
r148 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.136 $X2=0.999 $Y2=0.2025
r149 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.136
r150 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.135 $X2=0.837
+ $Y2=0.135
r151 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.2295
r152 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.0405 $X2=0.837 $Y2=0.135
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%11 2 7 10 15 18 23 26 29 31 33 34 38 39 42 43 46
+ 48 54 55 58 59 63 66 68 VSS
c43 68 VSS 3.78938e-19 $X=1.089 $Y=0.136
c44 66 VSS 4.82002e-21 $X=1.143 $Y=0.136
c45 65 VSS 7.16275e-19 $X=1.125 $Y=0.136
c46 63 VSS 1.52274e-19 $X=1.161 $Y=0.136
c47 60 VSS 0.00141149f $X=1.089 $Y=0.201
c48 59 VSS 8.53779e-19 $X=1.089 $Y=0.167
c49 58 VSS 6.05349e-19 $X=1.089 $Y=0.225
c50 56 VSS 0.00227099f $X=1.089 $Y=0.122
c51 55 VSS 7.78235e-19 $X=1.089 $Y=0.069
c52 54 VSS 3.06947e-19 $X=1.089 $Y=0.127
c53 48 VSS 0.0110409f $X=1.08 $Y=0.234
c54 46 VSS 0.00899572f $X=1.026 $Y=0.036
c55 43 VSS 0.0110409f $X=1.08 $Y=0.036
c56 42 VSS 0.00937164f $X=1.026 $Y=0.2025
c57 38 VSS 5.72268e-19 $X=1.043 $Y=0.2025
c58 33 VSS 5.72268e-19 $X=1.043 $Y=0.0675
c59 29 VSS 0.0143997f $X=1.269 $Y=0.136
c60 26 VSS 0.0615048f $X=1.269 $Y=0.0675
c61 18 VSS 0.0615873f $X=1.215 $Y=0.0675
c62 10 VSS 0.061355f $X=1.161 $Y=0.0675
c63 2 VSS 0.0588241f $X=1.107 $Y=0.0675
r64 65 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.125
+ $Y=0.136 $X2=1.143 $Y2=0.136
r65 63 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.136 $X2=1.143 $Y2=0.136
r66 61 68 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.136 $X2=1.089 $Y2=0.136
r67 61 65 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.136 $X2=1.125 $Y2=0.136
r68 59 60 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.167 $X2=1.089 $Y2=0.201
r69 58 60 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.225 $X2=1.089 $Y2=0.201
r70 57 68 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.145 $X2=1.089 $Y2=0.136
r71 57 59 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.145 $X2=1.089 $Y2=0.167
r72 55 56 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.069 $X2=1.089 $Y2=0.122
r73 54 68 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.127 $X2=1.089 $Y2=0.136
r74 54 56 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.127 $X2=1.089 $Y2=0.122
r75 53 55 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.089
+ $Y=0.045 $X2=1.089 $Y2=0.069
r76 48 58 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.08 $Y=0.234 $X2=1.089 $Y2=0.225
r77 48 50 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.026 $Y2=0.234
r78 45 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.036 $X2=1.026
+ $Y2=0.036
r79 43 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.08 $Y=0.036 $X2=1.089 $Y2=0.045
r80 43 45 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.036 $X2=1.026 $Y2=0.036
r81 42 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.234 $X2=1.026
+ $Y2=0.234
r82 39 42 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.2025 $X2=1.026 $Y2=0.2025
r83 38 42 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.043 $Y=0.2025 $X2=1.026 $Y2=0.2025
r84 37 46 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.026
+ $Y=0.0675 $X2=1.026 $Y2=0.036
r85 34 37 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.0675 $X2=1.026 $Y2=0.0675
r86 33 37 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.043 $Y=0.0675 $X2=1.026 $Y2=0.0675
r87 29 31 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.269
+ $Y=0.136 $X2=1.269 $Y2=0.2025
r88 26 29 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.269
+ $Y=0.0675 $X2=1.269 $Y2=0.136
r89 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.215
+ $Y=0.136 $X2=1.269 $Y2=0.136
r90 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.215
+ $Y=0.136 $X2=1.215 $Y2=0.2025
r91 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.215
+ $Y=0.0675 $X2=1.215 $Y2=0.136
r92 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.161
+ $Y=0.136 $X2=1.215 $Y2=0.136
r93 13 63 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.161 $Y=0.136 $X2=1.161
+ $Y2=0.136
r94 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.161
+ $Y=0.136 $X2=1.161 $Y2=0.2025
r95 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.161
+ $Y=0.0675 $X2=1.161 $Y2=0.136
r96 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.107
+ $Y=0.136 $X2=1.161 $Y2=0.136
r97 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.107
+ $Y=0.136 $X2=1.107 $Y2=0.2025
r98 2 5 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.107
+ $Y=0.0675 $X2=1.107 $Y2=0.136
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%Q 1 2 5 6 7 11 12 15 16 17 20 21 25 26 28 33 38
+ 40 43 46 49 52 VSS
c27 55 VSS 0.00197453f $X=1.134 $Y=0.234
c28 52 VSS 8.50672e-19 $X=1.134 $Y=0.216
c29 49 VSS 1.39487e-19 $X=1.134 $Y=0.0495
c30 46 VSS 6.94854e-19 $X=1.134 $Y=0.054
c31 43 VSS 0.00199537f $X=1.134 $Y=0.036
c32 42 VSS 0.00435712f $X=1.323 $Y=0.201
c33 40 VSS 0.0045092f $X=1.323 $Y=0.127
c34 39 VSS 0.0010981f $X=1.323 $Y=0.069
c35 38 VSS 9.20903e-19 $X=1.329 $Y=0.134
c36 36 VSS 0.0010981f $X=1.323 $Y=0.225
c37 34 VSS 0.00545672f $X=1.2085 $Y=0.234
c38 33 VSS 0.00256929f $X=1.175 $Y=0.234
c39 28 VSS 0.0155121f $X=1.313 $Y=0.234
c40 27 VSS 0.0054658f $X=1.2085 $Y=0.036
c41 26 VSS 0.0025515f $X=1.175 $Y=0.036
c42 25 VSS 0.00926069f $X=1.242 $Y=0.036
c43 21 VSS 0.0155121f $X=1.313 $Y=0.036
c44 20 VSS 0.00929505f $X=1.242 $Y=0.2025
c45 16 VSS 5.38922e-19 $X=1.259 $Y=0.2025
c46 15 VSS 0.0105438f $X=1.134 $Y=0.2025
c47 11 VSS 5.945e-19 $X=1.151 $Y=0.2025
c48 6 VSS 5.38922e-19 $X=1.259 $Y=0.0675
c49 5 VSS 0.010566f $X=1.134 $Y=0.0675
c50 1 VSS 5.945e-19 $X=1.151 $Y=0.0675
r51 56 57 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.225 $X2=1.134 $Y2=0.2295
r52 55 57 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.234 $X2=1.134 $Y2=0.2295
r53 52 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.216 $X2=1.134 $Y2=0.225
r54 48 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.045 $X2=1.134 $Y2=0.0495
r55 46 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.054 $X2=1.134 $Y2=0.0495
r56 43 48 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.036 $X2=1.134 $Y2=0.045
r57 41 42 3.3358 $w=2e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.145 $X2=1.323 $Y2=0.201
r58 39 40 3.45494 $w=2e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.069 $X2=1.323 $Y2=0.127
r59 38 41 0.655247 $w=2e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.134 $X2=1.323 $Y2=0.145
r60 38 40 0.416975 $w=2e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.134 $X2=1.323 $Y2=0.127
r61 36 42 1.42963 $w=2e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.225 $X2=1.323 $Y2=0.201
r62 35 39 1.42963 $w=2e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.045 $X2=1.323 $Y2=0.069
r63 33 34 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.175
+ $Y=0.234 $X2=1.2085 $Y2=0.234
r64 31 34 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.242
+ $Y=0.234 $X2=1.2085 $Y2=0.234
r65 29 55 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.143
+ $Y=0.234 $X2=1.134 $Y2=0.234
r66 29 33 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.143
+ $Y=0.234 $X2=1.175 $Y2=0.234
r67 28 36 0.685354 $w=2e-08 $l=1.3784e-08 $layer=M1 $thickness=3.6e-08 $X=1.313
+ $Y=0.234 $X2=1.323 $Y2=0.225
r68 28 31 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.313
+ $Y=0.234 $X2=1.242 $Y2=0.234
r69 26 27 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.175
+ $Y=0.036 $X2=1.2085 $Y2=0.036
r70 24 27 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=1.242
+ $Y=0.036 $X2=1.2085 $Y2=0.036
r71 24 25 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.242 $Y=0.036 $X2=1.242
+ $Y2=0.036
r72 22 43 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.143
+ $Y=0.036 $X2=1.134 $Y2=0.036
r73 22 26 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.143
+ $Y=0.036 $X2=1.175 $Y2=0.036
r74 21 35 0.685354 $w=2e-08 $l=1.3784e-08 $layer=M1 $thickness=3.6e-08 $X=1.313
+ $Y=0.036 $X2=1.323 $Y2=0.045
r75 21 24 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.313
+ $Y=0.036 $X2=1.242 $Y2=0.036
r76 20 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.242 $Y=0.234 $X2=1.242
+ $Y2=0.234
r77 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.225 $Y=0.2025 $X2=1.242 $Y2=0.2025
r78 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.259 $Y=0.2025 $X2=1.242 $Y2=0.2025
r79 15 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.134 $Y=0.216 $X2=1.134
+ $Y2=0.216
r80 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.117 $Y=0.2025 $X2=1.134 $Y2=0.2025
r81 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.151 $Y=0.2025 $X2=1.134 $Y2=0.2025
r82 10 25 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.242
+ $Y=0.0675 $X2=1.242 $Y2=0.036
r83 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.225 $Y=0.0675 $X2=1.242 $Y2=0.0675
r84 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.259 $Y=0.0675 $X2=1.242 $Y2=0.0675
r85 5 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.134 $Y=0.054 $X2=1.134
+ $Y2=0.054
r86 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.117
+ $Y=0.0675 $X2=1.134 $Y2=0.0675
r87 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.151
+ $Y=0.0675 $X2=1.134 $Y2=0.0675
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%13 1 6 9 VSS
c6 9 VSS 0.0277158f $X=0.38 $Y=0.0675
c7 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c8 4 VSS 3.22674e-19 $X=0.322 $Y=0.0675
r9 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r10 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%14 1 6 9 VSS
c10 9 VSS 0.022088f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.69239e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%15 1 6 9 VSS
c8 9 VSS 0.0223923f $X=0.758 $Y=0.0405
c9 6 VSS 3.14771e-19 $X=0.773 $Y=0.0405
c10 4 VSS 2.61968e-19 $X=0.7 $Y=0.0405
r11 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r12 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.7
+ $Y=0.0405 $X2=0.758 $Y2=0.0405
r13 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.685
+ $Y=0.0405 $X2=0.7 $Y2=0.0405
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%16 1 2 VSS
c0 1 VSS 0.00225696f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%17 1 2 VSS
c1 1 VSS 0.00201018f $X=0.341 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends

.subckt PM_DFFLQX4_ASAP7_75T_SRAM%18 1 2 VSS
c0 1 VSS 0.00219822f $X=0.773 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2295 $X2=0.739 $Y2=0.2295
.ends


* END of "./DFFLQx4_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DFFLQx4_ASAP7_75t_SRAM  VSS VDD CLK D Q
* 
* Q	Q
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_13_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_6_M3_g N_13_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_16_M4_d N_4_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_16_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_10_M7_d N_4_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.611
+ $Y=0.027
M8 N_15_M8_d N_6_M8_g N_10_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M9 VSS N_9_M9_g N_15_M9_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_9_M10_d N_10_M10_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.027
M11 N_11_M11_d N_10_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M12 N_11_M12_d N_10_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.027
M13 N_Q_M13_d N_11_M13_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.027
M14 N_Q_M14_d N_11_M14_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.151
+ $Y=0.027
M15 N_Q_M15_d N_11_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.027
M16 N_Q_M16_d N_11_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M17 VDD N_CLK_M17_g N_4_M17_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M18 N_6_M18_d N_4_M18_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M19 N_17_M19_d N_D_M19_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M20 N_8_M20_d N_4_M20_g N_17_M20_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M21 N_14_M21_d N_6_M21_g N_8_M21_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M22 VDD N_7_M22_g N_14_M22_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M23 N_7_M23_d N_8_M23_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M24 N_10_M24_d N_6_M24_g N_7_M24_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.665 $Y=0.216
M25 N_18_M25_d N_4_M25_g N_10_M25_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.719 $Y=0.216
M26 VDD N_9_M26_g N_18_M26_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M27 N_9_M27_d N_10_M27_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.827
+ $Y=0.216
M28 N_11_M28_d N_10_M28_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
M29 N_11_M29_d N_10_M29_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.162
M30 N_Q_M30_d N_11_M30_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.162
M31 N_Q_M31_d N_11_M31_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.151
+ $Y=0.162
M32 N_Q_M32_d N_11_M32_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.162
M33 N_Q_M33_d N_11_M33_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
*
* 
* .include "DFFLQx4_ASAP7_75t_SRAM.pex.sp.DFFLQX4_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DFFLQx4_ASAP7_75t_SRAM.pex.sp.DFFLQX4_ASAP7_75T_SRAM.pxi"
* File: DFFLQx4_ASAP7_75t_SRAM.pex.sp.DFFLQX4_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:26:46 2017
* 
x_PM_DFFLQX4_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M17_g CLK N_CLK_c_4_p
+ N_CLK_c_10_p VSS PM_DFFLQX4_ASAP7_75T_SRAM%CLK
x_PM_DFFLQX4_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_20_n N_4_M18_g N_4_c_34_p N_4_M20_g
+ N_4_M4_g N_4_M7_g N_4_c_77_p N_4_c_43_p N_4_M25_g N_4_c_89_p N_4_c_44_p
+ N_4_M0_s N_4_c_21_n N_4_M17_s N_4_c_22_n N_4_c_23_n N_4_c_24_n N_4_c_25_n
+ N_4_c_26_n N_4_c_27_n N_4_c_47_p N_4_c_28_n N_4_c_29_n N_4_c_30_n N_4_c_31_n
+ N_4_c_32_n N_4_c_58_p N_4_c_33_n N_4_c_36_p N_4_c_37_p N_4_c_38_p N_4_c_61_p
+ N_4_c_94_p N_4_c_46_p VSS PM_DFFLQX4_ASAP7_75T_SRAM%4
x_PM_DFFLQX4_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_122_n N_D_M19_g D N_D_c_123_n
+ N_D_c_133_p VSS PM_DFFLQX4_ASAP7_75T_SRAM%D
x_PM_DFFLQX4_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_147_n N_6_M21_g N_6_M8_g N_6_c_151_n
+ N_6_M24_g N_6_M1_d N_6_M18_d N_6_c_152_n N_6_c_172_n N_6_c_142_n N_6_c_154_n
+ N_6_c_143_n N_6_c_158_n N_6_c_174_n N_6_c_159_n N_6_c_161_n N_6_c_162_n
+ N_6_c_183_p N_6_c_168_n N_6_c_170_n N_6_c_144_n N_6_c_180_n N_6_c_181_n VSS
+ PM_DFFLQX4_ASAP7_75T_SRAM%6
x_PM_DFFLQX4_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_239_p N_7_M22_g N_7_M7_s N_7_M6_d
+ N_7_c_218_n N_7_M23_d N_7_c_219_n N_7_M24_s N_7_c_221_n N_7_c_237_p
+ N_7_c_230_n N_7_c_258_p N_7_c_231_n N_7_c_238_p N_7_c_223_n N_7_c_242_p
+ N_7_c_224_n N_7_c_225_n N_7_c_226_n N_7_c_256_p N_7_c_228_n N_7_c_235_n VSS
+ PM_DFFLQX4_ASAP7_75T_SRAM%7
x_PM_DFFLQX4_ASAP7_75T_SRAM%8 N_8_M6_g N_8_c_283_n N_8_M23_g N_8_M3_d N_8_M4_s
+ N_8_M20_d N_8_c_263_n N_8_M21_s N_8_c_313_p N_8_c_265_n N_8_c_287_n
+ N_8_c_314_p N_8_c_289_n N_8_c_266_n N_8_c_267_n N_8_c_302_n N_8_c_290_n
+ N_8_c_315_p N_8_c_268_n N_8_c_269_n N_8_c_271_n N_8_c_303_n N_8_c_275_n
+ N_8_c_304_n N_8_c_276_n N_8_c_278_n N_8_c_295_n N_8_c_308_n N_8_c_281_n VSS
+ PM_DFFLQX4_ASAP7_75T_SRAM%8
x_PM_DFFLQX4_ASAP7_75T_SRAM%9 N_9_M9_g N_9_c_323_p N_9_M26_g N_9_M10_d N_9_M27_d
+ N_9_c_322_p N_9_c_334_p N_9_c_321_p N_9_c_326_p N_9_c_320_p N_9_c_330_p
+ N_9_c_332_p N_9_c_339_p N_9_c_331_p N_9_c_335_p N_9_c_325_p N_9_c_333_p
+ N_9_c_336_p VSS PM_DFFLQX4_ASAP7_75T_SRAM%9
x_PM_DFFLQX4_ASAP7_75T_SRAM%10 N_10_M10_g N_10_c_354_n N_10_M27_g N_10_M11_g
+ N_10_M28_g N_10_M12_g N_10_c_396_p N_10_M29_g N_10_M8_s N_10_M7_d N_10_c_342_n
+ N_10_M25_s N_10_M24_d N_10_c_344_n N_10_c_376_n N_10_c_356_n N_10_c_357_n
+ N_10_c_409_p N_10_c_359_n N_10_c_368_n N_10_c_345_n N_10_c_346_n N_10_c_347_n
+ N_10_c_348_n N_10_c_381_n N_10_c_350_n N_10_c_382_n N_10_c_384_n N_10_c_385_n
+ N_10_c_386_n N_10_c_351_n N_10_c_352_n N_10_c_387_n N_10_c_361_n N_10_c_392_n
+ VSS PM_DFFLQX4_ASAP7_75T_SRAM%10
x_PM_DFFLQX4_ASAP7_75T_SRAM%11 N_11_M13_g N_11_M30_g N_11_M14_g N_11_M31_g
+ N_11_M15_g N_11_M32_g N_11_M16_g N_11_c_417_n N_11_M33_g N_11_M12_d N_11_M11_d
+ N_11_M29_d N_11_M28_d N_11_c_420_n N_11_c_412_n N_11_c_423_n N_11_c_413_n
+ N_11_c_426_n N_11_c_452_p N_11_c_453_p N_11_c_434_p N_11_c_442_p N_11_c_451_p
+ N_11_c_427_n VSS PM_DFFLQX4_ASAP7_75T_SRAM%11
x_PM_DFFLQX4_ASAP7_75T_SRAM%Q N_Q_M14_d N_Q_M13_d N_Q_c_456_n N_Q_M16_d N_Q_M15_d
+ N_Q_M31_d N_Q_M30_d N_Q_c_460_n N_Q_M33_d N_Q_M32_d N_Q_c_463_n N_Q_c_464_n
+ N_Q_c_466_n N_Q_c_467_n N_Q_c_470_n N_Q_c_472_n Q N_Q_c_476_n N_Q_c_477_n
+ N_Q_c_478_n N_Q_c_479_n N_Q_c_480_n VSS PM_DFFLQX4_ASAP7_75T_SRAM%Q
x_PM_DFFLQX4_ASAP7_75T_SRAM%13 N_13_M2_d N_13_M3_s N_13_c_482_n VSS
+ PM_DFFLQX4_ASAP7_75T_SRAM%13
x_PM_DFFLQX4_ASAP7_75T_SRAM%14 N_14_M21_d N_14_M22_s N_14_c_489_n VSS
+ PM_DFFLQX4_ASAP7_75T_SRAM%14
x_PM_DFFLQX4_ASAP7_75T_SRAM%15 N_15_M8_d N_15_M9_s N_15_c_498_n VSS
+ PM_DFFLQX4_ASAP7_75T_SRAM%15
x_PM_DFFLQX4_ASAP7_75T_SRAM%16 N_16_M5_s N_16_M4_d VSS PM_DFFLQX4_ASAP7_75T_SRAM%16
x_PM_DFFLQX4_ASAP7_75T_SRAM%17 N_17_M20_s N_17_M19_d VSS PM_DFFLQX4_ASAP7_75T_SRAM%17
x_PM_DFFLQX4_ASAP7_75T_SRAM%18 N_18_M26_s N_18_M25_d VSS PM_DFFLQX4_ASAP7_75T_SRAM%18
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_CLK_c_2_p N_4_c_20_n 0.00118333f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 CLK N_4_c_21_n 3.57152e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_4 N_CLK_c_4_p N_4_c_22_n 0.00206543f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.18
cc_5 CLK N_4_c_23_n 2.75361e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.07
cc_6 CLK N_4_c_24_n 0.00206543f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.125
cc_7 N_CLK_c_4_p N_4_c_25_n 2.75361e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2125
cc_8 CLK N_4_c_26_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_4_p N_4_c_27_n 5.03453e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_10_p N_4_c_28_n 8.76278e-19 $X=0.081 $Y=0.1305 $X2=0.145 $Y2=0.135
cc_11 N_CLK_c_4_p N_4_c_29_n 3.53054e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.164
cc_12 N_CLK_c_4_p N_4_c_30_n 6.09474e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.172
cc_13 N_CLK_c_4_p N_4_c_31_n 0.00138527f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.189
cc_14 N_CLK_c_4_p N_4_c_32_n 9.65218e-19 $X=0.081 $Y=0.135 $X2=0.159 $Y2=0.189
cc_15 N_CLK_c_4_p N_4_c_33_n 0.00167589f $X=0.081 $Y=0.135 $X2=0.229 $Y2=0.189
cc_16 CLK N_6_c_142_n 6.45949e-19 $X=0.082 $Y=0.119 $X2=0 $Y2=0
cc_17 N_CLK_c_4_p N_6_c_143_n 6.54444e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_18 CLK N_6_c_144_n 6.16145e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.234
cc_19 N_4_c_34_p N_D_M2_g 0.00341068f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.054
cc_20 N_4_c_34_p N_D_c_122_n 9.93922e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 N_4_c_36_p N_D_c_123_n 2.29805e-19 $X=0.29 $Y=0.189 $X2=0.081 $Y2=0.135
cc_22 N_4_c_37_p N_D_c_123_n 0.00102387f $X=0.513 $Y=0.189 $X2=0.081 $Y2=0.135
cc_23 N_4_c_38_p N_D_c_123_n 0.00337064f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_4_c_34_p N_6_M3_g 0.00355599f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.054
cc_25 N_4_M4_g N_6_M3_g 0.00355599f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_26 N_4_c_34_p N_6_c_147_n 9.91316e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_27 N_4_M7_g N_6_M8_g 0.00355599f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_28 N_4_c_43_p N_6_M8_g 0.00355599f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_29 N_4_c_44_p N_6_M8_g 0.00250099f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_30 N_4_c_44_p N_6_c_151_n 0.00180656f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_31 N_4_c_46_p N_6_c_152_n 0.00135022f $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_32 N_4_c_47_p N_6_c_142_n 0.00107729f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_33 N_4_c_36_p N_6_c_154_n 4.24027e-19 $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_34 N_4_c_32_n N_6_c_143_n 0.00285023f $X=0.159 $Y=0.189 $X2=0 $Y2=0
cc_35 N_4_c_33_n N_6_c_143_n 6.46981e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_36 N_4_c_46_p N_6_c_143_n 2.904e-19 $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_37 N_4_c_33_n N_6_c_158_n 4.24027e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_38 N_4_c_47_p N_6_c_159_n 0.00351854f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_39 N_4_c_36_p N_6_c_159_n 0.00102595f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_40 N_4_c_44_p N_6_c_161_n 6.63386e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_41 N_4_c_44_p N_6_c_162_n 0.00187197f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_42 N_4_c_29_n N_6_c_162_n 3.52457e-19 $X=0.189 $Y=0.164 $X2=0 $Y2=0
cc_43 N_4_c_58_p N_6_c_162_n 2.46239e-19 $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_44 N_4_c_36_p N_6_c_162_n 0.0253778f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_45 N_4_c_38_p N_6_c_162_n 0.00115493f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_61_p N_6_c_162_n 2.81476e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_47 N_4_c_37_p N_6_c_168_n 2.98936e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_48 N_4_c_38_p N_6_c_168_n 0.00170246f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_49 N_4_c_44_p N_6_c_170_n 0.00124003f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_50 N_4_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_51 N_4_M7_g N_7_M5_g 2.13359e-19 $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_52 N_4_c_44_p N_7_M5_g 0.00205839f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_53 N_4_c_61_p N_7_M5_g 3.15189e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_54 N_4_c_44_p N_7_c_218_n 5.50331e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.135
cc_55 N_4_c_44_p N_7_c_219_n 2.12581e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.1305
cc_56 N_4_c_44_p N_7_M24_s 2.50995e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_57 N_4_M7_g N_7_c_221_n 0.00200088f $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_58 N_4_c_44_p N_7_c_221_n 0.00303373f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_59 N_4_M7_g N_7_c_223_n 2.97268e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_60 N_4_M7_g N_7_c_224_n 2.21692e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_61 N_4_c_61_p N_7_c_225_n 5.74745e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_62 N_4_c_77_p N_7_c_226_n 0.00193027f $X=0.621 $Y=0.178 $X2=0 $Y2=0
cc_63 N_4_c_44_p N_7_c_226_n 0.00189849f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_64 N_4_M7_g N_7_c_228_n 3.80981e-19 $X=0.621 $Y=0.0405 $X2=0 $Y2=0
cc_65 N_4_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_66 N_4_M7_g N_8_M6_g 0.00341068f $X=0.621 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_67 N_4_c_44_p N_8_M6_g 0.00303187f $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.054
cc_68 N_4_c_37_p N_8_c_263_n 3.15319e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_69 N_4_c_38_p N_8_c_263_n 0.00136448f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_70 N_4_c_37_p N_8_c_265_n 0.00161272f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_71 N_4_M4_g N_8_c_266_n 3.80535e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_72 N_4_M4_g N_8_c_267_n 2.08362e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_73 N_4_M4_g N_8_c_268_n 2.25982e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_74 N_4_c_89_p N_8_c_269_n 2.70413e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_75 N_4_c_61_p N_8_c_269_n 0.00174159f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_76 N_4_c_89_p N_8_c_271_n 0.0017128f $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_77 N_4_c_44_p N_8_c_271_n 5.88593e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_78 N_4_c_37_p N_8_c_271_n 0.00102123f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_79 N_4_c_94_p N_8_c_271_n 3.42482e-19 $X=0.351 $Y=0.178 $X2=0 $Y2=0
cc_80 N_4_c_44_p N_8_c_275_n 8.16411e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_81 N_4_c_44_p N_8_c_276_n 3.32592e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_82 N_4_c_61_p N_8_c_276_n 8.9822e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_83 N_4_c_44_p N_8_c_278_n 5.02733e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_84 N_4_c_43_p N_9_M9_g 0.00341068f $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_85 N_4_c_43_p N_10_M10_g 2.13359e-19 $X=0.729 $Y=0.178 $X2=0.081 $Y2=0.054
cc_86 N_4_c_44_p N_10_c_342_n 8.28378e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_87 N_4_c_44_p N_10_M25_s 3.37661e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_88 N_4_c_44_p N_10_c_344_n 0.00134632f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_89 N_4_c_43_p N_10_c_345_n 2.69517e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_90 N_4_c_43_p N_10_c_346_n 2.11116e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_91 N_4_c_43_p N_10_c_347_n 2.5872e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_92 N_4_c_43_p N_10_c_348_n 0.00229157f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_93 N_4_c_44_p N_10_c_348_n 7.89371e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_94 N_4_c_43_p N_10_c_350_n 3.99306e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_95 N_4_c_44_p N_10_c_351_n 4.45535e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_96 N_4_c_43_p N_10_c_352_n 4.71808e-19 $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_97 N_4_c_44_p N_10_c_352_n 2.2968e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_98 N_4_c_34_p N_13_c_482_n 0.00526789f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_99 N_4_c_44_p N_14_M22_s 2.36286e-19 $X=0.725 $Y=0.178 $X2=0.081 $Y2=0.216
cc_100 N_4_M4_g N_14_c_489_n 0.00200088f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_101 N_4_c_89_p N_14_c_489_n 5.41258e-19 $X=0.464 $Y=0.178 $X2=0 $Y2=0
cc_102 N_4_c_44_p N_14_c_489_n 0.00230928f $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_103 N_4_c_37_p N_14_c_489_n 7.09553e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_104 N_4_c_43_p N_15_c_498_n 0.0019841f $X=0.729 $Y=0.178 $X2=0 $Y2=0
cc_105 N_4_c_44_p N_15_c_498_n 4.3039e-19 $X=0.725 $Y=0.178 $X2=0 $Y2=0
cc_106 N_D_M2_g N_6_M3_g 2.82885e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_107 D N_6_c_172_n 0.00115224f $X=0.298 $Y=0.082 $X2=0 $Y2=0
cc_108 N_D_c_123_n N_6_c_154_n 0.00115224f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_109 N_D_c_123_n N_6_c_174_n 0.00115224f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_110 N_D_c_123_n N_6_c_159_n 0.00124565f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_111 D N_6_c_162_n 2.27807e-19 $X=0.298 $Y=0.082 $X2=0 $Y2=0
cc_112 N_D_c_123_n N_6_c_162_n 9.62099e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_113 N_D_c_133_p N_6_c_168_n 4.3159e-19 $X=0.297 $Y=0.126 $X2=0 $Y2=0
cc_114 D N_6_c_144_n 0.00115224f $X=0.298 $Y=0.082 $X2=0 $Y2=0
cc_115 N_D_c_133_p N_6_c_180_n 0.00115224f $X=0.297 $Y=0.126 $X2=0 $Y2=0
cc_116 N_D_c_123_n N_6_c_181_n 0.00115224f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_117 N_D_c_123_n N_8_c_263_n 3.88702e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_118 N_D_c_123_n N_8_c_265_n 8.77202e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_119 D N_8_c_281_n 2.04306e-19 $X=0.298 $Y=0.082 $X2=0 $Y2=0
cc_120 D N_13_c_482_n 0.00430488f $X=0.298 $Y=0.082 $X2=0 $Y2=0
cc_121 N_D_c_123_n N_17_M20_s 3.05674e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.054
cc_122 N_6_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_123 N_6_c_183_p N_7_c_230_n 2.96121e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_124 N_6_c_161_n N_7_c_231_n 2.61213e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_125 N_6_c_183_p N_7_c_231_n 2.61213e-19 $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_126 N_6_c_170_n N_7_c_223_n 0.00327734f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_127 N_6_c_161_n N_7_c_224_n 0.00115177f $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_128 N_6_c_161_n N_7_c_235_n 2.96121e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_129 N_6_M8_g N_8_M6_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_130 N_6_c_147_n N_8_c_283_n 2.04136e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_131 N_6_c_151_n N_8_c_283_n 4.12331e-19 $X=0.675 $Y=0.135 $X2=0.081 $Y2=0.135
cc_132 N_6_c_183_p N_8_c_283_n 2.64012e-19 $X=0.601 $Y=0.153 $X2=0.081 $Y2=0.135
cc_133 N_6_c_168_n N_8_c_263_n 2.25088e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_134 N_6_M3_g N_8_c_287_n 3.49806e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_135 N_6_c_168_n N_8_c_287_n 3.83282e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_136 N_6_c_168_n N_8_c_289_n 9.7435e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_137 N_6_c_168_n N_8_c_290_n 9.7435e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_138 N_6_c_162_n N_8_c_268_n 0.00118282f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_139 N_6_c_168_n N_8_c_268_n 0.00106776f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_140 N_6_c_162_n N_8_c_275_n 0.00138951f $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_141 N_6_c_183_p N_8_c_278_n 0.00138951f $X=0.601 $Y=0.153 $X2=0 $Y2=0
cc_142 N_6_c_162_n N_8_c_295_n 2.54113e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_143 N_6_c_162_n N_8_c_281_n 3.92135e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_144 N_6_M8_g N_9_M9_g 2.82885e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_145 N_6_c_151_n N_10_c_354_n 2.73247e-19 $X=0.675 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_146 N_6_c_161_n N_10_c_342_n 2.24654e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_147 N_6_c_161_n N_10_c_356_n 5.06919e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_148 N_6_M8_g N_10_c_357_n 3.43727e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_149 N_6_c_170_n N_10_c_357_n 5.96743e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_150 N_6_c_161_n N_10_c_359_n 2.34004e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_151 N_6_c_170_n N_10_c_346_n 0.00329665f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_152 N_6_c_161_n N_10_c_361_n 2.83245e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_153 N_6_c_162_n N_13_c_482_n 8.35084e-19 $X=0.527 $Y=0.153 $X2=0 $Y2=0
cc_154 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_155 N_7_c_237_p N_8_M6_g 3.91159e-19 $X=0.581 $Y=0.09 $X2=0.135 $Y2=0.054
cc_156 N_7_c_238_p N_8_c_266_n 2.03196e-19 $X=0.594 $Y=0.054 $X2=0.464 $Y2=0.178
cc_157 N_7_c_239_p N_8_c_267_n 3.19692e-19 $X=0.513 $Y=0.09 $X2=0 $Y2=0
cc_158 N_7_c_237_p N_8_c_267_n 0.00107929f $X=0.581 $Y=0.09 $X2=0 $Y2=0
cc_159 N_7_c_223_n N_8_c_302_n 2.36738e-19 $X=0.621 $Y=0.122 $X2=0 $Y2=0
cc_160 N_7_c_242_p N_8_c_303_n 9.84729e-19 $X=0.621 $Y=0.14 $X2=0.056 $Y2=0.054
cc_161 N_7_c_237_p N_8_c_304_n 0.00507595f $X=0.581 $Y=0.09 $X2=0 $Y2=0
cc_162 N_7_M5_g N_8_c_276_n 3.12986e-19 $X=0.513 $Y=0.0405 $X2=0.071 $Y2=0.216
cc_163 N_7_c_239_p N_8_c_295_n 5.2508e-19 $X=0.513 $Y=0.09 $X2=0.018 $Y2=0.18
cc_164 N_7_c_218_n N_8_c_295_n 3.88009e-19 $X=0.594 $Y=0.0405 $X2=0.018 $Y2=0.18
cc_165 N_7_c_238_p N_8_c_308_n 2.03196e-19 $X=0.594 $Y=0.054 $X2=0.018 $Y2=0.125
cc_166 N_7_c_218_n N_10_c_342_n 0.00311119f $X=0.594 $Y=0.0405 $X2=0 $Y2=0
cc_167 N_7_c_238_p N_10_c_342_n 3.00222e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_168 N_7_c_228_n N_10_c_342_n 2.2454e-19 $X=0.621 $Y=0.09 $X2=0 $Y2=0
cc_169 N_7_c_221_n N_10_c_344_n 0.00207384f $X=0.65 $Y=0.2295 $X2=0 $Y2=0
cc_170 N_7_c_218_n N_10_c_356_n 3.50513e-19 $X=0.594 $Y=0.0405 $X2=0 $Y2=0
cc_171 N_7_c_238_p N_10_c_356_n 5.0339e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_172 N_7_c_238_p N_10_c_368_n 2.21141e-19 $X=0.594 $Y=0.054 $X2=0 $Y2=0
cc_173 N_7_c_228_n N_10_c_345_n 4.33699e-19 $X=0.621 $Y=0.09 $X2=0.071 $Y2=0.054
cc_174 N_7_c_256_p N_10_c_348_n 4.33699e-19 $X=0.621 $Y=0.214 $X2=0 $Y2=0
cc_175 N_7_c_221_n N_10_c_351_n 3.64454e-19 $X=0.65 $Y=0.2295 $X2=0.054
+ $Y2=0.234
cc_176 N_7_c_258_p N_10_c_351_n 4.86017e-19 $X=0.612 $Y=0.234 $X2=0.054
+ $Y2=0.234
cc_177 N_7_c_226_n N_10_c_352_n 4.33699e-19 $X=0.621 $Y=0.203 $X2=0.0505
+ $Y2=0.234
cc_178 N_8_c_263_n N_13_c_482_n 0.00119636f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.135
cc_179 N_8_c_295_n N_13_c_482_n 0.00362439f $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_180 N_8_c_281_n N_13_c_482_n 4.41747e-19 $X=0.45 $Y=0.036 $X2=0.351 $Y2=0.135
cc_181 N_8_c_263_n N_14_c_489_n 0.0018138f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.135
cc_182 N_8_c_313_p N_14_c_489_n 0.00209454f $X=0.45 $Y=0.234 $X2=0.351 $Y2=0.135
cc_183 N_8_c_314_p N_14_c_489_n 0.0013184f $X=0.434 $Y=0.234 $X2=0.351 $Y2=0.135
cc_184 N_8_c_315_p N_14_c_489_n 0.00116161f $X=0.459 $Y=0.225 $X2=0.351
+ $Y2=0.135
cc_185 N_8_c_295_n N_14_c_489_n 6.06615e-19 $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_186 N_9_M9_g N_10_M10_g 0.00268443f $X=0.783 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_187 N_9_c_320_p N_10_M10_g 3.74489e-19 $X=0.846 $Y=0.036 $X2=0.135 $Y2=0.054
cc_188 N_9_c_321_p N_10_c_376_n 0.00141609f $X=0.792 $Y=0.036 $X2=0.464
+ $Y2=0.178
cc_189 N_9_c_322_p N_10_c_368_n 0.00141609f $X=0.783 $Y=0.105 $X2=0 $Y2=0
cc_190 N_9_c_323_p N_10_c_345_n 3.34766e-19 $X=0.783 $Y=0.1055 $X2=0.071
+ $Y2=0.054
cc_191 N_9_c_322_p N_10_c_345_n 0.00141609f $X=0.783 $Y=0.105 $X2=0.071
+ $Y2=0.054
cc_192 N_9_c_325_p N_10_c_348_n 2.26874e-19 $X=0.945 $Y=0.225 $X2=0 $Y2=0
cc_193 N_9_c_326_p N_10_c_381_n 2.61208e-19 $X=0.828 $Y=0.036 $X2=0.071
+ $Y2=0.216
cc_194 N_9_M9_g N_10_c_382_n 6.3699e-19 $X=0.783 $Y=0.0405 $X2=0.056 $Y2=0.216
cc_195 N_9_c_322_p N_10_c_382_n 9.0998e-19 $X=0.783 $Y=0.105 $X2=0.056 $Y2=0.216
cc_196 N_9_c_320_p N_10_c_384_n 4.40983e-19 $X=0.846 $Y=0.036 $X2=0.018 $Y2=0.18
cc_197 N_9_c_330_p N_10_c_385_n 5.09066e-19 $X=0.882 $Y=0.036 $X2=0.027
+ $Y2=0.036
cc_198 N_9_c_331_p N_10_c_386_n 0.00148937f $X=0.9 $Y=0.234 $X2=0.054 $Y2=0.036
cc_199 N_9_c_332_p N_10_c_387_n 4.52584e-19 $X=0.9 $Y=0.036 $X2=0.135 $Y2=0.135
cc_200 N_9_c_333_p N_10_c_387_n 0.00280793f $X=0.945 $Y=0.122 $X2=0.135
+ $Y2=0.135
cc_201 N_9_c_334_p N_10_c_361_n 2.40515e-19 $X=0.936 $Y=0.036 $X2=0.145
+ $Y2=0.135
cc_202 N_9_c_335_p N_10_c_361_n 7.44774e-19 $X=0.918 $Y=0.234 $X2=0.145
+ $Y2=0.135
cc_203 N_9_c_336_p N_10_c_361_n 8.84468e-19 $X=0.945 $Y=0.167 $X2=0.145
+ $Y2=0.135
cc_204 N_9_c_336_p N_10_c_392_n 0.00213032f $X=0.945 $Y=0.167 $X2=0.033
+ $Y2=0.189
cc_205 N_9_c_334_p N_11_c_412_n 4.57392e-19 $X=0.936 $Y=0.036 $X2=0.725
+ $Y2=0.178
cc_206 N_9_c_339_p N_11_c_413_n 4.495e-19 $X=0.936 $Y=0.234 $X2=0.056 $Y2=0.054
cc_207 N_9_c_321_p N_15_c_498_n 7.33799e-19 $X=0.792 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_208 N_10_M11_g N_11_M13_g 2.13359e-19 $X=0.999 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_209 N_10_M12_g N_11_M13_g 0.00268443f $X=1.053 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_210 N_10_M12_g N_11_M14_g 2.13359e-19 $X=1.053 $Y=0.0675 $X2=0.351 $Y2=0.135
cc_211 N_10_c_396_p N_11_c_417_n 0.00102658f $X=1.053 $Y=0.136 $X2=0 $Y2=0
cc_212 N_10_c_396_p N_11_M12_d 3.7444e-19 $X=1.053 $Y=0.136 $X2=0.459 $Y2=0.178
cc_213 N_10_c_396_p N_11_M29_d 3.85232e-19 $X=1.053 $Y=0.136 $X2=0 $Y2=0
cc_214 N_10_c_396_p N_11_c_420_n 8.43851e-19 $X=1.053 $Y=0.136 $X2=0.725
+ $Y2=0.178
cc_215 N_10_M12_g N_11_c_412_n 4.61823e-19 $X=1.053 $Y=0.0675 $X2=0.725
+ $Y2=0.178
cc_216 N_10_c_396_p N_11_c_412_n 5.30021e-19 $X=1.053 $Y=0.136 $X2=0.725
+ $Y2=0.178
cc_217 N_10_c_396_p N_11_c_423_n 7.60428e-19 $X=1.053 $Y=0.136 $X2=0 $Y2=0
cc_218 N_10_M12_g N_11_c_413_n 4.56718e-19 $X=1.053 $Y=0.0675 $X2=0.056
+ $Y2=0.054
cc_219 N_10_c_396_p N_11_c_413_n 5.38938e-19 $X=1.053 $Y=0.136 $X2=0.056
+ $Y2=0.054
cc_220 N_10_c_392_n N_11_c_426_n 0.00103215f $X=0.999 $Y=0.136 $X2=0 $Y2=0
cc_221 N_10_c_361_n N_11_c_427_n 3.06386e-19 $X=0.999 $Y=0.153 $X2=0.054
+ $Y2=0.036
cc_222 N_10_c_342_n N_15_c_498_n 0.0018138f $X=0.648 $Y=0.0405 $X2=0.351
+ $Y2=0.135
cc_223 N_10_c_376_n N_15_c_498_n 0.00205226f $X=0.72 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_224 N_10_c_409_p N_15_c_498_n 0.0013184f $X=0.704 $Y=0.036 $X2=0.351
+ $Y2=0.135
cc_225 N_10_c_368_n N_15_c_498_n 0.00103564f $X=0.729 $Y=0.081 $X2=0.351
+ $Y2=0.135
cc_226 N_10_c_350_n N_15_c_498_n 4.47528e-19 $X=0.774 $Y=0.162 $X2=0.351
+ $Y2=0.135
cc_227 N_11_c_417_n N_Q_M14_d 3.73731e-19 $X=1.269 $Y=0.136 $X2=0.783 $Y2=0.0405
cc_228 N_11_c_412_n N_Q_c_456_n 0.00118764f $X=1.08 $Y=0.036 $X2=0.783
+ $Y2=0.1055
cc_229 N_11_c_423_n N_Q_c_456_n 2.62013e-19 $X=1.026 $Y=0.036 $X2=0.783
+ $Y2=0.1055
cc_230 N_11_c_417_n N_Q_M16_d 3.7444e-19 $X=1.269 $Y=0.136 $X2=0.783 $Y2=0.2295
cc_231 N_11_c_417_n N_Q_M31_d 3.8685e-19 $X=1.269 $Y=0.136 $X2=0 $Y2=0
cc_232 N_11_c_420_n N_Q_c_460_n 2.68378e-19 $X=1.026 $Y=0.2025 $X2=0.862
+ $Y2=0.2295
cc_233 N_11_c_434_p N_Q_c_460_n 0.00118419f $X=1.089 $Y=0.167 $X2=0.862
+ $Y2=0.2295
cc_234 N_11_c_417_n N_Q_M33_d 3.87022e-19 $X=1.269 $Y=0.136 $X2=0 $Y2=0
cc_235 N_11_c_417_n N_Q_c_463_n 8.43851e-19 $X=1.269 $Y=0.136 $X2=0.783
+ $Y2=0.105
cc_236 N_11_M15_g N_Q_c_464_n 3.57913e-19 $X=1.215 $Y=0.0675 $X2=0.783 $Y2=0.105
cc_237 N_11_M16_g N_Q_c_464_n 4.61823e-19 $X=1.269 $Y=0.0675 $X2=0.783 $Y2=0.105
cc_238 N_11_c_417_n N_Q_c_466_n 7.60428e-19 $X=1.269 $Y=0.136 $X2=0.936
+ $Y2=0.036
cc_239 N_11_M14_g N_Q_c_467_n 4.31409e-19 $X=1.161 $Y=0.0675 $X2=0.792 $Y2=0.036
cc_240 N_11_c_417_n N_Q_c_467_n 0.00142439f $X=1.269 $Y=0.136 $X2=0.792
+ $Y2=0.036
cc_241 N_11_c_442_p N_Q_c_467_n 5.02824e-19 $X=1.161 $Y=0.136 $X2=0.792
+ $Y2=0.036
cc_242 N_11_M15_g N_Q_c_470_n 3.53956e-19 $X=1.215 $Y=0.0675 $X2=0.864 $Y2=0.036
cc_243 N_11_M16_g N_Q_c_470_n 4.56718e-19 $X=1.269 $Y=0.0675 $X2=0.864 $Y2=0.036
cc_244 N_11_M14_g N_Q_c_472_n 3.94108e-19 $X=1.161 $Y=0.0675 $X2=0.9 $Y2=0.036
cc_245 N_11_c_417_n N_Q_c_472_n 0.00145408f $X=1.269 $Y=0.136 $X2=0.9 $Y2=0.036
cc_246 N_11_c_413_n N_Q_c_472_n 0.0013429f $X=1.08 $Y=0.234 $X2=0.9 $Y2=0.036
cc_247 N_11_c_442_p N_Q_c_472_n 5.18971e-19 $X=1.161 $Y=0.136 $X2=0.9 $Y2=0.036
cc_248 N_11_c_417_n N_Q_c_476_n 4.1631e-19 $X=1.269 $Y=0.136 $X2=0.918 $Y2=0.234
cc_249 N_11_c_412_n N_Q_c_477_n 0.00134363f $X=1.08 $Y=0.036 $X2=0.945 $Y2=0.117
cc_250 N_11_c_451_p N_Q_c_478_n 2.95672e-19 $X=1.143 $Y=0.136 $X2=0.945
+ $Y2=0.171
cc_251 N_11_c_452_p N_Q_c_479_n 0.00134363f $X=1.089 $Y=0.069 $X2=0 $Y2=0
cc_252 N_11_c_453_p N_Q_c_480_n 0.0013429f $X=1.089 $Y=0.225 $X2=0 $Y2=0
cc_253 N_11_c_451_p N_Q_c_480_n 3.06781e-19 $X=1.143 $Y=0.136 $X2=0 $Y2=0

* END of "./DFFLQx4_ASAP7_75t_SRAM.pex.sp.DFFLQX4_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: SDFHx1_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 13:03:02 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "SDFHx1_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./SDFHx1_ASAP7_75t_SRAM.pex.sp.pex"
* File: SDFHx1_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 13:03:02 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_SDFHX1_ASAP7_75T_SRAM%CLK 2 5 7 11 16 18 19 20 VSS
c19 20 VSS 1.17072e-19 $X=0.081 $Y=0.1785
c20 19 VSS 3.55344e-20 $X=0.081 $Y=0.167
c21 18 VSS 9.34089e-20 $X=0.081 $Y=0.162
c22 16 VSS 0.00100628f $X=0.078 $Y=0.19
c23 11 VSS 0.00681069f $X=0.081 $Y=0.135
c24 5 VSS 0.00208806f $X=0.081 $Y=0.135
c25 2 VSS 0.0627545f $X=0.081 $Y=0.054
r26 19 20 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.167 $X2=0.081 $Y2=0.1785
r27 18 19 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.162 $X2=0.081 $Y2=0.167
r28 17 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.144 $X2=0.081 $Y2=0.162
r29 16 20 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.19 $X2=0.081 $Y2=0.1785
r30 11 17 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.144
r31 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r32 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r33 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%4 2 5 7 10 13 15 18 21 23 25 28 30 36 37 38 41 45
+ 52 59 64 71 72 73 74 75 77 79 80 84 92 VSS
c66 111 VSS 1.06551e-19 $X=0.03 $Y=0.153
c67 110 VSS 6.89947e-19 $X=0.027 $Y=0.153
c68 92 VSS 0.001222f $X=0.891 $Y=0.135
c69 84 VSS 0.00111816f $X=0.135 $Y=0.135
c70 80 VSS 0.0020506f $X=0.817 $Y=0.153
c71 79 VSS 0.00159119f $X=0.743 $Y=0.153
c72 77 VSS 0.00276317f $X=0.891 $Y=0.153
c73 75 VSS 0.0014306f $X=0.479 $Y=0.153
c74 74 VSS 0.00120845f $X=0.337 $Y=0.153
c75 73 VSS 9.39788e-19 $X=0.211 $Y=0.153
c76 72 VSS 0.00665478f $X=0.175 $Y=0.153
c77 71 VSS 9.40943e-19 $X=0.621 $Y=0.153
c78 64 VSS 6.72589e-19 $X=0.033 $Y=0.153
c79 59 VSS 5.26559e-19 $X=0.621 $Y=0.135
c80 55 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c81 54 VSS 0.00180216f $X=0.047 $Y=0.234
c82 52 VSS 0.00253483f $X=0.054 $Y=0.234
c83 50 VSS 0.00305101f $X=0.027 $Y=0.234
c84 48 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c85 47 VSS 0.00199699f $X=0.047 $Y=0.036
c86 45 VSS 0.00239525f $X=0.054 $Y=0.036
c87 43 VSS 0.00305101f $X=0.027 $Y=0.036
c88 42 VSS 5.16336e-19 $X=0.018 $Y=0.2125
c89 41 VSS 0.00180713f $X=0.018 $Y=0.2
c90 40 VSS 4.96914e-19 $X=0.018 $Y=0.225
c91 38 VSS 0.00159315f $X=0.018 $Y=0.1125
c92 37 VSS 0.00142827f $X=0.018 $Y=0.081
c93 36 VSS 0.00143809f $X=0.018 $Y=0.144
c94 33 VSS 0.0049466f $X=0.056 $Y=0.216
c95 30 VSS 2.98509e-19 $X=0.071 $Y=0.216
c96 28 VSS 0.00460164f $X=0.056 $Y=0.054
c97 25 VSS 2.98509e-19 $X=0.071 $Y=0.054
c98 21 VSS 0.00216055f $X=0.891 $Y=0.135
c99 18 VSS 0.0585656f $X=0.891 $Y=0.0405
c100 13 VSS 0.00201792f $X=0.621 $Y=0.135
c101 10 VSS 0.0601628f $X=0.621 $Y=0.0675
c102 5 VSS 0.00199564f $X=0.135 $Y=0.135
c103 2 VSS 0.0630095f $X=0.135 $Y=0.054
r104 110 111 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r105 107 110 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r106 79 80 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.743
+ $Y=0.153 $X2=0.817 $Y2=0.153
r107 77 80 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.817 $Y2=0.153
r108 77 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r109 74 75 9.64198 $w=1.8e-08 $l=1.42e-07 $layer=M2 $thickness=3.6e-08 $X=0.337
+ $Y=0.153 $X2=0.479 $Y2=0.153
r110 73 74 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.211
+ $Y=0.153 $X2=0.337 $Y2=0.153
r111 72 73 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.175
+ $Y=0.153 $X2=0.211 $Y2=0.153
r112 70 79 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.743 $Y2=0.153
r113 70 75 9.64198 $w=1.8e-08 $l=1.42e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.479 $Y2=0.153
r114 70 71 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.621 $Y=0.153 $X2=0.621
+ $Y2=0.153
r115 67 72 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.153 $X2=0.175 $Y2=0.153
r116 67 84 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.135 $Y=0.153 $X2=0.135
+ $Y2=0.153
r117 64 111 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r118 63 67 6.92593 $w=1.8e-08 $l=1.02e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.135 $Y2=0.153
r119 63 64 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r120 59 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.153
r121 54 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r122 52 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r123 50 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r124 47 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r125 45 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r126 43 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r127 41 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r128 40 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r129 40 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r130 39 107 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r131 39 41 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.2
r132 37 38 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.1125
r133 36 107 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r134 36 38 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1125
r135 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r136 35 37 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r137 33 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r138 30 33 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r139 28 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r140 25 28 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r141 21 92 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.135 $X2=0.891
+ $Y2=0.135
r142 21 23 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.135 $X2=0.891 $Y2=0.2295
r143 18 21 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.0405 $X2=0.891 $Y2=0.135
r144 13 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r145 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2295
r146 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r147 5 84 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r148 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r149 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%SE 2 5 7 10 13 15 19 22 23 24 31 33 41 44 45 46 47
+ 54 58 59 62 63 VSS
c79 63 VSS 2.09605e-19 $X=1.215 $Y=0.113
c80 62 VSS 0.0013442f $X=1.215 $Y=0.09
c81 59 VSS 2.63823e-19 $X=0.225 $Y=0.099
c82 58 VSS 5.90201e-19 $X=0.225 $Y=0.081
c83 54 VSS 0.001241f $X=1.215 $Y=0.136
c84 47 VSS 0.0382892f $X=1.175 $Y=0.045
c85 46 VSS 0.00642311f $X=0.337 $Y=0.045
c86 45 VSS 0.00708959f $X=1.215 $Y=0.045
c87 44 VSS 0.00320338f $X=1.215 $Y=0.045
c88 41 VSS 0.00531f $X=0.225 $Y=0.045
c89 31 VSS 0.00110873f $X=0.225 $Y=0.126
c90 24 VSS 2.51525e-19 $X=0.279 $Y=0.135
c91 23 VSS 1.48251e-19 $X=0.261 $Y=0.135
c92 22 VSS 6.38823e-20 $X=0.258 $Y=0.135
c93 21 VSS 0.00134071f $X=0.255 $Y=0.135
c94 19 VSS 6.89032e-19 $X=0.297 $Y=0.135
c95 13 VSS 0.00257518f $X=1.215 $Y=0.136
c96 10 VSS 0.0624472f $X=1.215 $Y=0.0405
c97 5 VSS 0.00319967f $X=0.297 $Y=0.135
c98 2 VSS 0.063344f $X=0.297 $Y=0.0675
r99 62 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.09 $X2=1.215 $Y2=0.113
r100 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.081 $X2=0.225 $Y2=0.099
r101 54 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.136 $X2=1.215 $Y2=0.113
r102 46 47 56.9012 $w=1.8e-08 $l=8.38e-07 $layer=M2 $thickness=3.6e-08 $X=0.337
+ $Y=0.045 $X2=1.175 $Y2=0.045
r103 45 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.215 $Y2=0.09
r104 44 47 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.175 $Y2=0.045
r105 44 45 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.215 $Y=0.045 $X2=1.215
+ $Y2=0.045
r106 41 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.081
r107 40 46 7.60494 $w=1.8e-08 $l=1.12e-07 $layer=M2 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.337 $Y2=0.045
r108 40 41 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.225 $Y=0.045 $X2=0.225
+ $Y2=0.045
r109 31 59 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.099
r110 31 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r111 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.135 $X2=0.279 $Y2=0.135
r112 22 23 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.258
+ $Y=0.135 $X2=0.261 $Y2=0.135
r113 21 22 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.255
+ $Y=0.135 $X2=0.258 $Y2=0.135
r114 19 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.279 $Y2=0.135
r115 17 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.225 $Y2=0.135
r116 17 21 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.255 $Y2=0.135
r117 13 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.215 $Y=0.136 $X2=1.215
+ $Y2=0.136
r118 13 15 350.298 $w=2e-08 $l=9.35e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.136 $X2=1.215 $Y2=0.2295
r119 10 13 357.791 $w=2e-08 $l=9.55e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.0405 $X2=1.215 $Y2=0.136
r120 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r121 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r122 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%6 2 5 7 9 12 14 17 23 26 28 29 33 36 38 39 43 51
+ 57 58 65 VSS
c69 65 VSS 3.41193e-19 $X=1.161 $Y=0.2125
c70 58 VSS 5.45782e-19 $X=0.351 $Y=0.126
c71 57 VSS 8.0335e-19 $X=0.351 $Y=0.099
c72 51 VSS 0.00325146f $X=1.161 $Y=0.049
c73 43 VSS 3.66031e-19 $X=0.351 $Y=0.135
c74 39 VSS 9.89222e-19 $X=0.936 $Y=0.081
c75 38 VSS 0.00675922f $X=0.9 $Y=0.081
c76 36 VSS 0.00169093f $X=1.161 $Y=0.081
c77 33 VSS 8.10983e-19 $X=0.351 $Y=0.081
c78 29 VSS 7.48824e-19 $X=1.179 $Y=0.234
c79 28 VSS 0.00240687f $X=1.17 $Y=0.234
c80 26 VSS 0.00328115f $X=1.188 $Y=0.234
c81 23 VSS 8.98553e-20 $X=1.161 $Y=0.225
c82 17 VSS 0.0040579f $X=1.19 $Y=0.2295
c83 14 VSS 2.95772e-19 $X=1.205 $Y=0.2295
c84 12 VSS 0.0608204f $X=1.19 $Y=0.0405
c85 9 VSS 3.14771e-19 $X=1.205 $Y=0.0405
c86 5 VSS 0.00125227f $X=0.351 $Y=0.135
c87 2 VSS 0.0585837f $X=0.351 $Y=0.0675
r88 64 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.2 $X2=1.161 $Y2=0.2125
r89 57 58 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.099 $X2=0.351 $Y2=0.126
r90 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.161 $Y=0.049 $X2=1.161
+ $Y2=0.049
r91 43 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.126
r92 38 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.9
+ $Y=0.081 $X2=0.936 $Y2=0.081
r93 37 64 8.08025 $w=1.8e-08 $l=1.19e-07 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.2
r94 37 51 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.049
r95 36 39 15.2778 $w=1.8e-08 $l=2.25e-07 $layer=M2 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=0.936 $Y2=0.081
r96 36 37 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.161 $Y=0.081 $X2=1.161
+ $Y2=0.081
r97 33 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.099
r98 32 38 37.2778 $w=1.8e-08 $l=5.49e-07 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.9 $Y2=0.081
r99 32 33 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.081 $X2=0.351
+ $Y2=0.081
r100 28 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.17
+ $Y=0.234 $X2=1.179 $Y2=0.234
r101 26 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.188
+ $Y=0.234 $X2=1.179 $Y2=0.234
r102 23 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.225 $X2=1.161 $Y2=0.2125
r103 22 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.17 $Y2=0.234
r104 22 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.161 $Y2=0.225
r105 17 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.188 $Y=0.234
+ $X2=1.188 $Y2=0.234
r106 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.2295 $X2=1.19 $Y2=0.2295
r107 12 50 16.2355 $w=3.7e-08 $l=2.9e-08 $layer=LISD $thickness=2.8e-08 $X=1.19
+ $Y=0.0455 $X2=1.161 $Y2=0.0455
r108 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.0405 $X2=1.19 $Y2=0.0405
r109 5 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r110 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r111 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%D 2 5 7 11 VSS
c18 11 VSS 0.00145113f $X=0.405 $Y=0.134
c19 5 VSS 0.00106786f $X=0.405 $Y=0.135
c20 2 VSS 0.0589243f $X=0.405 $Y=0.0675
r21 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%SI 2 7 11 14 VSS
c21 14 VSS 0.0032805f $X=0.475 $Y=0.135
c22 11 VSS 0.0035781f $X=0.473 $Y=0.135
c23 2 VSS 0.0640988f $X=0.459 $Y=0.0675
r24 11 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.475 $Y=0.135 $X2=0.475
+ $Y2=0.135
r25 5 14 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.475 $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%9 2 5 8 11 14 17 20 23 37 40 42 45 49 53 58 60 67
+ 69 74 78 80 96 101 102 103 104 106 VSS
c120 108 VSS 7.92414e-20 $X=0.189 $Y=0.207
c121 106 VSS 2.53862e-19 $X=0.189 $Y=0.178
c122 105 VSS 3.91706e-20 $X=0.189 $Y=0.167
c123 104 VSS 6.6467e-19 $X=0.189 $Y=0.164
c124 103 VSS 3.3761e-19 $X=0.189 $Y=0.144
c125 102 VSS 4.92067e-19 $X=0.189 $Y=0.121
c126 101 VSS 8.32677e-19 $X=0.189 $Y=0.099
c127 96 VSS 6.49238e-19 $X=0.729 $Y=0.18
c128 80 VSS 0.0152374f $X=0.729 $Y=0.189
c129 78 VSS 0.0013748f $X=0.567 $Y=0.189
c130 74 VSS 6.28429e-19 $X=0.189 $Y=0.189
c131 69 VSS 0.00386366f $X=0.18 $Y=0.234
c132 68 VSS 4.87314e-19 $X=0.189 $Y=0.225
c133 67 VSS 0.00199636f $X=0.189 $Y=0.234
c134 60 VSS 0.00373046f $X=0.18 $Y=0.036
c135 58 VSS 0.00194932f $X=0.189 $Y=0.036
c136 53 VSS 9.61695e-20 $X=0.567 $Y=0.18
c137 49 VSS 5.76385e-19 $X=0.567 $Y=0.135
c138 45 VSS 0.00566559f $X=0.16 $Y=0.216
c139 40 VSS 0.0055918f $X=0.16 $Y=0.054
c140 20 VSS 0.108004f $X=0.945 $Y=0.178
c141 17 VSS 1.08457e-19 $X=0.837 $Y=0.178
c142 14 VSS 0.060017f $X=0.837 $Y=0.0405
c143 11 VSS 2.24613e-19 $X=0.675 $Y=0.178
c144 8 VSS 0.0602569f $X=0.675 $Y=0.0405
c145 2 VSS 0.0660345f $X=0.567 $Y=0.1355
r146 107 108 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.2 $X2=0.189 $Y2=0.207
r147 105 106 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.167 $X2=0.189 $Y2=0.178
r148 104 105 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.167
r149 103 104 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.164
r150 102 103 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.121 $X2=0.189 $Y2=0.144
r151 101 102 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.099 $X2=0.189 $Y2=0.121
r152 95 96 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.729 $Y=0.18 $X2=0.729
+ $Y2=0.18
r153 80 96 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.729 $Y=0.189 $X2=0.729
+ $Y2=0.189
r154 77 80 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.729 $Y2=0.189
r155 77 78 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.567 $Y=0.189 $X2=0.567
+ $Y2=0.189
r156 74 107 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.2
r157 74 106 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.178
r158 73 77 25.6667 $w=1.8e-08 $l=3.78e-07 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.567 $Y2=0.189
r159 73 74 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.189 $X2=0.189
+ $Y2=0.189
r160 69 70 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r161 68 108 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.207
r162 67 70 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r163 67 68 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.189 $Y2=0.225
r164 64 69 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r165 60 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r166 59 101 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.099
r167 58 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r168 58 59 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r169 55 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r170 53 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.18 $X2=0.567 $Y2=0.189
r171 52 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.171 $X2=0.567 $Y2=0.18
r172 49 52 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.171
r173 45 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r174 42 45 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r175 40 55 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r176 37 40 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r177 20 23 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.178 $X2=0.945 $Y2=0.2295
r178 17 20 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08 $X=0.837
+ $Y=0.178 $X2=0.945 $Y2=0.178
r179 17 95 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08 $X=0.837
+ $Y=0.178 $X2=0.729 $Y2=0.178
r180 14 17 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0405 $X2=0.837 $Y2=0.178
r181 11 95 43.022 $w=2.6e-08 $l=5.4e-08 $layer=LISD $thickness=2.8e-08 $X=0.675
+ $Y=0.178 $X2=0.729 $Y2=0.178
r182 8 11 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.178
r183 2 49 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r184 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1355 $X2=0.567 $Y2=0.2025
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%10 2 7 9 10 13 14 17 19 22 27 28 29 31 33 38 40 46
+ 47 48 49 50 51 52 56 VSS
c49 58 VSS 5.19568e-19 $X=0.828 $Y=0.09
c50 57 VSS 3.9329e-19 $X=0.819 $Y=0.09
c51 56 VSS 4.29e-19 $X=0.837 $Y=0.09
c52 52 VSS 5.92866e-19 $X=0.837 $Y=0.207
c53 51 VSS 1.19762e-19 $X=0.837 $Y=0.167
c54 50 VSS 1.86299e-19 $X=0.837 $Y=0.165
c55 49 VSS 3.05662e-19 $X=0.837 $Y=0.14
c56 48 VSS 4.69487e-19 $X=0.837 $Y=0.122
c57 47 VSS 1.91116e-19 $X=0.837 $Y=0.101
c58 46 VSS 4.02479e-19 $X=0.837 $Y=0.225
c59 44 VSS 3.58124e-20 $X=0.81 $Y=0.0715
c60 40 VSS 0.00112276f $X=0.81 $Y=0.054
c61 33 VSS 0.00268883f $X=0.81 $Y=0.234
c62 31 VSS 0.00427376f $X=0.828 $Y=0.234
c63 30 VSS 2.64081e-19 $X=0.799 $Y=0.09
c64 29 VSS 0.00133552f $X=0.797 $Y=0.09
c65 28 VSS 0.00410211f $X=0.747 $Y=0.09
c66 27 VSS 4.49532e-19 $X=0.747 $Y=0.09
c67 24 VSS 4.45336e-20 $X=0.801 $Y=0.09
c68 22 VSS 0.0178238f $X=0.866 $Y=0.2295
c69 19 VSS 3.14771e-19 $X=0.881 $Y=0.2295
c70 17 VSS 2.5391e-19 $X=0.808 $Y=0.2295
c71 13 VSS 0.0201369f $X=0.81 $Y=0.0405
c72 9 VSS 6.29543e-19 $X=0.827 $Y=0.0405
c73 2 VSS 0.0580179f $X=0.729 $Y=0.0405
r74 57 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.819
+ $Y=0.09 $X2=0.828 $Y2=0.09
r75 56 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.09 $X2=0.828 $Y2=0.09
r76 55 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.09 $X2=0.819 $Y2=0.09
r77 51 52 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.167 $X2=0.837 $Y2=0.207
r78 50 51 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.165 $X2=0.837 $Y2=0.167
r79 49 50 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.14 $X2=0.837 $Y2=0.165
r80 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.122 $X2=0.837 $Y2=0.14
r81 47 48 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.101 $X2=0.837 $Y2=0.122
r82 46 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.207
r83 45 56 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.09
r84 45 47 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.101
r85 43 44 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.062 $X2=0.81 $Y2=0.0715
r86 40 43 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.054 $X2=0.81 $Y2=0.062
r87 38 55 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.09
r88 38 44 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.0715
r89 31 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r90 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.81 $Y2=0.234
r91 29 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.797
+ $Y=0.09 $X2=0.799 $Y2=0.09
r92 27 29 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.09 $X2=0.797 $Y2=0.09
r93 27 28 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.747 $Y=0.09 $X2=0.747
+ $Y2=0.09
r94 24 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.81 $Y2=0.09
r95 24 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.799 $Y2=0.09
r96 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2295 $X2=0.866 $Y2=0.2295
r97 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.808
+ $Y=0.2295 $X2=0.866 $Y2=0.2295
r98 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.234 $X2=0.81
+ $Y2=0.234
r99 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2295 $X2=0.808 $Y2=0.2295
r100 13 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.054 $X2=0.81
+ $Y2=0.054
r101 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.0405 $X2=0.81 $Y2=0.0405
r102 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.0405 $X2=0.81 $Y2=0.0405
r103 5 28 16.3636 $w=2.2e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.09 $X2=0.747 $Y2=0.09
r104 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.09 $X2=0.729 $Y2=0.2295
r105 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0405 $X2=0.729 $Y2=0.09
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%11 2 5 7 9 14 17 21 22 25 30 31 33 34 37 39 40 43
+ 44 45 46 48 50 51 52 53 54 55 56 59 61 62 65 VSS
c72 65 VSS 1.00162e-19 $X=0.693 $Y=0.131
c73 61 VSS 9.09188e-19 $X=0.72 $Y=0.131
c74 59 VSS 8.5526e-19 $X=0.783 $Y=0.131
c75 56 VSS 1.82087e-19 $X=0.693 $Y=0.216
c76 55 VSS 1.40959e-19 $X=0.693 $Y=0.207
c77 54 VSS 1.07888e-19 $X=0.693 $Y=0.189
c78 53 VSS 1.66071e-19 $X=0.693 $Y=0.171
c79 52 VSS 2.71272e-19 $X=0.693 $Y=0.165
c80 51 VSS 3.53682e-19 $X=0.693 $Y=0.153
c81 50 VSS 2.11704e-19 $X=0.693 $Y=0.225
c82 48 VSS 4.15228e-19 $X=0.693 $Y=0.114
c83 47 VSS 2.7378e-19 $X=0.693 $Y=0.106
c84 46 VSS 5.46003e-20 $X=0.693 $Y=0.099
c85 45 VSS 5.96385e-20 $X=0.693 $Y=0.081
c86 43 VSS 1.65771e-19 $X=0.693 $Y=0.062
c87 42 VSS 2.30403e-19 $X=0.693 $Y=0.122
c88 40 VSS 0.00145015f $X=0.6665 $Y=0.036
c89 39 VSS 0.00201121f $X=0.649 $Y=0.036
c90 37 VSS 0.00303728f $X=0.648 $Y=0.036
c91 34 VSS 0.00412969f $X=0.684 $Y=0.036
c92 33 VSS 0.00297725f $X=0.649 $Y=0.234
c93 32 VSS 2.2805e-19 $X=0.612 $Y=0.234
c94 31 VSS 0.00126734f $X=0.609 $Y=0.234
c95 30 VSS 0.0016591f $X=0.595 $Y=0.234
c96 25 VSS 0.00558865f $X=0.684 $Y=0.234
c97 24 VSS 5.62656e-19 $X=0.594 $Y=0.2295
c98 21 VSS 0.00254121f $X=0.594 $Y=0.2025
c99 18 VSS 1.02475e-19 $X=0.5895 $Y=0.216
c100 16 VSS 5.70081e-19 $X=0.648 $Y=0.0405
c101 10 VSS 7.61325e-20 $X=0.6435 $Y=0.054
c102 5 VSS 0.00231049f $X=0.783 $Y=0.131
c103 2 VSS 0.0591968f $X=0.783 $Y=0.0405
r104 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.131 $X2=0.738 $Y2=0.131
r105 59 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.131 $X2=0.738 $Y2=0.131
r106 57 65 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.693 $Y2=0.131
r107 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.72 $Y2=0.131
r108 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.207 $X2=0.693 $Y2=0.216
r109 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.189 $X2=0.693 $Y2=0.207
r110 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.171 $X2=0.693 $Y2=0.189
r111 52 53 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.165 $X2=0.693 $Y2=0.171
r112 51 52 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.153 $X2=0.693 $Y2=0.165
r113 50 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.225 $X2=0.693 $Y2=0.216
r114 49 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.131
r115 49 51 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.153
r116 47 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.106 $X2=0.693 $Y2=0.114
r117 46 47 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.099 $X2=0.693 $Y2=0.106
r118 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.081 $X2=0.693 $Y2=0.099
r119 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.063 $X2=0.693 $Y2=0.081
r120 43 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.062 $X2=0.693 $Y2=0.063
r121 42 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.131
r122 42 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.114
r123 41 43 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.045 $X2=0.693 $Y2=0.062
r124 39 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.649
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r125 36 39 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.649 $Y2=0.036
r126 36 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r127 34 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.036 $X2=0.693 $Y2=0.045
r128 34 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r129 32 33 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.649 $Y2=0.234
r130 31 32 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.609
+ $Y=0.234 $X2=0.612 $Y2=0.234
r131 30 31 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.595
+ $Y=0.234 $X2=0.609 $Y2=0.234
r132 27 30 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.595 $Y2=0.234
r133 25 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.234 $X2=0.693 $Y2=0.225
r134 25 33 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.234 $X2=0.649 $Y2=0.234
r135 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2295 $X2=0.594 $Y2=0.2295
r136 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r137 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.594 $Y2=0.2295
r138 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.5895 $Y2=0.189
r139 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.189 $X2=0.5895 $Y2=0.189
r140 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r141 13 37 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r142 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.648 $Y2=0.0405
r143 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.6435 $Y2=0.081
r144 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.081 $X2=0.6435 $Y2=0.081
r145 5 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.131 $X2=0.783
+ $Y2=0.131
r146 5 7 369.03 $w=2e-08 $l=9.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.131 $X2=0.783 $Y2=0.2295
r147 2 5 339.058 $w=2e-08 $l=9.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.131
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%12 2 5 7 9 12 14 17 21 25 26 30 31 35 36 37 43 VSS
c33 43 VSS 0.00419842f $X=1.098 $Y=0.234
c34 42 VSS 0.00204425f $X=1.107 $Y=0.234
c35 37 VSS 0.00106194f $X=1.107 $Y=0.171
c36 36 VSS 0.00114954f $X=1.107 $Y=0.117
c37 35 VSS 0.00158518f $X=1.107 $Y=0.225
c38 33 VSS 7.70286e-19 $X=1.073 $Y=0.036
c39 32 VSS 4.41014e-19 $X=1.066 $Y=0.036
c40 31 VSS 0.00146362f $X=1.062 $Y=0.036
c41 30 VSS 0.00481311f $X=1.044 $Y=0.036
c42 26 VSS 0.00226308f $X=1.008 $Y=0.036
c43 25 VSS 0.00460331f $X=1.098 $Y=0.036
c44 21 VSS 7.16657e-19 $X=0.999 $Y=0.105
c45 17 VSS 0.00426839f $X=1.078 $Y=0.2295
c46 12 VSS 0.00485453f $X=1.078 $Y=0.0405
c47 5 VSS 0.00233254f $X=0.999 $Y=0.1055
c48 2 VSS 0.0590816f $X=0.999 $Y=0.0405
r49 43 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r50 42 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r51 39 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.098 $Y2=0.234
r52 36 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.117 $X2=1.107 $Y2=0.171
r53 35 42 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.234
r54 35 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.171
r55 34 36 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.045 $X2=1.107 $Y2=0.117
r56 32 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.066
+ $Y=0.036 $X2=1.073 $Y2=0.036
r57 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=1.062
+ $Y=0.036 $X2=1.066 $Y2=0.036
r58 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=1.062 $Y2=0.036
r59 28 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.036 $X2=1.073 $Y2=0.036
r60 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.008
+ $Y=0.036 $X2=1.044 $Y2=0.036
r61 25 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.098 $Y=0.036 $X2=1.107 $Y2=0.045
r62 25 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.036 $X2=1.08 $Y2=0.036
r63 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.999 $Y=0.045 $X2=1.008 $Y2=0.036
r64 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.045 $X2=0.999 $Y2=0.105
r65 17 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234 $X2=1.08
+ $Y2=0.234
r66 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2295 $X2=1.078 $Y2=0.2295
r67 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.036 $X2=1.08
+ $Y2=0.036
r68 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.0405 $X2=1.078 $Y2=0.0405
r69 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.105 $X2=0.999
+ $Y2=0.105
r70 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.1055 $X2=0.999 $Y2=0.2295
r71 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.0405 $X2=0.999 $Y2=0.1055
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%13 2 7 10 13 15 17 18 21 22 23 26 27 32 33 35 38
+ 39 40 41 43 46 47 50 60 65 68 70 71 78 VSS
c70 78 VSS 0.00312516f $X=1.269 $Y=0.136
c71 71 VSS 0.00160638f $X=1.229 $Y=0.153
c72 70 VSS 0.00791219f $X=1.175 $Y=0.153
c73 68 VSS 0.00415759f $X=1.269 $Y=0.153
c74 65 VSS 1.90597e-19 $X=0.945 $Y=0.153
c75 60 VSS 0.0033916f $X=0.936 $Y=0.234
c76 59 VSS 0.00253671f $X=0.945 $Y=0.234
c77 50 VSS 4.04001e-19 $X=1.053 $Y=0.14
c78 47 VSS 3.26354e-19 $X=1.008 $Y=0.162
c79 46 VSS 0.00199114f $X=0.99 $Y=0.162
c80 44 VSS 0.0023929f $X=1.044 $Y=0.162
c81 43 VSS 0.00104404f $X=0.945 $Y=0.225
c82 41 VSS 2.07499e-19 $X=0.945 $Y=0.136
c83 40 VSS 2.77769e-19 $X=0.945 $Y=0.119
c84 39 VSS 2.61356e-19 $X=0.945 $Y=0.101
c85 38 VSS 6.393e-19 $X=0.945 $Y=0.081
c86 37 VSS 3.04212e-19 $X=0.945 $Y=0.153
c87 35 VSS 0.00136569f $X=0.92 $Y=0.036
c88 34 VSS 4.8751e-19 $X=0.904 $Y=0.036
c89 33 VSS 0.00146362f $X=0.9 $Y=0.036
c90 32 VSS 0.00358427f $X=0.882 $Y=0.036
c91 27 VSS 0.00347893f $X=0.936 $Y=0.036
c92 26 VSS 0.00276615f $X=0.918 $Y=0.2295
c93 22 VSS 5.63046e-19 $X=0.935 $Y=0.2295
c94 21 VSS 0.0201056f $X=0.864 $Y=0.0405
c95 17 VSS 5.63046e-19 $X=0.881 $Y=0.0405
c96 13 VSS 0.00278011f $X=1.269 $Y=0.136
c97 10 VSS 0.0625639f $X=1.269 $Y=0.0675
c98 5 VSS 0.00302777f $X=1.053 $Y=0.14
c99 2 VSS 0.0627731f $X=1.053 $Y=0.0405
r100 70 71 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=1.175
+ $Y=0.153 $X2=1.229 $Y2=0.153
r101 68 71 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.269
+ $Y=0.153 $X2=1.229 $Y2=0.153
r102 68 78 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.269 $Y=0.153 $X2=1.269
+ $Y2=0.153
r103 64 70 15.6173 $w=1.8e-08 $l=2.3e-07 $layer=M2 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=1.175 $Y2=0.153
r104 64 65 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.945 $Y=0.153 $X2=0.945
+ $Y2=0.153
r105 60 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r106 59 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r107 56 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.234 $X2=0.936 $Y2=0.234
r108 48 50 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.153 $X2=1.053 $Y2=0.14
r109 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.99
+ $Y=0.162 $X2=1.008 $Y2=0.162
r110 45 65 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.945 $Y2=0.162
r111 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.99 $Y2=0.162
r112 44 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.162 $X2=1.053 $Y2=0.153
r113 44 47 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.162 $X2=1.008 $Y2=0.162
r114 43 59 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.234
r115 42 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.162
r116 42 43 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.225
r117 40 41 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.119 $X2=0.945 $Y2=0.136
r118 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.101 $X2=0.945 $Y2=0.119
r119 38 39 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.081 $X2=0.945 $Y2=0.101
r120 37 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.162
r121 37 41 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.136
r122 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.081
r123 34 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.904
+ $Y=0.036 $X2=0.92 $Y2=0.036
r124 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.036 $X2=0.904 $Y2=0.036
r125 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r126 29 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r127 27 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r128 27 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.92 $Y2=0.036
r129 26 56 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.234
+ $X2=0.918 $Y2=0.234
r130 23 26 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.2295 $X2=0.918 $Y2=0.2295
r131 22 26 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.935 $Y=0.2295 $X2=0.918 $Y2=0.2295
r132 21 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036
+ $X2=0.864 $Y2=0.036
r133 18 21 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.864 $Y2=0.0405
r134 17 21 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0405 $X2=0.864 $Y2=0.0405
r135 13 78 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.269 $Y=0.136 $X2=1.269
+ $Y2=0.136
r136 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.136 $X2=1.269 $Y2=0.2025
r137 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.0675 $X2=1.269 $Y2=0.136
r138 5 50 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.053 $Y=0.14 $X2=1.053
+ $Y2=0.14
r139 5 7 335.312 $w=2e-08 $l=8.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.14 $X2=1.053 $Y2=0.2295
r140 2 5 372.777 $w=2e-08 $l=9.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.0405 $X2=1.053 $Y2=0.14
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%14 1 4 6 11 14 21 23 24 25 VSS
c29 26 VSS 0.00225803f $X=0.485 $Y=0.234
c30 25 VSS 0.0014167f $X=0.461 $Y=0.234
c31 24 VSS 0.0134342f $X=0.447 $Y=0.234
c32 23 VSS 0.00523898f $X=0.309 $Y=0.234
c33 21 VSS 0.00168783f $X=0.486 $Y=0.234
c34 14 VSS 0.0195485f $X=0.542 $Y=0.2025
c35 11 VSS 3.25039e-19 $X=0.557 $Y=0.2025
c36 9 VSS 4.57278e-19 $X=0.484 $Y=0.2025
c37 4 VSS 0.00250857f $X=0.272 $Y=0.2025
c38 1 VSS 3.31752e-19 $X=0.287 $Y=0.2025
r39 25 26 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.461
+ $Y=0.234 $X2=0.485 $Y2=0.234
r40 24 25 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.234 $X2=0.461 $Y2=0.234
r41 23 24 9.37037 $w=1.8e-08 $l=1.38e-07 $layer=M1 $thickness=3.6e-08 $X=0.309
+ $Y=0.234 $X2=0.447 $Y2=0.234
r42 21 26 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.485 $Y2=0.234
r43 17 23 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.309 $Y2=0.234
r44 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.542 $Y2=0.2025
r45 9 14 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.484
+ $Y=0.2025 $X2=0.542 $Y2=0.2025
r46 9 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r47 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.2025 $X2=0.484 $Y2=0.2025
r48 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r49 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.272 $Y2=0.2025
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%16 1 2 5 6 7 10 12 18 20 21 22 23 24 25 VSS
c21 25 VSS 3.8923e-20 $X=0.423 $Y=0.198
c22 24 VSS 8.46035e-21 $X=0.414 $Y=0.198
c23 23 VSS 0.00116854f $X=0.396 $Y=0.198
c24 22 VSS 0.00134991f $X=0.379 $Y=0.198
c25 21 VSS 8.46035e-21 $X=0.36 $Y=0.198
c26 20 VSS 2.61077e-19 $X=0.342 $Y=0.198
c27 18 VSS 3.31089e-19 $X=0.432 $Y=0.198
c28 12 VSS 5.44897e-19 $X=0.324 $Y=0.198
c29 10 VSS 0.00631853f $X=0.432 $Y=0.2025
c30 6 VSS 5.67296e-19 $X=0.449 $Y=0.2025
c31 5 VSS 0.00790786f $X=0.324 $Y=0.2025
c32 1 VSS 6.05629e-19 $X=0.341 $Y=0.2025
r33 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.423 $Y2=0.198
r34 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.414 $Y2=0.198
r35 22 23 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.198 $X2=0.396 $Y2=0.198
r36 21 22 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.198 $X2=0.379 $Y2=0.198
r37 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r38 18 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.423 $Y2=0.198
r39 12 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.342 $Y2=0.198
r40 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r41 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r42 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r43 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198 $X2=0.324
+ $Y2=0.198
r44 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
r45 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%QN 1 6 9 14 15 16 19 22 30 VSS
c7 30 VSS 0.0042609f $X=1.314 $Y=0.234
c8 29 VSS 0.00278493f $X=1.323 $Y=0.234
c9 22 VSS 0.00408512f $X=1.314 $Y=0.036
c10 21 VSS 0.00278493f $X=1.323 $Y=0.036
c11 19 VSS 0.00664444f $X=1.296 $Y=0.036
c12 16 VSS 0.00487569f $X=1.323 $Y=0.2
c13 15 VSS 0.00226847f $X=1.323 $Y=0.09
c14 12 VSS 0.0013947f $X=1.323 $Y=0.225
c15 9 VSS 0.00691625f $X=1.294 $Y=0.2025
c16 4 VSS 3.77696e-19 $X=1.294 $Y=0.0675
r17 30 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.314
+ $Y=0.234 $X2=1.3185 $Y2=0.234
r18 29 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.234 $X2=1.3185 $Y2=0.234
r19 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.234 $X2=1.314 $Y2=0.234
r20 22 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.314
+ $Y=0.036 $X2=1.3185 $Y2=0.036
r21 21 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.036 $X2=1.3185 $Y2=0.036
r22 18 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.036 $X2=1.314 $Y2=0.036
r23 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.036 $X2=1.296
+ $Y2=0.036
r24 15 16 7.46914 $w=1.8e-08 $l=1.1e-07 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.09 $X2=1.323 $Y2=0.2
r25 14 16 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.223 $X2=1.323 $Y2=0.2
r26 12 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.225 $X2=1.323 $Y2=0.234
r27 12 14 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.225 $X2=1.323 $Y2=0.223
r28 11 21 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.045 $X2=1.323 $Y2=0.036
r29 11 15 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.045 $X2=1.323 $Y2=0.09
r30 9 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.234 $X2=1.296
+ $Y2=0.234
r31 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=1.279
+ $Y=0.2025 $X2=1.294 $Y2=0.2025
r32 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.296
+ $Y=0.0675 $X2=1.296 $Y2=0.036
r33 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.279
+ $Y=0.0675 $X2=1.294 $Y2=0.0675
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%19 1 6 9 VSS
c10 9 VSS 0.0140217f $X=0.704 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.719 $Y=0.2295
c12 4 VSS 2.70811e-19 $X=0.646 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.646
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.631
+ $Y=0.2295 $X2=0.646 $Y2=0.2295
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%20 1 6 9 VSS
c9 9 VSS 0.0145746f $X=0.974 $Y=0.0405
c10 6 VSS 3.14771e-19 $X=0.989 $Y=0.0405
c11 4 VSS 2.65708e-19 $X=0.916 $Y=0.0405
r12 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r13 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.916
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r14 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.901
+ $Y=0.0405 $X2=0.916 $Y2=0.0405
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%22 1 2 VSS
c2 1 VSS 0.00203573f $X=0.719 $Y=0.0405
r3 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0405 $X2=0.685 $Y2=0.0405
.ends

.subckt PM_SDFHX1_ASAP7_75T_SRAM%23 1 2 VSS
c0 1 VSS 0.00214045f $X=0.989 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.2295 $X2=0.955 $Y2=0.2295
.ends


* END of "./SDFHx1_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt SDFHx1_ASAP7_75t_SRAM  VSS VDD CLK SE D SI QN
* 
* QN	QN
* SI	SI
* D	D
* SE	SE
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_9_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_SE_M2_g noxref_15 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 noxref_21 N_6_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 noxref_17 N_D_M4_g noxref_21 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 noxref_15 N_SI_M5_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 N_11_M6_d N_4_M6_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M7 N_22_M7_d N_9_M7_g N_11_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M8 VSS N_10_M8_g N_22_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.027
M9 N_10_M9_d N_11_M9_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_13_M10_d N_9_M10_g N_10_M10_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.827 $Y=0.027
M11 N_20_M11_d N_4_M11_g N_13_M11_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.027
M12 VSS N_12_M12_g N_20_M12_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.027
M13 N_12_M13_d N_13_M13_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.027
M14 VSS N_SE_M14_g N_6_M14_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.205
+ $Y=0.027
M15 N_QN_M15_d N_13_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M16 VDD N_CLK_M16_g N_4_M16_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M17 N_9_M17_d N_4_M17_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M18 N_16_M18_d N_SE_M18_g N_14_M18_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M19 VDD N_6_M19_g N_16_M19_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M20 N_16_M20_d N_D_M20_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M21 N_14_M21_d N_SI_M21_g N_16_M21_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M22 N_11_M22_d N_9_M22_g N_14_M22_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M23 N_19_M23_d N_4_M23_g N_11_M23_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.611 $Y=0.216
M24 VDD N_10_M24_g N_19_M24_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.216
M25 N_10_M25_d N_11_M25_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M26 N_13_M26_d N_4_M26_g N_10_M26_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.216
M27 N_23_M27_d N_9_M27_g N_13_M27_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.935 $Y=0.216
M28 VDD N_12_M28_g N_23_M28_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.216
M29 N_12_M29_d N_13_M29_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.216
M30 VDD N_SE_M30_g N_6_M30_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.205
+ $Y=0.216
M31 N_QN_M31_d N_13_M31_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
*
* 
* .include "SDFHx1_ASAP7_75t_SRAM.pex.sp.SDFHX1_ASAP7_75T_SRAM.pxi"
* BEGIN of "./SDFHx1_ASAP7_75t_SRAM.pex.sp.SDFHX1_ASAP7_75T_SRAM.pxi"
* File: SDFHx1_ASAP7_75t_SRAM.pex.sp.SDFHX1_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 13:03:02 2017
* 
x_PM_SDFHX1_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M16_g N_CLK_c_3_p CLK
+ N_CLK_c_9_p N_CLK_c_7_p N_CLK_c_19_p VSS PM_SDFHX1_ASAP7_75T_SRAM%CLK
x_PM_SDFHX1_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_21_n N_4_M17_g N_4_M6_g N_4_c_41_p
+ N_4_M23_g N_4_M11_g N_4_c_45_p N_4_M26_g N_4_M0_s N_4_c_22_n N_4_M16_s
+ N_4_c_23_n N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_54_p N_4_c_35_p
+ N_4_c_28_n N_4_c_58_p N_4_c_29_n N_4_c_56_p N_4_c_32_p N_4_c_36_p N_4_c_46_p
+ N_4_c_34_p N_4_c_65_p N_4_c_31_n N_4_c_48_p VSS PM_SDFHX1_ASAP7_75T_SRAM%4
x_PM_SDFHX1_ASAP7_75T_SRAM%SE N_SE_M2_g N_SE_c_91_p N_SE_M18_g N_SE_M14_g
+ N_SE_c_126_p N_SE_M30_g N_SE_c_96_p N_SE_c_140_p N_SE_c_138_p N_SE_c_156_p
+ N_SE_c_87_n SE N_SE_c_86_n N_SE_c_92_p N_SE_c_93_p N_SE_c_88_n N_SE_c_89_n
+ N_SE_c_136_p N_SE_c_105_p N_SE_c_109_p N_SE_c_94_p N_SE_c_137_p VSS
+ PM_SDFHX1_ASAP7_75T_SRAM%SE
x_PM_SDFHX1_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_169_n N_6_M19_g N_6_M14_s N_6_c_170_n
+ N_6_M30_s N_6_c_199_p N_6_c_206_p N_6_c_216_p N_6_c_203_p N_6_c_212_p
+ N_6_c_220_p N_6_c_172_n N_6_c_165_n N_6_c_187_p N_6_c_167_n N_6_c_175_n
+ N_6_c_178_n N_6_c_179_n N_6_c_205_p VSS PM_SDFHX1_ASAP7_75T_SRAM%6
x_PM_SDFHX1_ASAP7_75T_SRAM%D N_D_M4_g N_D_c_237_n N_D_M20_g D VSS
+ PM_SDFHX1_ASAP7_75T_SRAM%D
x_PM_SDFHX1_ASAP7_75T_SRAM%SI N_SI_M5_g N_SI_M21_g SI N_SI_c_257_n VSS
+ PM_SDFHX1_ASAP7_75T_SRAM%SI
x_PM_SDFHX1_ASAP7_75T_SRAM%9 N_9_c_279_n N_9_M22_g N_9_M7_g N_9_c_346_p N_9_M10_g
+ N_9_c_330_p N_9_c_283_n N_9_M27_g N_9_M1_d N_9_c_288_n N_9_M17_d N_9_c_289_n
+ N_9_c_290_n N_9_c_315_n N_9_c_302_n N_9_c_273_n N_9_c_374_p N_9_c_293_n
+ N_9_c_274_n N_9_c_296_n N_9_c_275_n N_9_c_299_n N_9_c_276_n N_9_c_277_n
+ N_9_c_300_n N_9_c_301_n N_9_c_278_n VSS PM_SDFHX1_ASAP7_75T_SRAM%9
x_PM_SDFHX1_ASAP7_75T_SRAM%10 N_10_M8_g N_10_M24_g N_10_M10_s N_10_M9_d
+ N_10_c_398_n N_10_M25_d N_10_c_411_n N_10_M26_s N_10_c_413_n N_10_c_401_n
+ N_10_c_402_n N_10_c_399_n N_10_c_440_p N_10_c_394_n N_10_c_404_n N_10_c_400_n
+ N_10_c_427_p N_10_c_441_p N_10_c_396_n N_10_c_429_p N_10_c_397_n N_10_c_417_n
+ N_10_c_418_n N_10_c_405_n VSS PM_SDFHX1_ASAP7_75T_SRAM%10
x_PM_SDFHX1_ASAP7_75T_SRAM%11 N_11_M9_g N_11_c_443_n N_11_M25_g N_11_M6_d N_11_M7_s
+ N_11_M22_d N_11_c_444_n N_11_M23_s N_11_c_507_p N_11_c_466_n N_11_c_467_n
+ N_11_c_445_n N_11_c_453_n N_11_c_454_n N_11_c_455_n N_11_c_456_n N_11_c_457_n
+ N_11_c_490_n N_11_c_459_n N_11_c_460_n N_11_c_447_n N_11_c_510_p N_11_c_448_n
+ N_11_c_449_n N_11_c_472_n N_11_c_474_n N_11_c_477_n N_11_c_511_p N_11_c_451_n
+ N_11_c_452_n N_11_c_484_n N_11_c_486_n VSS PM_SDFHX1_ASAP7_75T_SRAM%11
x_PM_SDFHX1_ASAP7_75T_SRAM%12 N_12_M12_g N_12_c_536_p N_12_M28_g N_12_M13_d
+ N_12_c_521_n N_12_M29_d N_12_c_523_n N_12_c_515_n N_12_c_516_n N_12_c_517_n
+ N_12_c_518_n N_12_c_519_n N_12_c_527_n N_12_c_520_n N_12_c_530_n N_12_c_545_p
+ VSS PM_SDFHX1_ASAP7_75T_SRAM%12
x_PM_SDFHX1_ASAP7_75T_SRAM%13 N_13_M13_g N_13_M29_g N_13_M15_g N_13_c_553_n
+ N_13_M31_g N_13_M11_s N_13_M10_d N_13_c_554_n N_13_M27_s N_13_M26_d
+ N_13_c_578_n N_13_c_555_n N_13_c_556_n N_13_c_547_n N_13_c_558_n N_13_c_559_n
+ N_13_c_567_n N_13_c_549_n N_13_c_580_n N_13_c_581_n N_13_c_616_p N_13_c_601_n
+ N_13_c_603_n N_13_c_568_n N_13_c_550_n N_13_c_560_n N_13_c_551_n N_13_c_562_n
+ N_13_c_564_n VSS PM_SDFHX1_ASAP7_75T_SRAM%13
x_PM_SDFHX1_ASAP7_75T_SRAM%14 N_14_M18_s N_14_c_618_n N_14_M21_d N_14_M22_s
+ N_14_c_617_n N_14_c_624_n N_14_c_619_n N_14_c_621_n N_14_c_625_n VSS
+ PM_SDFHX1_ASAP7_75T_SRAM%14
x_PM_SDFHX1_ASAP7_75T_SRAM%16 N_16_M19_s N_16_M18_d N_16_c_660_n N_16_M21_s
+ N_16_M20_d N_16_c_662_n N_16_c_652_n N_16_c_651_n N_16_c_654_n N_16_c_646_n
+ N_16_c_656_n N_16_c_657_n N_16_c_648_n N_16_c_650_n VSS
+ PM_SDFHX1_ASAP7_75T_SRAM%16
x_PM_SDFHX1_ASAP7_75T_SRAM%QN N_QN_M15_d N_QN_M31_d N_QN_c_670_n QN N_QN_c_667_n
+ N_QN_c_671_n N_QN_c_673_n N_QN_c_668_n N_QN_c_669_n VSS
+ PM_SDFHX1_ASAP7_75T_SRAM%QN
x_PM_SDFHX1_ASAP7_75T_SRAM%19 N_19_M23_d N_19_M24_s N_19_c_675_n VSS
+ PM_SDFHX1_ASAP7_75T_SRAM%19
x_PM_SDFHX1_ASAP7_75T_SRAM%20 N_20_M11_d N_20_M12_s N_20_c_684_n VSS
+ PM_SDFHX1_ASAP7_75T_SRAM%20
x_PM_SDFHX1_ASAP7_75T_SRAM%22 N_22_M8_s N_22_M7_d VSS PM_SDFHX1_ASAP7_75T_SRAM%22
x_PM_SDFHX1_ASAP7_75T_SRAM%23 N_23_M28_s N_23_M27_d VSS PM_SDFHX1_ASAP7_75T_SRAM%23
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_CLK_c_2_p N_4_c_21_n 0.00105598f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_CLK_c_3_p N_4_c_22_n 2.66516e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.054
cc_4 N_CLK_c_3_p N_4_c_23_n 0.0012473f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.144
cc_5 N_CLK_c_3_p N_4_c_24_n 3.97017e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.081
cc_6 N_CLK_c_3_p N_4_c_25_n 0.0012473f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.1125
cc_7 N_CLK_c_7_p N_4_c_26_n 0.00140648f $X=0.081 $Y=0.167 $X2=0.018 $Y2=0.2
cc_8 N_CLK_c_3_p N_4_c_27_n 4.97741e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_9_p N_4_c_28_n 0.00123168f $X=0.081 $Y=0.162 $X2=0.033 $Y2=0.153
cc_10 N_CLK_c_3_p N_4_c_29_n 5.36602e-19 $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_11 N_CLK_c_9_p N_4_c_29_n 8.66987e-19 $X=0.081 $Y=0.162 $X2=0.175 $Y2=0.153
cc_12 N_CLK_c_3_p N_4_c_31_n 0.00203815f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_13 N_CLK_c_3_p N_SE_c_86_n 2.45198e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2
cc_14 N_CLK_c_3_p N_9_c_273_n 6.32319e-19 $X=0.081 $Y=0.135 $X2=0.621 $Y2=0.135
cc_15 CLK N_9_c_274_n 3.23206e-19 $X=0.078 $Y=0.19 $X2=0.337 $Y2=0.153
cc_16 CLK N_9_c_275_n 2.57347e-19 $X=0.078 $Y=0.19 $X2=0.817 $Y2=0.153
cc_17 N_CLK_c_3_p N_9_c_276_n 0.00114506f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_18 N_CLK_c_3_p N_9_c_277_n 3.05593e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_19 N_CLK_c_19_p N_9_c_278_n 3.05593e-19 $X=0.081 $Y=0.1785 $X2=0 $Y2=0
cc_20 N_4_c_32_p N_SE_c_87_n 8.13669e-19 $X=0.337 $Y=0.153 $X2=0 $Y2=0
cc_21 N_4_c_32_p N_SE_c_88_n 0.00228328f $X=0.337 $Y=0.153 $X2=0 $Y2=0
cc_22 N_4_c_34_p N_SE_c_89_n 0.00228328f $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_23 N_4_c_35_p N_6_c_165_n 3.98881e-19 $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_24 N_4_c_36_p N_6_c_165_n 0.0176013f $X=0.479 $Y=0.153 $X2=0 $Y2=0
cc_25 N_4_c_36_p N_6_c_167_n 0.00114531f $X=0.479 $Y=0.153 $X2=0 $Y2=0
cc_26 N_4_c_36_p D 0.00102191f $X=0.479 $Y=0.153 $X2=0.081 $Y2=0.135
cc_27 N_4_c_34_p SI 0.00113575f $X=0.743 $Y=0.153 $X2=0.081 $Y2=0.135
cc_28 N_4_M6_g N_9_c_279_n 0.00365763f $X=0.621 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_29 N_4_c_41_p N_9_c_279_n 9.97803e-19 $X=0.621 $Y=0.135 $X2=0.081 $Y2=0.054
cc_30 N_4_M6_g N_9_M7_g 0.00355599f $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_4_M11_g N_9_M10_g 0.00355599f $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_32 N_4_M11_g N_9_c_283_n 0.00605856f $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.1785
cc_33 N_4_c_45_p N_9_c_283_n 0.00180656f $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.1785
cc_34 N_4_c_46_p N_9_c_283_n 5.51712e-19 $X=0.891 $Y=0.153 $X2=0.081 $Y2=0.1785
cc_35 N_4_c_34_p N_9_c_283_n 0.00168667f $X=0.743 $Y=0.153 $X2=0.081 $Y2=0.1785
cc_36 N_4_c_48_p N_9_c_283_n 0.00123876f $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.1785
cc_37 N_4_c_29_n N_9_c_288_n 2.18034e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_38 N_4_c_29_n N_9_c_289_n 2.58357e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_35_p N_9_c_290_n 0.00279251f $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_34_p N_9_c_290_n 9.87747e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_41 N_4_c_29_n N_9_c_273_n 3.93085e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_42 N_4_c_54_p N_9_c_293_n 2.66501e-19 $X=0.054 $Y=0.234 $X2=0 $Y2=0
cc_43 N_4_c_29_n N_9_c_293_n 4.19323e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_44 N_4_c_56_p N_9_c_274_n 2.46239e-19 $X=0.211 $Y=0.153 $X2=0 $Y2=0
cc_45 N_4_c_34_p N_9_c_296_n 2.46239e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_46 N_4_c_58_p N_9_c_275_n 3.80004e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_56_p N_9_c_275_n 0.0471484f $X=0.211 $Y=0.153 $X2=0 $Y2=0
cc_48 N_4_c_34_p N_9_c_299_n 2.81643e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_49 N_4_c_31_n N_9_c_300_n 0.00218805f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_50 N_4_c_56_p N_9_c_301_n 0.00116576f $X=0.211 $Y=0.153 $X2=0 $Y2=0
cc_51 N_4_M6_g N_10_M8_g 2.82885e-19 $X=0.621 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_52 N_4_c_46_p N_10_c_394_n 2.61213e-19 $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_53 N_4_c_65_p N_10_c_394_n 2.61213e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_54 N_4_c_48_p N_10_c_396_n 0.00318254f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_55 N_4_c_46_p N_10_c_397_n 0.00128311f $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_56 N_4_M11_g N_11_M9_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_57 N_4_c_45_p N_11_c_443_n 3.1781e-19 $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.135
cc_58 N_4_c_58_p N_11_c_444_n 3.24488e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_59 N_4_M6_g N_11_c_445_n 3.41974e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_60 N_4_c_58_p N_11_c_445_n 0.00102727f $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_61 N_4_c_35_p N_11_c_447_n 0.00133858f $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_62 N_4_c_34_p N_11_c_448_n 7.726e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_63 N_4_c_58_p N_11_c_449_n 8.63476e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_64 N_4_c_34_p N_11_c_449_n 5.92766e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_65 N_4_c_65_p N_11_c_451_n 3.86765e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_66 N_4_c_34_p N_11_c_452_n 3.86765e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_67 N_4_M11_g N_12_M12_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_68 N_4_M11_g N_13_c_547_n 3.18506e-19 $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_69 N_4_c_48_p N_13_c_547_n 4.09234e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_70 N_4_c_48_p N_13_c_549_n 0.00320381f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_71 N_4_c_48_p N_13_c_550_n 3.56772e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_72 N_4_c_46_p N_13_c_551_n 9.47997e-19 $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_73 N_4_c_36_p N_14_c_617_n 4.23942e-19 $X=0.479 $Y=0.153 $X2=0 $Y2=0
cc_74 N_SE_M2_g N_6_M3_g 0.00304756f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_75 N_SE_c_91_p N_6_c_169_n 0.00126421f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_76 N_SE_c_92_p N_6_c_170_n 2.11282e-19 $X=1.215 $Y=0.045 $X2=0.081 $Y2=0.135
cc_77 N_SE_c_93_p N_6_c_170_n 8.20809e-19 $X=1.215 $Y=0.045 $X2=0.081 $Y2=0.135
cc_78 N_SE_c_94_p N_6_c_172_n 3.53759e-19 $X=1.215 $Y=0.09 $X2=0 $Y2=0
cc_79 N_SE_c_89_n N_6_c_165_n 0.0680793f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_80 N_SE_c_96_p N_6_c_167_n 8.79603e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_81 N_SE_c_93_p N_6_c_175_n 0.00733801f $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_82 N_SE_c_89_n N_6_c_175_n 0.00103045f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_83 N_SE_c_94_p N_6_c_175_n 3.73635e-19 $X=1.215 $Y=0.09 $X2=0 $Y2=0
cc_84 N_SE_c_89_n N_6_c_178_n 2.46239e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_85 N_SE_c_87_n N_6_c_179_n 3.24594e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_86 N_SE_M2_g N_D_M4_g 2.13359e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_87 N_SE_c_86_n N_9_c_302_n 0.00266639f $X=0.225 $Y=0.045 $X2=0 $Y2=0
cc_88 N_SE_c_88_n N_9_c_302_n 4.45368e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_89 N_SE_c_105_p N_9_c_302_n 2.64176e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_90 N_SE_c_87_n N_9_c_275_n 4.53301e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_91 N_SE_c_88_n N_9_c_275_n 3.907e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_92 N_SE_c_105_p N_9_c_276_n 0.00292661f $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_93 N_SE_c_109_p N_9_c_277_n 0.00266639f $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_94 N_SE_c_87_n N_9_c_300_n 0.00266639f $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_95 N_SE_c_89_n N_10_c_398_n 4.38905e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_96 N_SE_c_89_n N_10_c_399_n 3.0053e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_97 N_SE_c_89_n N_10_c_400_n 7.16568e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_98 N_SE_c_89_n N_11_c_453_n 0.00113636f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_99 N_SE_c_89_n N_11_c_454_n 2.78297e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_100 N_SE_c_89_n N_11_c_455_n 5.99401e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_101 N_SE_c_89_n N_11_c_456_n 4.8504e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_102 N_SE_c_89_n N_11_c_457_n 4.65038e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_103 N_SE_c_89_n N_12_c_515_n 5.48108e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_104 N_SE_c_89_n N_12_c_516_n 0.00109158f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_105 N_SE_c_89_n N_12_c_517_n 5.50727e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_106 N_SE_c_89_n N_12_c_518_n 9.11285e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_107 N_SE_c_89_n N_12_c_519_n 4.62125e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_108 N_SE_c_89_n N_12_c_520_n 5.48546e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_109 N_SE_M14_g N_13_M15_g 0.00268443f $X=1.215 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_110 N_SE_c_126_p N_13_c_553_n 0.00112344f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_111 N_SE_c_89_n N_13_c_554_n 2.30689e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_112 N_SE_c_89_n N_13_c_555_n 9.08574e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_113 N_SE_c_89_n N_13_c_556_n 0.00124317f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_114 N_SE_c_89_n N_13_c_547_n 4.54245e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_115 N_SE_c_89_n N_13_c_558_n 4.39544e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_116 N_SE_c_89_n N_13_c_559_n 5.37888e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_117 N_SE_c_93_p N_13_c_560_n 3.26078e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_118 N_SE_c_89_n N_13_c_551_n 9.36021e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_119 N_SE_c_92_p N_13_c_562_n 9.36021e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_120 N_SE_c_136_p N_13_c_562_n 0.00114818f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_121 N_SE_c_137_p N_13_c_564_n 0.00409247f $X=1.215 $Y=0.113 $X2=0 $Y2=0
cc_122 N_SE_c_138_p N_14_c_618_n 2.31793e-19 $X=0.261 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_123 N_SE_M2_g N_14_c_619_n 3.83731e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_124 N_SE_c_140_p N_14_c_619_n 6.51345e-19 $X=0.258 $Y=0.135 $X2=0 $Y2=0
cc_125 VSS N_SE_c_86_n 2.40719e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.135
cc_126 VSS N_SE_c_88_n 5.30841e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.135
cc_127 VSS N_SE_c_105_p 9.86432e-19 $X=0.225 $Y=0.081 $X2=0.081 $Y2=0.135
cc_128 VSS N_SE_c_96_p 0.00129447f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_129 VSS N_SE_c_88_n 7.061e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_130 VSS N_SE_c_105_p 7.68051e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_131 VSS N_SE_c_86_n 8.44602e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.19
cc_132 VSS N_SE_c_88_n 5.36527e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.19
cc_133 VSS N_SE_c_89_n 0.00141783f $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.144
cc_134 VSS N_SE_c_89_n 2.35788e-19 $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.162
cc_135 VSS N_SE_c_88_n 6.93145e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.1785
cc_136 VSS N_SE_c_89_n 9.13621e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_137 VSS N_SE_c_89_n 4.6862e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_138 VSS N_SE_c_89_n 5.41611e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_139 VSS N_SE_c_89_n 8.51044e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_140 VSS N_SE_c_156_p 0.00129447f $X=0.279 $Y=0.135 $X2=0 $Y2=0
cc_141 VSS N_SE_c_88_n 3.48715e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_142 VSS N_SE_c_109_p 9.77595e-19 $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_143 VSS N_SE_c_89_n 2.40178e-19 $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.135
cc_144 VSS N_SE_c_89_n 6.42719e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_145 VSS N_SE_c_89_n 0.00110738f $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.162
cc_146 N_SE_c_94_p N_QN_c_667_n 3.2291e-19 $X=1.215 $Y=0.09 $X2=0.081 $Y2=0.19
cc_147 N_SE_c_93_p N_QN_c_668_n 8.07872e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_148 N_SE_c_89_n N_20_c_684_n 4.98441e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_149 N_6_M3_g N_D_M4_g 0.00304756f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_150 N_6_c_169_n N_D_c_237_n 9.71463e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_151 N_6_c_165_n D 3.33994e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_152 N_6_c_167_n D 0.00195518f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_153 N_6_c_179_n D 9.77589e-19 $X=0.351 $Y=0.126 $X2=0 $Y2=0
cc_154 N_6_M3_g N_SI_M5_g 2.48122e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_155 N_6_c_165_n SI 3.40688e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_156 N_6_c_187_p N_9_c_283_n 3.37164e-19 $X=0.936 $Y=0.081 $X2=0.891 $Y2=0.135
cc_157 N_6_c_165_n N_9_c_275_n 0.0011956f $X=0.9 $Y=0.081 $X2=0.817 $Y2=0.153
cc_158 N_6_c_165_n N_10_c_401_n 5.04077e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_159 N_6_c_165_n N_10_c_402_n 2.53924e-19 $X=0.9 $Y=0.081 $X2=0.056 $Y2=0.054
cc_160 N_6_c_165_n N_10_c_399_n 9.03945e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_161 N_6_c_165_n N_10_c_404_n 5.75824e-19 $X=0.9 $Y=0.081 $X2=0.018 $Y2=0.1125
cc_162 N_6_c_165_n N_10_c_405_n 7.91051e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_163 N_6_c_165_n N_11_c_454_n 4.20387e-19 $X=0.9 $Y=0.081 $X2=0.018 $Y2=0.081
cc_164 N_6_c_165_n N_11_c_459_n 4.92006e-19 $X=0.9 $Y=0.081 $X2=0.054 $Y2=0.036
cc_165 N_6_c_165_n N_11_c_460_n 7.19039e-19 $X=0.9 $Y=0.081 $X2=0.054 $Y2=0.036
cc_166 N_6_c_170_n N_12_c_521_n 0.00124414f $X=1.19 $Y=0.0405 $X2=0.621
+ $Y2=0.135
cc_167 N_6_c_172_n N_12_c_521_n 2.40393e-19 $X=1.161 $Y=0.081 $X2=0.621
+ $Y2=0.135
cc_168 N_6_c_199_p N_12_c_523_n 5.25714e-19 $X=1.19 $Y=0.2295 $X2=0.891
+ $Y2=0.0405
cc_169 N_6_c_172_n N_12_c_515_n 9.95523e-19 $X=1.161 $Y=0.081 $X2=0.891
+ $Y2=0.135
cc_170 N_6_c_170_n N_12_c_516_n 3.43147e-19 $X=1.19 $Y=0.0405 $X2=0.071
+ $Y2=0.054
cc_171 N_6_c_175_n N_12_c_516_n 0.00251979f $X=1.161 $Y=0.049 $X2=0.071
+ $Y2=0.054
cc_172 N_6_c_203_p N_12_c_527_n 0.00251979f $X=1.17 $Y=0.234 $X2=0.018 $Y2=0.045
cc_173 N_6_c_172_n N_12_c_520_n 0.0012739f $X=1.161 $Y=0.081 $X2=0.018 $Y2=0.144
cc_174 N_6_c_205_p N_12_c_520_n 0.00251979f $X=1.161 $Y=0.2125 $X2=0.018
+ $Y2=0.144
cc_175 N_6_c_206_p N_12_c_530_n 0.00251979f $X=1.161 $Y=0.225 $X2=0.018
+ $Y2=0.081
cc_176 N_6_c_187_p N_13_c_556_n 6.23859e-19 $X=0.936 $Y=0.081 $X2=0 $Y2=0
cc_177 N_6_c_172_n N_13_c_559_n 3.66836e-19 $X=1.161 $Y=0.081 $X2=0.018
+ $Y2=0.1125
cc_178 N_6_c_172_n N_13_c_567_n 5.24665e-19 $X=1.161 $Y=0.081 $X2=0.018
+ $Y2=0.162
cc_179 N_6_c_187_p N_13_c_568_n 3.12147e-19 $X=0.936 $Y=0.081 $X2=0.621
+ $Y2=0.135
cc_180 N_6_c_170_n N_13_c_551_n 2.50315e-19 $X=1.19 $Y=0.0405 $X2=0.621
+ $Y2=0.153
cc_181 N_6_c_212_p N_13_c_551_n 3.14624e-19 $X=1.179 $Y=0.234 $X2=0.621
+ $Y2=0.153
cc_182 N_6_c_172_n N_13_c_551_n 0.00815696f $X=1.161 $Y=0.081 $X2=0.621
+ $Y2=0.153
cc_183 N_6_c_175_n N_13_c_551_n 0.00110082f $X=1.161 $Y=0.049 $X2=0.621
+ $Y2=0.153
cc_184 N_6_c_199_p N_13_c_562_n 2.19627e-19 $X=1.19 $Y=0.2295 $X2=0.621
+ $Y2=0.153
cc_185 N_6_c_216_p N_13_c_562_n 3.14624e-19 $X=1.188 $Y=0.234 $X2=0.621
+ $Y2=0.153
cc_186 N_6_M3_g N_14_c_621_n 2.37298e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_187 VSS N_6_c_165_n 3.90811e-19 $X=0.9 $Y=0.081 $X2=0.621 $Y2=0.135
cc_188 VSS N_6_c_178_n 7.35661e-19 $X=0.351 $Y=0.099 $X2=0.621 $Y2=0.135
cc_189 VSS N_6_c_220_p 6.42252e-19 $X=0.351 $Y=0.081 $X2=0.621 $Y2=0.2295
cc_190 VSS N_6_c_220_p 0.00369658f $X=0.351 $Y=0.081 $X2=0.891 $Y2=0.135
cc_191 N_6_M3_g N_16_c_646_n 2.50526e-19 $X=0.351 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_192 N_6_c_167_n N_16_c_646_n 0.00110314f $X=0.351 $Y=0.135 $X2=0.891
+ $Y2=0.135
cc_193 VSS N_6_c_178_n 2.30452e-19 $X=0.351 $Y=0.099 $X2=0.135 $Y2=0.135
cc_194 VSS N_6_c_165_n 7.92007e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_195 VSS N_6_c_220_p 8.14481e-19 $X=0.351 $Y=0.081 $X2=0.891 $Y2=0.0405
cc_196 VSS N_6_c_165_n 2.67459e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_197 VSS N_6_c_165_n 3.16736e-19 $X=0.9 $Y=0.081 $X2=0.891 $Y2=0.135
cc_198 VSS N_6_c_165_n 2.43408e-19 $X=0.9 $Y=0.081 $X2=0.891 $Y2=0.135
cc_199 VSS N_6_c_165_n 5.19239e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_200 N_6_c_216_p N_QN_c_669_n 2.64332e-19 $X=1.188 $Y=0.234 $X2=0.071
+ $Y2=0.216
cc_201 N_6_c_187_p N_20_c_684_n 5.02041e-19 $X=0.936 $Y=0.081 $X2=0.621
+ $Y2=0.0675
cc_202 VSS N_6_c_220_p 2.73492e-19 $X=0.351 $Y=0.081 $X2=0.135 $Y2=0.054
cc_203 N_D_M4_g N_SI_M5_g 0.00348334f $X=0.405 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_204 D SI 7.00288e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_205 N_D_c_237_n N_SI_c_257_n 0.00109838f $X=0.405 $Y=0.135 $X2=0.621
+ $Y2=0.2295
cc_206 N_D_M4_g N_14_c_621_n 2.37298e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_207 VSS N_D_M4_g 3.08888e-19 $X=0.405 $Y=0.0675 $X2=0.891 $Y2=0.2295
cc_208 VSS D 5.77345e-19 $X=0.405 $Y=0.134 $X2=0.891 $Y2=0.2295
cc_209 N_D_M4_g N_16_c_648_n 2.43567e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_210 D N_16_c_648_n 0.00108212f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_211 D N_16_c_650_n 3.4434e-19 $X=0.405 $Y=0.134 $X2=0.071 $Y2=0.054
cc_212 VSS D 8.86227e-19 $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.135
cc_213 VSS D 0.00161923f $X=0.405 $Y=0.134 $X2=0.891 $Y2=0.0405
cc_214 N_SI_M5_g N_9_c_279_n 2.94371e-19 $X=0.459 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_215 N_SI_c_257_n N_9_c_279_n 5.18435e-19 $X=0.475 $Y=0.135 $X2=0.135
+ $Y2=0.054
cc_216 SI N_9_c_290_n 0.00114959f $X=0.473 $Y=0.135 $X2=0 $Y2=0
cc_217 SI N_9_c_315_n 0.00114959f $X=0.473 $Y=0.135 $X2=0.054 $Y2=0.234
cc_218 SI N_9_c_296_n 0.00239259f $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.153
cc_219 SI N_9_c_275_n 0.00167124f $X=0.473 $Y=0.135 $X2=0.817 $Y2=0.153
cc_220 SI N_14_c_617_n 0.00560919f $X=0.473 $Y=0.135 $X2=0.621 $Y2=0.2295
cc_221 SI N_14_c_624_n 0.00167456f $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.135
cc_222 N_SI_M5_g N_14_c_625_n 2.70361e-19 $X=0.459 $Y=0.0675 $X2=0.071 $Y2=0.054
cc_223 SI N_16_c_651_n 6.69571e-19 $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.0405
cc_224 VSS N_SI_M5_g 3.10987e-19 $X=0.459 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_225 VSS N_SI_c_257_n 2.08525e-19 $X=0.475 $Y=0.135 $X2=0.891 $Y2=0.135
cc_226 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.135
cc_227 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.2295
cc_228 VSS SI 0.00110314f $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.2295
cc_229 N_9_M7_g N_10_M8_g 0.00341068f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_230 N_9_M10_g N_10_M8_g 2.13359e-19 $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_231 N_9_c_283_n N_10_M8_g 0.00205997f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_232 N_9_c_299_n N_10_M8_g 3.19768e-19 $X=0.729 $Y=0.18 $X2=0.081 $Y2=0.054
cc_233 N_9_c_283_n N_10_c_398_n 5.49754e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_234 N_9_c_283_n N_10_c_411_n 2.12581e-19 $X=0.945 $Y=0.178 $X2=0.081
+ $Y2=0.144
cc_235 N_9_c_283_n N_10_M26_s 2.50995e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.167
cc_236 N_9_M10_g N_10_c_413_n 0.00200065f $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_237 N_9_c_283_n N_10_c_413_n 0.00303373f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_238 N_9_M10_g N_10_c_396_n 2.74825e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_239 N_9_M10_g N_10_c_397_n 2.10136e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_240 N_9_c_299_n N_10_c_417_n 6.73839e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_241 N_9_c_330_p N_10_c_418_n 0.00195059f $X=0.837 $Y=0.178 $X2=0 $Y2=0
cc_242 N_9_c_283_n N_10_c_418_n 0.00191847f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_243 N_9_M10_g N_10_c_405_n 3.61755e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_244 N_9_M7_g N_11_M9_g 2.13359e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_245 N_9_M10_g N_11_M9_g 0.00341068f $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_246 N_9_c_283_n N_11_M9_g 0.00302156f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_247 N_9_c_290_n N_11_c_444_n 7.70794e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_248 N_9_c_296_n N_11_c_444_n 0.001307f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_249 N_9_c_296_n N_11_c_466_n 0.00138499f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_250 N_9_c_275_n N_11_c_467_n 0.00160025f $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_251 N_9_M7_g N_11_c_453_n 4.38308e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_252 N_9_M7_g N_11_c_459_n 2.0845e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_253 N_9_M7_g N_11_c_460_n 2.27141e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_254 N_9_c_283_n N_11_c_449_n 0.0361494f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_255 N_9_c_283_n N_11_c_472_n 2.38252e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_256 N_9_c_299_n N_11_c_472_n 0.00386452f $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_257 N_9_c_346_p N_11_c_474_n 7.00743e-19 $X=0.675 $Y=0.178 $X2=0 $Y2=0
cc_258 N_9_c_283_n N_11_c_474_n 7.89771e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_259 N_9_c_275_n N_11_c_474_n 4.88732e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_260 N_9_M7_g N_11_c_477_n 2.5554e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_261 N_9_c_283_n N_11_c_477_n 3.47488e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_262 N_9_c_296_n N_11_c_477_n 2.13133e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_263 N_9_c_275_n N_11_c_477_n 4.32971e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_264 N_9_c_299_n N_11_c_477_n 2.60223e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_265 N_9_c_283_n N_11_c_451_n 4.76652e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_266 N_9_c_283_n N_11_c_452_n 4.41163e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_267 N_9_c_283_n N_11_c_484_n 3.33141e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_268 N_9_c_299_n N_11_c_484_n 9.1388e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_269 N_9_M7_g N_11_c_486_n 2.12062e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_270 N_9_c_283_n N_12_M12_g 0.00341068f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_271 N_9_c_283_n N_13_M13_g 2.13359e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_272 N_9_c_283_n N_13_c_554_n 8.27183e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_273 N_9_c_283_n N_13_M27_s 3.37661e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_274 N_9_c_283_n N_13_c_578_n 0.00145657f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_275 N_9_c_283_n N_13_c_567_n 3.13444e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_276 N_9_c_283_n N_13_c_580_n 2.6418e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_277 N_9_c_283_n N_13_c_581_n 0.00294656f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_278 N_9_c_283_n N_13_c_568_n 3.75802e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_279 N_9_c_283_n N_13_c_550_n 5.46321e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_280 N_9_c_289_n N_14_c_618_n 9.65806e-19 $X=0.16 $Y=0.216 $X2=0.081 $Y2=0.135
cc_281 N_9_c_275_n N_14_c_618_n 4.65646e-19 $X=0.729 $Y=0.189 $X2=0.081
+ $Y2=0.135
cc_282 N_9_c_301_n N_14_c_618_n 0.00109797f $X=0.189 $Y=0.164 $X2=0.081
+ $Y2=0.135
cc_283 N_9_c_290_n N_14_c_617_n 9.68946e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_284 N_9_c_275_n N_14_c_617_n 6.49405e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_285 N_9_c_374_p N_14_c_619_n 7.61293e-19 $X=0.189 $Y=0.234 $X2=0 $Y2=0
cc_286 N_9_c_275_n N_14_c_619_n 7.84624e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_287 N_9_c_275_n N_14_c_625_n 6.22262e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_288 VSS N_9_c_288_n 9.30745e-19 $X=0.16 $Y=0.054 $X2=0.081 $Y2=0.135
cc_289 N_9_c_275_n N_16_c_652_n 2.13751e-19 $X=0.729 $Y=0.189 $X2=0.081
+ $Y2=0.135
cc_290 N_9_c_275_n N_16_c_651_n 7.1298e-19 $X=0.729 $Y=0.189 $X2=0.081 $Y2=0.162
cc_291 N_9_c_275_n N_16_c_654_n 6.46208e-19 $X=0.729 $Y=0.189 $X2=0.081
+ $Y2=0.1785
cc_292 N_9_c_275_n N_16_c_646_n 4.50553e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_293 N_9_c_275_n N_16_c_656_n 4.86474e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_294 N_9_c_275_n N_16_c_657_n 4.60071e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_295 N_9_c_275_n N_16_c_648_n 4.38038e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_296 N_9_c_275_n N_16_c_650_n 2.31538e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_297 VSS N_9_c_279_n 3.33061e-19 $X=0.567 $Y=0.1355 $X2=0 $Y2=0
cc_298 VSS N_9_c_290_n 0.00110314f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_299 N_9_c_283_n N_19_M24_s 2.33161e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.216
cc_300 N_9_M7_g N_19_c_675_n 0.00248549f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_301 N_9_c_283_n N_19_c_675_n 0.00208457f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_302 N_9_c_275_n N_19_c_675_n 7.88525e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_303 N_9_c_283_n N_20_c_684_n 0.00250239f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_304 N_10_M8_g N_11_M9_g 0.00268443f $X=0.729 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_305 N_10_c_399_n N_11_M9_g 3.80603e-19 $X=0.797 $Y=0.09 $X2=0.135 $Y2=0.054
cc_306 N_10_c_400_n N_11_c_457_n 2.46574e-19 $X=0.81 $Y=0.054 $X2=0.027
+ $Y2=0.036
cc_307 N_10_c_401_n N_11_c_490_n 0.00360624f $X=0.747 $Y=0.09 $X2=0.054
+ $Y2=0.036
cc_308 N_10_c_402_n N_11_c_459_n 3.99428e-19 $X=0.747 $Y=0.09 $X2=0.054
+ $Y2=0.036
cc_309 N_10_c_397_n N_11_c_448_n 2.22221e-19 $X=0.837 $Y=0.165 $X2=0.054
+ $Y2=0.234
cc_310 N_10_c_427_p N_11_c_477_n 2.22221e-19 $X=0.837 $Y=0.225 $X2=0.0505
+ $Y2=0.234
cc_311 N_10_c_399_n N_11_c_451_n 0.00219679f $X=0.797 $Y=0.09 $X2=0.621
+ $Y2=0.135
cc_312 N_10_c_429_p N_11_c_451_n 9.66928e-19 $X=0.837 $Y=0.14 $X2=0.621
+ $Y2=0.135
cc_313 N_10_M8_g N_11_c_484_n 3.21351e-19 $X=0.729 $Y=0.0405 $X2=0.033 $Y2=0.153
cc_314 N_10_c_401_n N_11_c_484_n 0.00219679f $X=0.747 $Y=0.09 $X2=0.033
+ $Y2=0.153
cc_315 N_10_c_398_n N_13_c_554_n 0.00379158f $X=0.81 $Y=0.0405 $X2=0.891
+ $Y2=0.135
cc_316 N_10_c_400_n N_13_c_554_n 2.84891e-19 $X=0.81 $Y=0.054 $X2=0.891
+ $Y2=0.135
cc_317 N_10_c_405_n N_13_c_554_n 2.08929e-19 $X=0.837 $Y=0.09 $X2=0.891
+ $Y2=0.135
cc_318 N_10_c_413_n N_13_c_578_n 0.00222825f $X=0.866 $Y=0.2295 $X2=0.056
+ $Y2=0.054
cc_319 N_10_c_398_n N_13_c_556_n 3.41768e-19 $X=0.81 $Y=0.0405 $X2=0 $Y2=0
cc_320 N_10_c_405_n N_13_c_567_n 4.2911e-19 $X=0.837 $Y=0.09 $X2=0.018 $Y2=0.162
cc_321 N_10_c_418_n N_13_c_581_n 4.2911e-19 $X=0.837 $Y=0.207 $X2=0.027
+ $Y2=0.036
cc_322 N_10_c_413_n N_13_c_568_n 3.64454e-19 $X=0.866 $Y=0.2295 $X2=0.621
+ $Y2=0.135
cc_323 N_10_c_440_p N_13_c_568_n 4.86017e-19 $X=0.828 $Y=0.234 $X2=0.621
+ $Y2=0.135
cc_324 N_10_c_441_p N_13_c_550_n 4.2911e-19 $X=0.837 $Y=0.101 $X2=0 $Y2=0
cc_325 N_11_c_444_n N_14_c_617_n 0.00424458f $X=0.594 $Y=0.2025 $X2=0.621
+ $Y2=0.2295
cc_326 N_11_c_466_n N_14_c_617_n 4.3429e-19 $X=0.595 $Y=0.234 $X2=0.621
+ $Y2=0.2295
cc_327 N_11_c_466_n N_14_c_624_n 2.8677e-19 $X=0.595 $Y=0.234 $X2=0.891
+ $Y2=0.135
cc_328 VSS N_11_c_444_n 0.0016174f $X=0.594 $Y=0.2025 $X2=0.621 $Y2=0.0675
cc_329 VSS N_11_c_454_n 0.00414127f $X=0.648 $Y=0.036 $X2=0.621 $Y2=0.0675
cc_330 VSS N_11_c_455_n 3.30384e-19 $X=0.649 $Y=0.036 $X2=0.621 $Y2=0.0675
cc_331 VSS N_11_c_454_n 2.79363e-19 $X=0.648 $Y=0.036 $X2=0 $Y2=0
cc_332 VSS N_11_c_459_n 2.70508e-19 $X=0.693 $Y=0.081 $X2=0 $Y2=0
cc_333 N_11_c_444_n N_19_c_675_n 0.00167238f $X=0.594 $Y=0.2025 $X2=0.621
+ $Y2=0.0675
cc_334 N_11_c_507_p N_19_c_675_n 0.00315491f $X=0.684 $Y=0.234 $X2=0.621
+ $Y2=0.0675
cc_335 N_11_c_445_n N_19_c_675_n 0.00111131f $X=0.649 $Y=0.234 $X2=0.621
+ $Y2=0.0675
cc_336 N_11_c_454_n N_19_c_675_n 5.67227e-19 $X=0.648 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_337 N_11_c_510_p N_19_c_675_n 4.0515e-19 $X=0.693 $Y=0.225 $X2=0.621
+ $Y2=0.0675
cc_338 N_11_c_511_p N_19_c_675_n 0.0409693f $X=0.693 $Y=0.216 $X2=0.621
+ $Y2=0.0675
cc_339 N_11_c_453_n N_22_M8_s 2.44135e-19 $X=0.684 $Y=0.036 $X2=0.135 $Y2=0.054
cc_340 N_11_c_457_n N_22_M8_s 3.62465e-19 $X=0.693 $Y=0.062 $X2=0.135 $Y2=0.054
cc_341 N_12_M12_g N_13_M13_g 0.00268443f $X=0.999 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_342 N_12_c_519_n N_13_M13_g 3.55314e-19 $X=1.062 $Y=0.036 $X2=0.135 $Y2=0.054
cc_343 N_12_c_517_n N_13_c_555_n 0.00136796f $X=1.008 $Y=0.036 $X2=0 $Y2=0
cc_344 N_12_c_515_n N_13_c_559_n 0.00136796f $X=0.999 $Y=0.105 $X2=0.018
+ $Y2=0.1125
cc_345 N_12_c_536_p N_13_c_567_n 3.34766e-19 $X=0.999 $Y=0.1055 $X2=0.018
+ $Y2=0.162
cc_346 N_12_c_515_n N_13_c_567_n 0.00136796f $X=0.999 $Y=0.105 $X2=0.018
+ $Y2=0.162
cc_347 N_12_c_527_n N_13_c_581_n 5.28703e-19 $X=1.107 $Y=0.225 $X2=0.027
+ $Y2=0.036
cc_348 N_12_M12_g N_13_c_601_n 6.35734e-19 $X=0.999 $Y=0.0405 $X2=0.047
+ $Y2=0.036
cc_349 N_12_c_515_n N_13_c_601_n 7.99759e-19 $X=0.999 $Y=0.105 $X2=0.047
+ $Y2=0.036
cc_350 N_12_c_519_n N_13_c_603_n 2.75024e-19 $X=1.062 $Y=0.036 $X2=0.027
+ $Y2=0.234
cc_351 N_12_c_530_n N_13_c_603_n 0.00266666f $X=1.107 $Y=0.171 $X2=0.027
+ $Y2=0.234
cc_352 N_12_c_523_n N_13_c_551_n 2.19627e-19 $X=1.078 $Y=0.2295 $X2=0.621
+ $Y2=0.153
cc_353 N_12_c_530_n N_13_c_551_n 0.00106087f $X=1.107 $Y=0.171 $X2=0.621
+ $Y2=0.153
cc_354 N_12_c_545_p N_13_c_551_n 5.80975e-19 $X=1.098 $Y=0.234 $X2=0.621
+ $Y2=0.153
cc_355 N_12_c_517_n N_20_c_684_n 5.06067e-19 $X=1.008 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_356 N_13_c_564_n N_QN_c_670_n 0.00114532f $X=1.269 $Y=0.136 $X2=0.621
+ $Y2=0.0675
cc_357 N_13_c_560_n N_QN_c_671_n 2.31819e-19 $X=1.269 $Y=0.153 $X2=0 $Y2=0
cc_358 N_13_c_564_n N_QN_c_671_n 0.00431194f $X=1.269 $Y=0.136 $X2=0 $Y2=0
cc_359 N_13_c_564_n N_QN_c_673_n 5.42522e-19 $X=1.269 $Y=0.136 $X2=0 $Y2=0
cc_360 N_13_c_554_n N_20_c_684_n 0.00210698f $X=0.864 $Y=0.0405 $X2=0.621
+ $Y2=0.0675
cc_361 N_13_c_555_n N_20_c_684_n 0.00203632f $X=0.936 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_362 N_13_c_558_n N_20_c_684_n 0.00129774f $X=0.92 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_363 N_13_c_559_n N_20_c_684_n 0.00104094f $X=0.945 $Y=0.081 $X2=0.621
+ $Y2=0.0675
cc_364 N_13_c_616_p N_20_c_684_n 2.5109e-19 $X=0.99 $Y=0.162 $X2=0.621
+ $Y2=0.0675
cc_365 VSS N_14_c_618_n 0.00156967f $X=0.272 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_366 VSS N_14_c_617_n 0.00145555f $X=0.542 $Y=0.2025 $X2=0.891 $Y2=0.0405
cc_367 N_14_c_618_n N_16_c_660_n 0.003872f $X=0.272 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_368 N_14_c_621_n N_16_c_660_n 0.00248801f $X=0.447 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_369 N_14_c_617_n N_16_c_662_n 0.00434154f $X=0.542 $Y=0.2025 $X2=0.621
+ $Y2=0.0675
cc_370 N_14_c_621_n N_16_c_662_n 0.0025506f $X=0.447 $Y=0.234 $X2=0.621
+ $Y2=0.0675
cc_371 N_14_c_618_n N_16_c_652_n 3.19827e-19 $X=0.272 $Y=0.2025 $X2=0.621
+ $Y2=0.135
cc_372 N_14_c_621_n N_16_c_652_n 0.0113176f $X=0.447 $Y=0.234 $X2=0.621
+ $Y2=0.135
cc_373 VSS N_14_c_617_n 4.53012e-19 $X=0.542 $Y=0.2025 $X2=0 $Y2=0
cc_374 VSS N_16_c_662_n 0.00141703f $X=0.432 $Y=0.2025 $X2=0.135 $Y2=0.135

* END of "./SDFHx1_ASAP7_75t_SRAM.pex.sp.SDFHX1_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: SDFHx2_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 13:03:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "SDFHx2_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./SDFHx2_ASAP7_75t_SRAM.pex.sp.pex"
* File: SDFHx2_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 13:03:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_SDFHX2_ASAP7_75T_SRAM%CLK 2 5 7 11 16 18 19 20 VSS
c19 20 VSS 1.17072e-19 $X=0.081 $Y=0.1785
c20 19 VSS 3.55344e-20 $X=0.081 $Y=0.167
c21 18 VSS 9.34089e-20 $X=0.081 $Y=0.162
c22 16 VSS 0.00100628f $X=0.078 $Y=0.19
c23 11 VSS 0.00681069f $X=0.081 $Y=0.135
c24 5 VSS 0.00208806f $X=0.081 $Y=0.135
c25 2 VSS 0.0627545f $X=0.081 $Y=0.054
r26 19 20 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.167 $X2=0.081 $Y2=0.1785
r27 18 19 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.162 $X2=0.081 $Y2=0.167
r28 17 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.144 $X2=0.081 $Y2=0.162
r29 16 20 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.19 $X2=0.081 $Y2=0.1785
r30 11 17 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.144
r31 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r32 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r33 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%4 2 5 7 10 13 15 18 21 23 25 28 30 36 37 38 41 45
+ 52 59 64 71 72 73 74 75 77 79 80 84 92 VSS
c65 111 VSS 1.06551e-19 $X=0.03 $Y=0.153
c66 110 VSS 6.89947e-19 $X=0.027 $Y=0.153
c67 92 VSS 0.001222f $X=0.891 $Y=0.135
c68 84 VSS 0.00111816f $X=0.135 $Y=0.135
c69 80 VSS 0.00209834f $X=0.817 $Y=0.153
c70 79 VSS 0.00159119f $X=0.743 $Y=0.153
c71 77 VSS 0.00277988f $X=0.891 $Y=0.153
c72 75 VSS 0.0014306f $X=0.479 $Y=0.153
c73 74 VSS 0.00120845f $X=0.337 $Y=0.153
c74 73 VSS 9.39788e-19 $X=0.211 $Y=0.153
c75 72 VSS 0.00665478f $X=0.175 $Y=0.153
c76 71 VSS 9.40943e-19 $X=0.621 $Y=0.153
c77 64 VSS 6.72589e-19 $X=0.033 $Y=0.153
c78 59 VSS 5.26559e-19 $X=0.621 $Y=0.135
c79 55 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c80 54 VSS 0.00180216f $X=0.047 $Y=0.234
c81 52 VSS 0.00253483f $X=0.054 $Y=0.234
c82 50 VSS 0.00305101f $X=0.027 $Y=0.234
c83 48 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c84 47 VSS 0.00199699f $X=0.047 $Y=0.036
c85 45 VSS 0.00239525f $X=0.054 $Y=0.036
c86 43 VSS 0.00305101f $X=0.027 $Y=0.036
c87 42 VSS 5.16336e-19 $X=0.018 $Y=0.2125
c88 41 VSS 0.00180713f $X=0.018 $Y=0.2
c89 40 VSS 4.96914e-19 $X=0.018 $Y=0.225
c90 38 VSS 0.00159315f $X=0.018 $Y=0.1125
c91 37 VSS 0.00142827f $X=0.018 $Y=0.081
c92 36 VSS 0.00143809f $X=0.018 $Y=0.144
c93 33 VSS 0.0049466f $X=0.056 $Y=0.216
c94 30 VSS 2.98509e-19 $X=0.071 $Y=0.216
c95 28 VSS 0.00460164f $X=0.056 $Y=0.054
c96 25 VSS 2.98509e-19 $X=0.071 $Y=0.054
c97 21 VSS 0.00216055f $X=0.891 $Y=0.135
c98 18 VSS 0.0585656f $X=0.891 $Y=0.0405
c99 13 VSS 0.00201785f $X=0.621 $Y=0.135
c100 10 VSS 0.0601628f $X=0.621 $Y=0.0675
c101 5 VSS 0.00199564f $X=0.135 $Y=0.135
c102 2 VSS 0.0630095f $X=0.135 $Y=0.054
r103 110 111 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r104 107 110 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r105 79 80 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.743
+ $Y=0.153 $X2=0.817 $Y2=0.153
r106 77 80 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.817 $Y2=0.153
r107 77 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r108 74 75 9.64198 $w=1.8e-08 $l=1.42e-07 $layer=M2 $thickness=3.6e-08 $X=0.337
+ $Y=0.153 $X2=0.479 $Y2=0.153
r109 73 74 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.211
+ $Y=0.153 $X2=0.337 $Y2=0.153
r110 72 73 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.175
+ $Y=0.153 $X2=0.211 $Y2=0.153
r111 70 79 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.743 $Y2=0.153
r112 70 75 9.64198 $w=1.8e-08 $l=1.42e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.479 $Y2=0.153
r113 70 71 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.621 $Y=0.153 $X2=0.621
+ $Y2=0.153
r114 67 72 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.153 $X2=0.175 $Y2=0.153
r115 67 84 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.135 $Y=0.153 $X2=0.135
+ $Y2=0.153
r116 64 111 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r117 63 67 6.92593 $w=1.8e-08 $l=1.02e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.135 $Y2=0.153
r118 63 64 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r119 59 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.153
r120 54 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r121 52 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r122 50 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r123 47 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r124 45 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r125 43 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r126 41 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r127 40 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r128 40 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r129 39 107 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r130 39 41 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.2
r131 37 38 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.1125
r132 36 107 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r133 36 38 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1125
r134 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r135 35 37 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r136 33 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r137 30 33 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r138 28 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r139 25 28 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r140 21 92 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.135 $X2=0.891
+ $Y2=0.135
r141 21 23 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.135 $X2=0.891 $Y2=0.2295
r142 18 21 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.0405 $X2=0.891 $Y2=0.135
r143 13 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r144 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2295
r145 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r146 5 84 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r147 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r148 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%SE 2 5 7 10 13 15 19 22 23 24 31 33 41 44 45 46 47
+ 54 58 59 62 63 VSS
c79 63 VSS 2.09605e-19 $X=1.215 $Y=0.113
c80 62 VSS 0.00191998f $X=1.215 $Y=0.09
c81 59 VSS 2.63823e-19 $X=0.225 $Y=0.099
c82 58 VSS 5.90201e-19 $X=0.225 $Y=0.081
c83 54 VSS 0.00128636f $X=1.215 $Y=0.136
c84 47 VSS 0.0383019f $X=1.175 $Y=0.045
c85 46 VSS 0.00642311f $X=0.337 $Y=0.045
c86 45 VSS 0.00700571f $X=1.215 $Y=0.045
c87 44 VSS 0.00307515f $X=1.215 $Y=0.045
c88 41 VSS 0.00531f $X=0.225 $Y=0.045
c89 31 VSS 0.00110873f $X=0.225 $Y=0.126
c90 24 VSS 2.51525e-19 $X=0.279 $Y=0.135
c91 23 VSS 1.48251e-19 $X=0.261 $Y=0.135
c92 22 VSS 6.38823e-20 $X=0.258 $Y=0.135
c93 21 VSS 0.00134071f $X=0.255 $Y=0.135
c94 19 VSS 6.89032e-19 $X=0.297 $Y=0.135
c95 13 VSS 0.00244398f $X=1.215 $Y=0.136
c96 10 VSS 0.0611074f $X=1.215 $Y=0.0405
c97 5 VSS 0.00319967f $X=0.297 $Y=0.135
c98 2 VSS 0.063344f $X=0.297 $Y=0.0675
r99 62 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.09 $X2=1.215 $Y2=0.113
r100 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.081 $X2=0.225 $Y2=0.099
r101 54 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.136 $X2=1.215 $Y2=0.113
r102 46 47 56.9012 $w=1.8e-08 $l=8.38e-07 $layer=M2 $thickness=3.6e-08 $X=0.337
+ $Y=0.045 $X2=1.175 $Y2=0.045
r103 45 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.215 $Y2=0.09
r104 44 47 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.175 $Y2=0.045
r105 44 45 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.215 $Y=0.045 $X2=1.215
+ $Y2=0.045
r106 41 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.081
r107 40 46 7.60494 $w=1.8e-08 $l=1.12e-07 $layer=M2 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.337 $Y2=0.045
r108 40 41 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.225 $Y=0.045 $X2=0.225
+ $Y2=0.045
r109 31 59 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.099
r110 31 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r111 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.135 $X2=0.279 $Y2=0.135
r112 22 23 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.258
+ $Y=0.135 $X2=0.261 $Y2=0.135
r113 21 22 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.255
+ $Y=0.135 $X2=0.258 $Y2=0.135
r114 19 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.279 $Y2=0.135
r115 17 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.225 $Y2=0.135
r116 17 21 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.255 $Y2=0.135
r117 13 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.215 $Y=0.136 $X2=1.215
+ $Y2=0.136
r118 13 15 350.298 $w=2e-08 $l=9.35e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.136 $X2=1.215 $Y2=0.2295
r119 10 13 357.791 $w=2e-08 $l=9.55e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.0405 $X2=1.215 $Y2=0.136
r120 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r121 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r122 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%6 2 5 7 9 12 14 17 23 26 28 29 33 36 38 39 43 51
+ 57 58 65 VSS
c69 65 VSS 3.21273e-19 $X=1.161 $Y=0.2125
c70 58 VSS 5.45782e-19 $X=0.351 $Y=0.126
c71 57 VSS 8.0335e-19 $X=0.351 $Y=0.099
c72 51 VSS 0.00324902f $X=1.161 $Y=0.049
c73 43 VSS 3.66031e-19 $X=0.351 $Y=0.135
c74 39 VSS 9.89222e-19 $X=0.936 $Y=0.081
c75 38 VSS 0.00685031f $X=0.9 $Y=0.081
c76 36 VSS 0.00169093f $X=1.161 $Y=0.081
c77 33 VSS 8.10983e-19 $X=0.351 $Y=0.081
c78 29 VSS 7.48824e-19 $X=1.179 $Y=0.234
c79 28 VSS 0.00240687f $X=1.17 $Y=0.234
c80 26 VSS 0.00328115f $X=1.188 $Y=0.234
c81 23 VSS 9.88154e-20 $X=1.161 $Y=0.225
c82 17 VSS 0.00404882f $X=1.19 $Y=0.2295
c83 14 VSS 2.95772e-19 $X=1.205 $Y=0.2295
c84 12 VSS 0.060801f $X=1.19 $Y=0.0405
c85 9 VSS 3.14771e-19 $X=1.205 $Y=0.0405
c86 5 VSS 0.00125227f $X=0.351 $Y=0.135
c87 2 VSS 0.0585837f $X=0.351 $Y=0.0675
r88 64 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.2 $X2=1.161 $Y2=0.2125
r89 57 58 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.099 $X2=0.351 $Y2=0.126
r90 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.161 $Y=0.049 $X2=1.161
+ $Y2=0.049
r91 43 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.126
r92 38 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.9
+ $Y=0.081 $X2=0.936 $Y2=0.081
r93 37 64 8.08025 $w=1.8e-08 $l=1.19e-07 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.2
r94 37 51 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.049
r95 36 39 15.2778 $w=1.8e-08 $l=2.25e-07 $layer=M2 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=0.936 $Y2=0.081
r96 36 37 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.161 $Y=0.081 $X2=1.161
+ $Y2=0.081
r97 33 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.099
r98 32 38 37.2778 $w=1.8e-08 $l=5.49e-07 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.9 $Y2=0.081
r99 32 33 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.081 $X2=0.351
+ $Y2=0.081
r100 28 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.17
+ $Y=0.234 $X2=1.179 $Y2=0.234
r101 26 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.188
+ $Y=0.234 $X2=1.179 $Y2=0.234
r102 23 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.225 $X2=1.161 $Y2=0.2125
r103 22 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.17 $Y2=0.234
r104 22 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.161 $Y2=0.225
r105 17 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.188 $Y=0.234
+ $X2=1.188 $Y2=0.234
r106 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.2295 $X2=1.19 $Y2=0.2295
r107 12 50 16.2355 $w=3.7e-08 $l=2.9e-08 $layer=LISD $thickness=2.8e-08 $X=1.19
+ $Y=0.0455 $X2=1.161 $Y2=0.0455
r108 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.0405 $X2=1.19 $Y2=0.0405
r109 5 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r110 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r111 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%D 2 5 7 11 VSS
c18 11 VSS 0.00145113f $X=0.405 $Y=0.134
c19 5 VSS 0.00106786f $X=0.405 $Y=0.135
c20 2 VSS 0.0589243f $X=0.405 $Y=0.0675
r21 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%SI 2 7 11 14 VSS
c21 14 VSS 0.0032805f $X=0.475 $Y=0.135
c22 11 VSS 0.0035781f $X=0.473 $Y=0.135
c23 2 VSS 0.0640988f $X=0.459 $Y=0.0675
r24 11 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.475 $Y=0.135 $X2=0.475
+ $Y2=0.135
r25 5 14 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.475 $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%9 2 5 8 11 14 17 20 23 37 40 42 45 49 53 58 60 67
+ 69 74 78 80 96 101 102 103 104 106 VSS
c121 108 VSS 7.92414e-20 $X=0.189 $Y=0.207
c122 106 VSS 2.53862e-19 $X=0.189 $Y=0.178
c123 105 VSS 3.91706e-20 $X=0.189 $Y=0.167
c124 104 VSS 6.6467e-19 $X=0.189 $Y=0.164
c125 103 VSS 3.3761e-19 $X=0.189 $Y=0.144
c126 102 VSS 4.92067e-19 $X=0.189 $Y=0.121
c127 101 VSS 8.32677e-19 $X=0.189 $Y=0.099
c128 96 VSS 6.49238e-19 $X=0.729 $Y=0.18
c129 80 VSS 0.0152374f $X=0.729 $Y=0.189
c130 78 VSS 0.0013748f $X=0.567 $Y=0.189
c131 74 VSS 6.28429e-19 $X=0.189 $Y=0.189
c132 69 VSS 0.00386366f $X=0.18 $Y=0.234
c133 68 VSS 4.87314e-19 $X=0.189 $Y=0.225
c134 67 VSS 0.00199636f $X=0.189 $Y=0.234
c135 60 VSS 0.00373046f $X=0.18 $Y=0.036
c136 58 VSS 0.00194932f $X=0.189 $Y=0.036
c137 53 VSS 9.61695e-20 $X=0.567 $Y=0.18
c138 49 VSS 5.76385e-19 $X=0.567 $Y=0.135
c139 45 VSS 0.00566559f $X=0.16 $Y=0.216
c140 40 VSS 0.0055918f $X=0.16 $Y=0.054
c141 20 VSS 0.108836f $X=0.945 $Y=0.178
c142 17 VSS 1.08457e-19 $X=0.837 $Y=0.178
c143 14 VSS 0.0600244f $X=0.837 $Y=0.0405
c144 11 VSS 2.24613e-19 $X=0.675 $Y=0.178
c145 8 VSS 0.0602569f $X=0.675 $Y=0.0405
c146 2 VSS 0.0660345f $X=0.567 $Y=0.1355
r147 107 108 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.2 $X2=0.189 $Y2=0.207
r148 105 106 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.167 $X2=0.189 $Y2=0.178
r149 104 105 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.167
r150 103 104 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.164
r151 102 103 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.121 $X2=0.189 $Y2=0.144
r152 101 102 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.099 $X2=0.189 $Y2=0.121
r153 95 96 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.729 $Y=0.18 $X2=0.729
+ $Y2=0.18
r154 80 96 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.729 $Y=0.189 $X2=0.729
+ $Y2=0.189
r155 77 80 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.729 $Y2=0.189
r156 77 78 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.567 $Y=0.189 $X2=0.567
+ $Y2=0.189
r157 74 107 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.2
r158 74 106 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.178
r159 73 77 25.6667 $w=1.8e-08 $l=3.78e-07 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.567 $Y2=0.189
r160 73 74 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.189 $X2=0.189
+ $Y2=0.189
r161 69 70 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r162 68 108 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.207
r163 67 70 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r164 67 68 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.189 $Y2=0.225
r165 64 69 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r166 60 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r167 59 101 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.099
r168 58 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r169 58 59 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r170 55 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r171 53 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.18 $X2=0.567 $Y2=0.189
r172 52 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.171 $X2=0.567 $Y2=0.18
r173 49 52 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.171
r174 45 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r175 42 45 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r176 40 55 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r177 37 40 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r178 20 23 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.178 $X2=0.945 $Y2=0.2295
r179 17 20 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08 $X=0.837
+ $Y=0.178 $X2=0.945 $Y2=0.178
r180 17 95 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08 $X=0.837
+ $Y=0.178 $X2=0.729 $Y2=0.178
r181 14 17 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0405 $X2=0.837 $Y2=0.178
r182 11 95 43.022 $w=2.6e-08 $l=5.4e-08 $layer=LISD $thickness=2.8e-08 $X=0.675
+ $Y=0.178 $X2=0.729 $Y2=0.178
r183 8 11 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.178
r184 2 49 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r185 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1355 $X2=0.567 $Y2=0.2025
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%10 2 7 9 10 13 14 17 19 22 27 28 29 31 36 38 44 45
+ 46 47 48 49 50 54 VSS
c49 56 VSS 5.19568e-19 $X=0.828 $Y=0.09
c50 55 VSS 4.09996e-19 $X=0.819 $Y=0.09
c51 54 VSS 4.29e-19 $X=0.837 $Y=0.09
c52 50 VSS 5.92866e-19 $X=0.837 $Y=0.207
c53 49 VSS 1.19762e-19 $X=0.837 $Y=0.167
c54 48 VSS 1.59501e-19 $X=0.837 $Y=0.165
c55 47 VSS 3.13056e-19 $X=0.837 $Y=0.14
c56 46 VSS 5.61414e-19 $X=0.837 $Y=0.122
c57 45 VSS 1.91116e-19 $X=0.837 $Y=0.101
c58 44 VSS 4.02479e-19 $X=0.837 $Y=0.225
c59 42 VSS 3.58124e-20 $X=0.81 $Y=0.0715
c60 38 VSS 0.00112276f $X=0.81 $Y=0.054
c61 31 VSS 0.00670205f $X=0.828 $Y=0.234
c62 30 VSS 4.74851e-19 $X=0.7965 $Y=0.09
c63 29 VSS 0.00125276f $X=0.792 $Y=0.09
c64 28 VSS 0.00410211f $X=0.747 $Y=0.09
c65 27 VSS 4.49532e-19 $X=0.747 $Y=0.09
c66 24 VSS 1.65079e-19 $X=0.801 $Y=0.09
c67 22 VSS 0.0178177f $X=0.866 $Y=0.2295
c68 19 VSS 3.14771e-19 $X=0.881 $Y=0.2295
c69 17 VSS 2.67274e-19 $X=0.808 $Y=0.2295
c70 13 VSS 0.020153f $X=0.81 $Y=0.0405
c71 9 VSS 6.29543e-19 $X=0.827 $Y=0.0405
c72 2 VSS 0.0580179f $X=0.729 $Y=0.0405
r73 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.819
+ $Y=0.09 $X2=0.828 $Y2=0.09
r74 54 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.09 $X2=0.828 $Y2=0.09
r75 53 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.09 $X2=0.819 $Y2=0.09
r76 49 50 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.167 $X2=0.837 $Y2=0.207
r77 48 49 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.165 $X2=0.837 $Y2=0.167
r78 47 48 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.14 $X2=0.837 $Y2=0.165
r79 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.122 $X2=0.837 $Y2=0.14
r80 45 46 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.101 $X2=0.837 $Y2=0.122
r81 44 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.207
r82 43 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.09
r83 43 45 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.101
r84 41 42 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.062 $X2=0.81 $Y2=0.0715
r85 38 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.054 $X2=0.81 $Y2=0.062
r86 36 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.09
r87 36 42 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.0715
r88 31 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r89 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.81 $Y2=0.234
r90 29 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.09 $X2=0.7965 $Y2=0.09
r91 27 29 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.09 $X2=0.792 $Y2=0.09
r92 27 28 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.747 $Y=0.09 $X2=0.747
+ $Y2=0.09
r93 24 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.81 $Y2=0.09
r94 24 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.7965 $Y2=0.09
r95 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2295 $X2=0.866 $Y2=0.2295
r96 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.808
+ $Y=0.2295 $X2=0.866 $Y2=0.2295
r97 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.234 $X2=0.81
+ $Y2=0.234
r98 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2295 $X2=0.808 $Y2=0.2295
r99 13 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.054 $X2=0.81
+ $Y2=0.054
r100 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.0405 $X2=0.81 $Y2=0.0405
r101 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.0405 $X2=0.81 $Y2=0.0405
r102 5 28 16.3636 $w=2.2e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.09 $X2=0.747 $Y2=0.09
r103 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.09 $X2=0.729 $Y2=0.2295
r104 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0405 $X2=0.729 $Y2=0.09
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%11 2 5 7 9 14 17 21 22 25 30 31 33 34 37 39 40 43
+ 44 45 46 48 50 51 52 53 54 55 56 59 61 62 64 VSS
c72 64 VSS 1.00092e-19 $X=0.693 $Y=0.131
c73 61 VSS 9.09188e-19 $X=0.72 $Y=0.131
c74 59 VSS 6.42979e-19 $X=0.783 $Y=0.131
c75 56 VSS 1.82087e-19 $X=0.693 $Y=0.216
c76 55 VSS 1.40959e-19 $X=0.693 $Y=0.207
c77 54 VSS 1.07888e-19 $X=0.693 $Y=0.189
c78 53 VSS 1.66071e-19 $X=0.693 $Y=0.171
c79 52 VSS 2.71272e-19 $X=0.693 $Y=0.165
c80 51 VSS 3.53682e-19 $X=0.693 $Y=0.153
c81 50 VSS 2.11704e-19 $X=0.693 $Y=0.225
c82 48 VSS 4.15228e-19 $X=0.693 $Y=0.114
c83 47 VSS 2.7378e-19 $X=0.693 $Y=0.106
c84 46 VSS 5.46003e-20 $X=0.693 $Y=0.099
c85 45 VSS 5.96385e-20 $X=0.693 $Y=0.081
c86 43 VSS 1.65771e-19 $X=0.693 $Y=0.062
c87 42 VSS 2.30403e-19 $X=0.693 $Y=0.122
c88 40 VSS 0.00145015f $X=0.6665 $Y=0.036
c89 39 VSS 0.00201121f $X=0.649 $Y=0.036
c90 37 VSS 0.00303728f $X=0.648 $Y=0.036
c91 34 VSS 0.00412969f $X=0.684 $Y=0.036
c92 33 VSS 0.00297725f $X=0.649 $Y=0.234
c93 32 VSS 2.2805e-19 $X=0.612 $Y=0.234
c94 31 VSS 0.00126734f $X=0.609 $Y=0.234
c95 30 VSS 0.0016591f $X=0.595 $Y=0.234
c96 25 VSS 0.00558865f $X=0.684 $Y=0.234
c97 24 VSS 5.62656e-19 $X=0.594 $Y=0.2295
c98 21 VSS 0.00254121f $X=0.594 $Y=0.2025
c99 18 VSS 1.02475e-19 $X=0.5895 $Y=0.216
c100 16 VSS 5.70081e-19 $X=0.648 $Y=0.0405
c101 10 VSS 7.61325e-20 $X=0.6435 $Y=0.054
c102 5 VSS 0.00241128f $X=0.783 $Y=0.131
c103 2 VSS 0.0591782f $X=0.783 $Y=0.0405
r104 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.131 $X2=0.738 $Y2=0.131
r105 59 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.131 $X2=0.738 $Y2=0.131
r106 57 64 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.693 $Y2=0.131
r107 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.72 $Y2=0.131
r108 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.207 $X2=0.693 $Y2=0.216
r109 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.189 $X2=0.693 $Y2=0.207
r110 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.171 $X2=0.693 $Y2=0.189
r111 52 53 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.165 $X2=0.693 $Y2=0.171
r112 51 52 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.153 $X2=0.693 $Y2=0.165
r113 50 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.225 $X2=0.693 $Y2=0.216
r114 49 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.131
r115 49 51 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.153
r116 47 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.106 $X2=0.693 $Y2=0.114
r117 46 47 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.099 $X2=0.693 $Y2=0.106
r118 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.081 $X2=0.693 $Y2=0.099
r119 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.063 $X2=0.693 $Y2=0.081
r120 43 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.062 $X2=0.693 $Y2=0.063
r121 42 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.131
r122 42 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.114
r123 41 43 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.045 $X2=0.693 $Y2=0.062
r124 39 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.649
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r125 36 39 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.649 $Y2=0.036
r126 36 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r127 34 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.036 $X2=0.693 $Y2=0.045
r128 34 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r129 32 33 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.649 $Y2=0.234
r130 31 32 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.609
+ $Y=0.234 $X2=0.612 $Y2=0.234
r131 30 31 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.595
+ $Y=0.234 $X2=0.609 $Y2=0.234
r132 27 30 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.595 $Y2=0.234
r133 25 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.234 $X2=0.693 $Y2=0.225
r134 25 33 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.234 $X2=0.649 $Y2=0.234
r135 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2295 $X2=0.594 $Y2=0.2295
r136 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r137 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.594 $Y2=0.2295
r138 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.5895 $Y2=0.189
r139 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.189 $X2=0.5895 $Y2=0.189
r140 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r141 13 37 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r142 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.648 $Y2=0.0405
r143 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.6435 $Y2=0.081
r144 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.081 $X2=0.6435 $Y2=0.081
r145 5 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.131 $X2=0.783
+ $Y2=0.131
r146 5 7 369.03 $w=2e-08 $l=9.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.131 $X2=0.783 $Y2=0.2295
r147 2 5 339.058 $w=2e-08 $l=9.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.131
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%12 2 5 7 9 12 14 17 21 25 26 30 31 35 36 37 43 VSS
c33 43 VSS 0.00419842f $X=1.098 $Y=0.234
c34 42 VSS 0.00204425f $X=1.107 $Y=0.234
c35 37 VSS 0.00106194f $X=1.107 $Y=0.171
c36 36 VSS 0.00114954f $X=1.107 $Y=0.117
c37 35 VSS 0.00158518f $X=1.107 $Y=0.225
c38 33 VSS 7.70286e-19 $X=1.073 $Y=0.036
c39 32 VSS 4.41014e-19 $X=1.066 $Y=0.036
c40 31 VSS 0.00146362f $X=1.062 $Y=0.036
c41 30 VSS 0.00481311f $X=1.044 $Y=0.036
c42 26 VSS 0.00226308f $X=1.008 $Y=0.036
c43 25 VSS 0.00460331f $X=1.098 $Y=0.036
c44 21 VSS 7.16657e-19 $X=0.999 $Y=0.105
c45 17 VSS 0.00426839f $X=1.078 $Y=0.2295
c46 12 VSS 0.00485453f $X=1.078 $Y=0.0405
c47 5 VSS 0.00233254f $X=0.999 $Y=0.1055
c48 2 VSS 0.0590816f $X=0.999 $Y=0.0405
r49 43 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r50 42 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r51 39 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.098 $Y2=0.234
r52 36 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.117 $X2=1.107 $Y2=0.171
r53 35 42 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.234
r54 35 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.171
r55 34 36 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.045 $X2=1.107 $Y2=0.117
r56 32 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.066
+ $Y=0.036 $X2=1.073 $Y2=0.036
r57 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=1.062
+ $Y=0.036 $X2=1.066 $Y2=0.036
r58 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=1.062 $Y2=0.036
r59 28 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.036 $X2=1.073 $Y2=0.036
r60 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.008
+ $Y=0.036 $X2=1.044 $Y2=0.036
r61 25 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.098 $Y=0.036 $X2=1.107 $Y2=0.045
r62 25 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.036 $X2=1.08 $Y2=0.036
r63 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.999 $Y=0.045 $X2=1.008 $Y2=0.036
r64 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.045 $X2=0.999 $Y2=0.105
r65 17 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234 $X2=1.08
+ $Y2=0.234
r66 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2295 $X2=1.078 $Y2=0.2295
r67 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.036 $X2=1.08
+ $Y2=0.036
r68 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.0405 $X2=1.078 $Y2=0.0405
r69 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.105 $X2=0.999
+ $Y2=0.105
r70 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.1055 $X2=0.999 $Y2=0.2295
r71 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.0405 $X2=0.999 $Y2=0.1055
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%13 2 7 10 15 18 21 23 25 26 29 30 31 34 35 40 41
+ 43 46 47 48 49 51 54 55 58 68 73 76 78 79 86 VSS
c79 86 VSS 0.00317836f $X=1.269 $Y=0.136
c80 79 VSS 0.00160638f $X=1.229 $Y=0.153
c81 78 VSS 0.00791219f $X=1.175 $Y=0.153
c82 76 VSS 0.00438571f $X=1.269 $Y=0.153
c83 73 VSS 1.90597e-19 $X=0.945 $Y=0.153
c84 68 VSS 0.0033916f $X=0.936 $Y=0.234
c85 67 VSS 0.00253671f $X=0.945 $Y=0.234
c86 58 VSS 4.04001e-19 $X=1.053 $Y=0.14
c87 55 VSS 3.26354e-19 $X=1.008 $Y=0.162
c88 54 VSS 0.00199114f $X=0.99 $Y=0.162
c89 52 VSS 0.0023929f $X=1.044 $Y=0.162
c90 51 VSS 0.00104404f $X=0.945 $Y=0.225
c91 49 VSS 2.07499e-19 $X=0.945 $Y=0.136
c92 48 VSS 2.77769e-19 $X=0.945 $Y=0.119
c93 47 VSS 2.61356e-19 $X=0.945 $Y=0.101
c94 46 VSS 6.393e-19 $X=0.945 $Y=0.081
c95 45 VSS 3.04212e-19 $X=0.945 $Y=0.153
c96 43 VSS 0.00136569f $X=0.92 $Y=0.036
c97 42 VSS 4.8751e-19 $X=0.904 $Y=0.036
c98 41 VSS 0.00146362f $X=0.9 $Y=0.036
c99 40 VSS 0.00358427f $X=0.882 $Y=0.036
c100 35 VSS 0.00347893f $X=0.936 $Y=0.036
c101 34 VSS 0.00276615f $X=0.918 $Y=0.2295
c102 30 VSS 5.63046e-19 $X=0.935 $Y=0.2295
c103 29 VSS 0.0201056f $X=0.864 $Y=0.0405
c104 25 VSS 5.63046e-19 $X=0.881 $Y=0.0405
c105 21 VSS 0.00431818f $X=1.323 $Y=0.136
c106 18 VSS 0.0615048f $X=1.323 $Y=0.0675
c107 10 VSS 0.0581342f $X=1.269 $Y=0.0675
c108 5 VSS 0.00302777f $X=1.053 $Y=0.14
c109 2 VSS 0.0627731f $X=1.053 $Y=0.0405
r110 78 79 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=1.175
+ $Y=0.153 $X2=1.229 $Y2=0.153
r111 76 79 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.269
+ $Y=0.153 $X2=1.229 $Y2=0.153
r112 76 86 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.269 $Y=0.153 $X2=1.269
+ $Y2=0.153
r113 72 78 15.6173 $w=1.8e-08 $l=2.3e-07 $layer=M2 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=1.175 $Y2=0.153
r114 72 73 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.945 $Y=0.153 $X2=0.945
+ $Y2=0.153
r115 68 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r116 67 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r117 64 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.234 $X2=0.936 $Y2=0.234
r118 56 58 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.153 $X2=1.053 $Y2=0.14
r119 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.99
+ $Y=0.162 $X2=1.008 $Y2=0.162
r120 53 73 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.945 $Y2=0.162
r121 53 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.99 $Y2=0.162
r122 52 56 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.162 $X2=1.053 $Y2=0.153
r123 52 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.162 $X2=1.008 $Y2=0.162
r124 51 67 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.234
r125 50 73 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.162
r126 50 51 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.225
r127 48 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.119 $X2=0.945 $Y2=0.136
r128 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.101 $X2=0.945 $Y2=0.119
r129 46 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.081 $X2=0.945 $Y2=0.101
r130 45 73 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.162
r131 45 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.136
r132 44 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.081
r133 42 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.904
+ $Y=0.036 $X2=0.92 $Y2=0.036
r134 41 42 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.036 $X2=0.904 $Y2=0.036
r135 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r136 37 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r137 35 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r138 35 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.92 $Y2=0.036
r139 34 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.234
+ $X2=0.918 $Y2=0.234
r140 31 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.2295 $X2=0.918 $Y2=0.2295
r141 30 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.935 $Y=0.2295 $X2=0.918 $Y2=0.2295
r142 29 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036
+ $X2=0.864 $Y2=0.036
r143 26 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.864 $Y2=0.0405
r144 25 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0405 $X2=0.864 $Y2=0.0405
r145 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.136 $X2=1.323 $Y2=0.2025
r146 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.0675 $X2=1.323 $Y2=0.136
r147 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.269
+ $Y=0.136 $X2=1.323 $Y2=0.136
r148 13 86 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.269 $Y=0.136 $X2=1.269
+ $Y2=0.136
r149 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.136 $X2=1.269 $Y2=0.2025
r150 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.0675 $X2=1.269 $Y2=0.136
r151 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.053 $Y=0.14 $X2=1.053
+ $Y2=0.14
r152 5 7 335.312 $w=2e-08 $l=8.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.14 $X2=1.053 $Y2=0.2295
r153 2 5 372.777 $w=2e-08 $l=9.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.0405 $X2=1.053 $Y2=0.14
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%14 1 4 6 11 14 21 23 24 25 VSS
c29 26 VSS 0.00225803f $X=0.485 $Y=0.234
c30 25 VSS 0.0014167f $X=0.461 $Y=0.234
c31 24 VSS 0.0134342f $X=0.447 $Y=0.234
c32 23 VSS 0.00523898f $X=0.309 $Y=0.234
c33 21 VSS 0.00168783f $X=0.486 $Y=0.234
c34 14 VSS 0.0195485f $X=0.542 $Y=0.2025
c35 11 VSS 3.25039e-19 $X=0.557 $Y=0.2025
c36 9 VSS 4.57278e-19 $X=0.484 $Y=0.2025
c37 4 VSS 0.00250857f $X=0.272 $Y=0.2025
c38 1 VSS 3.31752e-19 $X=0.287 $Y=0.2025
r39 25 26 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.461
+ $Y=0.234 $X2=0.485 $Y2=0.234
r40 24 25 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.234 $X2=0.461 $Y2=0.234
r41 23 24 9.37037 $w=1.8e-08 $l=1.38e-07 $layer=M1 $thickness=3.6e-08 $X=0.309
+ $Y=0.234 $X2=0.447 $Y2=0.234
r42 21 26 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.485 $Y2=0.234
r43 17 23 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.309 $Y2=0.234
r44 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.542 $Y2=0.2025
r45 9 14 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.484
+ $Y=0.2025 $X2=0.542 $Y2=0.2025
r46 9 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r47 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.2025 $X2=0.484 $Y2=0.2025
r48 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r49 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.272 $Y2=0.2025
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%16 1 2 5 6 7 10 12 18 20 21 22 23 24 25 VSS
c21 25 VSS 3.8923e-20 $X=0.423 $Y=0.198
c22 24 VSS 8.46035e-21 $X=0.414 $Y=0.198
c23 23 VSS 0.00116854f $X=0.396 $Y=0.198
c24 22 VSS 0.00134991f $X=0.379 $Y=0.198
c25 21 VSS 8.46035e-21 $X=0.36 $Y=0.198
c26 20 VSS 2.61077e-19 $X=0.342 $Y=0.198
c27 18 VSS 3.31089e-19 $X=0.432 $Y=0.198
c28 12 VSS 5.44897e-19 $X=0.324 $Y=0.198
c29 10 VSS 0.00631853f $X=0.432 $Y=0.2025
c30 6 VSS 5.67296e-19 $X=0.449 $Y=0.2025
c31 5 VSS 0.00790786f $X=0.324 $Y=0.2025
c32 1 VSS 6.05629e-19 $X=0.341 $Y=0.2025
r33 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.423 $Y2=0.198
r34 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.414 $Y2=0.198
r35 22 23 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.198 $X2=0.396 $Y2=0.198
r36 21 22 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.198 $X2=0.379 $Y2=0.198
r37 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r38 18 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.423 $Y2=0.198
r39 12 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.342 $Y2=0.198
r40 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r41 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r42 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r43 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198 $X2=0.324
+ $Y2=0.198
r44 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
r45 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%QN 1 2 6 7 10 11 14 16 24 26 VSS
c14 26 VSS 0.00603734f $X=1.377 $Y=0.2
c15 25 VSS 0.0025598f $X=1.377 $Y=0.09
c16 24 VSS 0.00130995f $X=1.379 $Y=0.223
c17 16 VSS 0.0146181f $X=1.368 $Y=0.234
c18 14 VSS 0.0097377f $X=1.296 $Y=0.036
c19 11 VSS 0.0144374f $X=1.368 $Y=0.036
c20 10 VSS 0.0101615f $X=1.296 $Y=0.2025
c21 6 VSS 5.72268e-19 $X=1.313 $Y=0.2025
c22 1 VSS 5.72268e-19 $X=1.313 $Y=0.0675
r23 25 26 7.46914 $w=1.8e-08 $l=1.1e-07 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.09 $X2=1.377 $Y2=0.2
r24 24 26 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.223 $X2=1.377 $Y2=0.2
r25 22 24 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.225 $X2=1.377 $Y2=0.223
r26 21 25 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.045 $X2=1.377 $Y2=0.09
r27 16 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.368 $Y=0.234 $X2=1.377 $Y2=0.225
r28 16 18 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.368
+ $Y=0.234 $X2=1.296 $Y2=0.234
r29 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.036 $X2=1.296
+ $Y2=0.036
r30 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.368 $Y=0.036 $X2=1.377 $Y2=0.045
r31 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.368
+ $Y=0.036 $X2=1.296 $Y2=0.036
r32 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.234 $X2=1.296
+ $Y2=0.234
r33 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.279 $Y=0.2025 $X2=1.296 $Y2=0.2025
r34 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.313 $Y=0.2025 $X2=1.296 $Y2=0.2025
r35 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.296
+ $Y=0.0675 $X2=1.296 $Y2=0.036
r36 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.279
+ $Y=0.0675 $X2=1.296 $Y2=0.0675
r37 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.313
+ $Y=0.0675 $X2=1.296 $Y2=0.0675
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%19 1 6 9 VSS
c10 9 VSS 0.0140217f $X=0.704 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.719 $Y=0.2295
c12 4 VSS 2.70811e-19 $X=0.646 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.646
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.631
+ $Y=0.2295 $X2=0.646 $Y2=0.2295
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%20 1 6 9 VSS
c9 9 VSS 0.0145746f $X=0.974 $Y=0.0405
c10 6 VSS 3.14771e-19 $X=0.989 $Y=0.0405
c11 4 VSS 2.65708e-19 $X=0.916 $Y=0.0405
r12 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r13 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.916
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r14 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.901
+ $Y=0.0405 $X2=0.916 $Y2=0.0405
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%22 1 2 VSS
c2 1 VSS 0.00203573f $X=0.719 $Y=0.0405
r3 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0405 $X2=0.685 $Y2=0.0405
.ends

.subckt PM_SDFHX2_ASAP7_75T_SRAM%23 1 2 VSS
c0 1 VSS 0.00214045f $X=0.989 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.2295 $X2=0.955 $Y2=0.2295
.ends


* END of "./SDFHx2_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt SDFHx2_ASAP7_75t_SRAM  VSS VDD CLK SE D SI QN
* 
* QN	QN
* SI	SI
* D	D
* SE	SE
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_9_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_SE_M2_g noxref_15 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 noxref_21 N_6_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 noxref_17 N_D_M4_g noxref_21 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 noxref_15 N_SI_M5_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 N_11_M6_d N_4_M6_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M7 N_22_M7_d N_9_M7_g N_11_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M8 VSS N_10_M8_g N_22_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.027
M9 N_10_M9_d N_11_M9_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_13_M10_d N_9_M10_g N_10_M10_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.827 $Y=0.027
M11 N_20_M11_d N_4_M11_g N_13_M11_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.027
M12 VSS N_12_M12_g N_20_M12_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.027
M13 N_12_M13_d N_13_M13_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.027
M14 VSS N_SE_M14_g N_6_M14_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.205
+ $Y=0.027
M15 N_QN_M15_d N_13_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M16 N_QN_M16_d N_13_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.027
M17 VDD N_CLK_M17_g N_4_M17_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M18 N_9_M18_d N_4_M18_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M19 N_16_M19_d N_SE_M19_g N_14_M19_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M20 VDD N_6_M20_g N_16_M20_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M21 N_16_M21_d N_D_M21_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M22 N_14_M22_d N_SI_M22_g N_16_M22_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M23 N_11_M23_d N_9_M23_g N_14_M23_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M24 N_19_M24_d N_4_M24_g N_11_M24_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.611 $Y=0.216
M25 VDD N_10_M25_g N_19_M25_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.216
M26 N_10_M26_d N_11_M26_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M27 N_13_M27_d N_4_M27_g N_10_M27_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.216
M28 N_23_M28_d N_9_M28_g N_13_M28_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.935 $Y=0.216
M29 VDD N_12_M29_g N_23_M29_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.216
M30 N_12_M30_d N_13_M30_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.216
M31 VDD N_SE_M31_g N_6_M31_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.205
+ $Y=0.216
M32 N_QN_M32_d N_13_M32_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
M33 N_QN_M33_d N_13_M33_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.162
*
* 
* .include "SDFHx2_ASAP7_75t_SRAM.pex.sp.SDFHX2_ASAP7_75T_SRAM.pxi"
* BEGIN of "./SDFHx2_ASAP7_75t_SRAM.pex.sp.SDFHX2_ASAP7_75T_SRAM.pxi"
* File: SDFHx2_ASAP7_75t_SRAM.pex.sp.SDFHX2_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 13:03:25 2017
* 
x_PM_SDFHX2_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M17_g N_CLK_c_3_p CLK
+ N_CLK_c_9_p N_CLK_c_7_p N_CLK_c_19_p VSS PM_SDFHX2_ASAP7_75T_SRAM%CLK
x_PM_SDFHX2_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_21_n N_4_M18_g N_4_M6_g N_4_c_41_p
+ N_4_M24_g N_4_M11_g N_4_c_45_p N_4_M27_g N_4_M0_s N_4_c_22_n N_4_M17_s
+ N_4_c_23_n N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_54_p N_4_c_35_p
+ N_4_c_28_n N_4_c_58_p N_4_c_29_n N_4_c_56_p N_4_c_32_p N_4_c_36_p N_4_c_46_p
+ N_4_c_34_p N_4_c_64_p N_4_c_31_n N_4_c_48_p VSS PM_SDFHX2_ASAP7_75T_SRAM%4
x_PM_SDFHX2_ASAP7_75T_SRAM%SE N_SE_M2_g N_SE_c_90_p N_SE_M19_g N_SE_M14_g
+ N_SE_c_126_p N_SE_M31_g N_SE_c_95_p N_SE_c_140_p N_SE_c_138_p N_SE_c_156_p
+ N_SE_c_86_n SE N_SE_c_85_n N_SE_c_91_p N_SE_c_92_p N_SE_c_87_n N_SE_c_88_n
+ N_SE_c_136_p N_SE_c_104_p N_SE_c_108_p N_SE_c_93_p N_SE_c_137_p VSS
+ PM_SDFHX2_ASAP7_75T_SRAM%SE
x_PM_SDFHX2_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_168_n N_6_M20_g N_6_M14_s N_6_c_169_n
+ N_6_M31_s N_6_c_198_p N_6_c_205_p N_6_c_215_p N_6_c_202_p N_6_c_211_p
+ N_6_c_219_p N_6_c_171_n N_6_c_164_n N_6_c_186_p N_6_c_166_n N_6_c_174_n
+ N_6_c_177_n N_6_c_178_n N_6_c_204_p VSS PM_SDFHX2_ASAP7_75T_SRAM%6
x_PM_SDFHX2_ASAP7_75T_SRAM%D N_D_M4_g N_D_c_236_n N_D_M21_g D VSS
+ PM_SDFHX2_ASAP7_75T_SRAM%D
x_PM_SDFHX2_ASAP7_75T_SRAM%SI N_SI_M5_g N_SI_M22_g SI N_SI_c_256_n VSS
+ PM_SDFHX2_ASAP7_75T_SRAM%SI
x_PM_SDFHX2_ASAP7_75T_SRAM%9 N_9_c_278_n N_9_M23_g N_9_M7_g N_9_c_346_p N_9_M10_g
+ N_9_c_330_p N_9_c_282_n N_9_M28_g N_9_M1_d N_9_c_287_n N_9_M18_d N_9_c_288_n
+ N_9_c_289_n N_9_c_314_n N_9_c_301_n N_9_c_272_n N_9_c_374_p N_9_c_292_n
+ N_9_c_273_n N_9_c_295_n N_9_c_274_n N_9_c_298_n N_9_c_275_n N_9_c_276_n
+ N_9_c_299_n N_9_c_300_n N_9_c_277_n VSS PM_SDFHX2_ASAP7_75T_SRAM%9
x_PM_SDFHX2_ASAP7_75T_SRAM%10 N_10_M8_g N_10_M25_g N_10_M10_s N_10_M9_d
+ N_10_c_397_n N_10_M26_d N_10_c_410_n N_10_M27_s N_10_c_412_n N_10_c_400_n
+ N_10_c_401_n N_10_c_398_n N_10_c_394_n N_10_c_403_n N_10_c_399_n N_10_c_427_p
+ N_10_c_441_p N_10_c_395_n N_10_c_429_p N_10_c_396_n N_10_c_417_n N_10_c_418_n
+ N_10_c_404_n VSS PM_SDFHX2_ASAP7_75T_SRAM%10
x_PM_SDFHX2_ASAP7_75T_SRAM%11 N_11_M9_g N_11_c_443_n N_11_M26_g N_11_M6_d N_11_M7_s
+ N_11_M23_d N_11_c_444_n N_11_M24_s N_11_c_507_p N_11_c_466_n N_11_c_467_n
+ N_11_c_445_n N_11_c_453_n N_11_c_454_n N_11_c_455_n N_11_c_456_n N_11_c_457_n
+ N_11_c_490_n N_11_c_459_n N_11_c_460_n N_11_c_447_n N_11_c_510_p N_11_c_448_n
+ N_11_c_449_n N_11_c_472_n N_11_c_474_n N_11_c_477_n N_11_c_511_p N_11_c_482_n
+ N_11_c_451_n N_11_c_452_n N_11_c_486_n VSS PM_SDFHX2_ASAP7_75T_SRAM%11
x_PM_SDFHX2_ASAP7_75T_SRAM%12 N_12_M12_g N_12_c_536_p N_12_M29_g N_12_M13_d
+ N_12_c_521_n N_12_M30_d N_12_c_523_n N_12_c_515_n N_12_c_516_n N_12_c_517_n
+ N_12_c_518_n N_12_c_519_n N_12_c_527_n N_12_c_520_n N_12_c_530_n N_12_c_545_p
+ VSS PM_SDFHX2_ASAP7_75T_SRAM%12
x_PM_SDFHX2_ASAP7_75T_SRAM%13 N_13_M13_g N_13_M30_g N_13_M15_g N_13_M32_g
+ N_13_M16_g N_13_c_554_n N_13_M33_g N_13_M11_s N_13_M10_d N_13_c_555_n
+ N_13_M28_s N_13_M27_d N_13_c_579_n N_13_c_556_n N_13_c_557_n N_13_c_547_n
+ N_13_c_559_n N_13_c_560_n N_13_c_568_n N_13_c_549_n N_13_c_581_n N_13_c_582_n
+ N_13_c_625_p N_13_c_602_n N_13_c_604_n N_13_c_569_n N_13_c_550_n N_13_c_561_n
+ N_13_c_551_n N_13_c_563_n N_13_c_565_n VSS PM_SDFHX2_ASAP7_75T_SRAM%13
x_PM_SDFHX2_ASAP7_75T_SRAM%14 N_14_M19_s N_14_c_627_n N_14_M22_d N_14_M23_s
+ N_14_c_626_n N_14_c_633_n N_14_c_628_n N_14_c_630_n N_14_c_634_n VSS
+ PM_SDFHX2_ASAP7_75T_SRAM%14
x_PM_SDFHX2_ASAP7_75T_SRAM%16 N_16_M20_s N_16_M19_d N_16_c_669_n N_16_M22_s
+ N_16_M21_d N_16_c_671_n N_16_c_661_n N_16_c_660_n N_16_c_663_n N_16_c_655_n
+ N_16_c_665_n N_16_c_666_n N_16_c_657_n N_16_c_659_n VSS
+ PM_SDFHX2_ASAP7_75T_SRAM%16
x_PM_SDFHX2_ASAP7_75T_SRAM%QN N_QN_M16_d N_QN_M15_d N_QN_M33_d N_QN_M32_d
+ N_QN_c_680_n N_QN_c_676_n N_QN_c_684_n N_QN_c_677_n QN N_QN_c_688_n VSS
+ PM_SDFHX2_ASAP7_75T_SRAM%QN
x_PM_SDFHX2_ASAP7_75T_SRAM%19 N_19_M24_d N_19_M25_s N_19_c_691_n VSS
+ PM_SDFHX2_ASAP7_75T_SRAM%19
x_PM_SDFHX2_ASAP7_75T_SRAM%20 N_20_M11_d N_20_M12_s N_20_c_700_n VSS
+ PM_SDFHX2_ASAP7_75T_SRAM%20
x_PM_SDFHX2_ASAP7_75T_SRAM%22 N_22_M8_s N_22_M7_d VSS PM_SDFHX2_ASAP7_75T_SRAM%22
x_PM_SDFHX2_ASAP7_75T_SRAM%23 N_23_M29_s N_23_M28_d VSS PM_SDFHX2_ASAP7_75T_SRAM%23
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_CLK_c_2_p N_4_c_21_n 0.00105598f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_CLK_c_3_p N_4_c_22_n 2.66516e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.054
cc_4 N_CLK_c_3_p N_4_c_23_n 0.0012473f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.144
cc_5 N_CLK_c_3_p N_4_c_24_n 3.97017e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.081
cc_6 N_CLK_c_3_p N_4_c_25_n 0.0012473f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.1125
cc_7 N_CLK_c_7_p N_4_c_26_n 0.00140648f $X=0.081 $Y=0.167 $X2=0.018 $Y2=0.2
cc_8 N_CLK_c_3_p N_4_c_27_n 4.97741e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_9_p N_4_c_28_n 0.00123168f $X=0.081 $Y=0.162 $X2=0.033 $Y2=0.153
cc_10 N_CLK_c_3_p N_4_c_29_n 5.36602e-19 $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_11 N_CLK_c_9_p N_4_c_29_n 8.66987e-19 $X=0.081 $Y=0.162 $X2=0.175 $Y2=0.153
cc_12 N_CLK_c_3_p N_4_c_31_n 0.00203815f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_13 N_CLK_c_3_p N_SE_c_85_n 2.45198e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2
cc_14 N_CLK_c_3_p N_9_c_272_n 6.32319e-19 $X=0.081 $Y=0.135 $X2=0.621 $Y2=0.135
cc_15 CLK N_9_c_273_n 3.23206e-19 $X=0.078 $Y=0.19 $X2=0.337 $Y2=0.153
cc_16 CLK N_9_c_274_n 2.57347e-19 $X=0.078 $Y=0.19 $X2=0.817 $Y2=0.153
cc_17 N_CLK_c_3_p N_9_c_275_n 0.00114506f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_18 N_CLK_c_3_p N_9_c_276_n 3.05593e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_19 N_CLK_c_19_p N_9_c_277_n 3.05593e-19 $X=0.081 $Y=0.1785 $X2=0 $Y2=0
cc_20 N_4_c_32_p N_SE_c_86_n 8.13669e-19 $X=0.337 $Y=0.153 $X2=0 $Y2=0
cc_21 N_4_c_32_p N_SE_c_87_n 0.0022834f $X=0.337 $Y=0.153 $X2=0 $Y2=0
cc_22 N_4_c_34_p N_SE_c_88_n 0.0022834f $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_23 N_4_c_35_p N_6_c_164_n 3.98881e-19 $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_24 N_4_c_36_p N_6_c_164_n 0.0176158f $X=0.479 $Y=0.153 $X2=0 $Y2=0
cc_25 N_4_c_36_p N_6_c_166_n 0.00114531f $X=0.479 $Y=0.153 $X2=0 $Y2=0
cc_26 N_4_c_36_p D 0.00102191f $X=0.479 $Y=0.153 $X2=0.081 $Y2=0.135
cc_27 N_4_c_34_p SI 0.00113575f $X=0.743 $Y=0.153 $X2=0.081 $Y2=0.135
cc_28 N_4_M6_g N_9_c_278_n 0.00365763f $X=0.621 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_29 N_4_c_41_p N_9_c_278_n 9.97803e-19 $X=0.621 $Y=0.135 $X2=0.081 $Y2=0.054
cc_30 N_4_M6_g N_9_M7_g 0.00355599f $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_4_M11_g N_9_M10_g 0.00355599f $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_32 N_4_M11_g N_9_c_282_n 0.00605856f $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.1785
cc_33 N_4_c_45_p N_9_c_282_n 0.00180656f $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.1785
cc_34 N_4_c_46_p N_9_c_282_n 5.51712e-19 $X=0.891 $Y=0.153 $X2=0.081 $Y2=0.1785
cc_35 N_4_c_34_p N_9_c_282_n 0.00168667f $X=0.743 $Y=0.153 $X2=0.081 $Y2=0.1785
cc_36 N_4_c_48_p N_9_c_282_n 0.00123876f $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.1785
cc_37 N_4_c_29_n N_9_c_287_n 2.18034e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_38 N_4_c_29_n N_9_c_288_n 2.58357e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_35_p N_9_c_289_n 0.00279251f $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_34_p N_9_c_289_n 9.87747e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_41 N_4_c_29_n N_9_c_272_n 3.93085e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_42 N_4_c_54_p N_9_c_292_n 2.66501e-19 $X=0.054 $Y=0.234 $X2=0 $Y2=0
cc_43 N_4_c_29_n N_9_c_292_n 4.19323e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_44 N_4_c_56_p N_9_c_273_n 2.46239e-19 $X=0.211 $Y=0.153 $X2=0 $Y2=0
cc_45 N_4_c_34_p N_9_c_295_n 2.46239e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_46 N_4_c_58_p N_9_c_274_n 3.80004e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_56_p N_9_c_274_n 0.0471484f $X=0.211 $Y=0.153 $X2=0 $Y2=0
cc_48 N_4_c_34_p N_9_c_298_n 2.81643e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_49 N_4_c_31_n N_9_c_299_n 0.00218805f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_50 N_4_c_56_p N_9_c_300_n 0.00116576f $X=0.211 $Y=0.153 $X2=0 $Y2=0
cc_51 N_4_M6_g N_10_M8_g 2.82885e-19 $X=0.621 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_52 N_4_c_64_p N_10_c_394_n 5.29207e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_53 N_4_c_48_p N_10_c_395_n 0.00318254f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_54 N_4_c_46_p N_10_c_396_n 0.00128311f $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_55 N_4_M11_g N_11_M9_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_56 N_4_c_45_p N_11_c_443_n 2.98891e-19 $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.135
cc_57 N_4_c_58_p N_11_c_444_n 3.24488e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_58 N_4_M6_g N_11_c_445_n 3.41974e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_59 N_4_c_58_p N_11_c_445_n 0.00102727f $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_60 N_4_c_35_p N_11_c_447_n 0.00133841f $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_61 N_4_c_34_p N_11_c_448_n 7.726e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_62 N_4_c_58_p N_11_c_449_n 8.63476e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_63 N_4_c_34_p N_11_c_449_n 5.92766e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_64 N_4_c_34_p N_11_c_451_n 3.70527e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_65 N_4_c_64_p N_11_c_452_n 3.70527e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_66 N_4_M11_g N_12_M12_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_67 N_4_M11_g N_13_c_547_n 3.18506e-19 $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_68 N_4_c_48_p N_13_c_547_n 4.09234e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_69 N_4_c_48_p N_13_c_549_n 0.00320381f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_70 N_4_c_48_p N_13_c_550_n 3.56772e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_71 N_4_c_46_p N_13_c_551_n 9.47997e-19 $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_72 N_4_c_36_p N_14_c_626_n 4.23942e-19 $X=0.479 $Y=0.153 $X2=0 $Y2=0
cc_73 N_SE_M2_g N_6_M3_g 0.00304756f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_74 N_SE_c_90_p N_6_c_168_n 0.00126421f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_75 N_SE_c_91_p N_6_c_169_n 2.11282e-19 $X=1.215 $Y=0.045 $X2=0.081 $Y2=0.135
cc_76 N_SE_c_92_p N_6_c_169_n 8.20809e-19 $X=1.215 $Y=0.045 $X2=0.081 $Y2=0.135
cc_77 N_SE_c_93_p N_6_c_171_n 3.53759e-19 $X=1.215 $Y=0.09 $X2=0 $Y2=0
cc_78 N_SE_c_88_n N_6_c_164_n 0.0680793f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_79 N_SE_c_95_p N_6_c_166_n 8.79603e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_80 N_SE_c_92_p N_6_c_174_n 0.00733801f $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_81 N_SE_c_88_n N_6_c_174_n 0.00103045f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_82 N_SE_c_93_p N_6_c_174_n 3.73635e-19 $X=1.215 $Y=0.09 $X2=0 $Y2=0
cc_83 N_SE_c_88_n N_6_c_177_n 2.46239e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_84 N_SE_c_86_n N_6_c_178_n 3.24594e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_85 N_SE_M2_g N_D_M4_g 2.13359e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_86 N_SE_c_85_n N_9_c_301_n 0.00266639f $X=0.225 $Y=0.045 $X2=0 $Y2=0
cc_87 N_SE_c_87_n N_9_c_301_n 4.45368e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_88 N_SE_c_104_p N_9_c_301_n 2.64176e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_89 N_SE_c_86_n N_9_c_274_n 4.53301e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_90 N_SE_c_87_n N_9_c_274_n 3.907e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_91 N_SE_c_104_p N_9_c_275_n 0.00292661f $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_92 N_SE_c_108_p N_9_c_276_n 0.00266639f $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_93 N_SE_c_86_n N_9_c_299_n 0.00266639f $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_94 N_SE_c_88_n N_10_c_397_n 4.38905e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_95 N_SE_c_88_n N_10_c_398_n 3.00479e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_96 N_SE_c_88_n N_10_c_399_n 7.16568e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_97 N_SE_c_88_n N_11_c_453_n 0.00113636f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_98 N_SE_c_88_n N_11_c_454_n 2.78297e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_99 N_SE_c_88_n N_11_c_455_n 5.99401e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_100 N_SE_c_88_n N_11_c_456_n 4.8504e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_101 N_SE_c_88_n N_11_c_457_n 4.65038e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_102 N_SE_c_88_n N_12_c_515_n 5.48108e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_103 N_SE_c_88_n N_12_c_516_n 0.00109158f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_104 N_SE_c_88_n N_12_c_517_n 5.50727e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_105 N_SE_c_88_n N_12_c_518_n 9.11285e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_106 N_SE_c_88_n N_12_c_519_n 4.62125e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_107 N_SE_c_88_n N_12_c_520_n 5.48546e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_108 N_SE_M14_g N_13_M15_g 0.00268443f $X=1.215 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_109 N_SE_M14_g N_13_M16_g 2.13359e-19 $X=1.215 $Y=0.0405 $X2=0.081 $Y2=0.162
cc_110 N_SE_c_126_p N_13_c_554_n 0.00114994f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_111 N_SE_c_88_n N_13_c_555_n 2.30689e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_112 N_SE_c_88_n N_13_c_556_n 9.08574e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_113 N_SE_c_88_n N_13_c_557_n 0.00124317f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_114 N_SE_c_88_n N_13_c_547_n 4.54245e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_115 N_SE_c_88_n N_13_c_559_n 4.39544e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_116 N_SE_c_88_n N_13_c_560_n 5.37888e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_117 N_SE_c_92_p N_13_c_561_n 3.26078e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_118 N_SE_c_88_n N_13_c_551_n 9.36021e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_119 N_SE_c_91_p N_13_c_563_n 9.36021e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_120 N_SE_c_136_p N_13_c_563_n 0.00114818f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_121 N_SE_c_137_p N_13_c_565_n 0.00409386f $X=1.215 $Y=0.113 $X2=0 $Y2=0
cc_122 N_SE_c_138_p N_14_c_627_n 2.31793e-19 $X=0.261 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_123 N_SE_M2_g N_14_c_628_n 3.83731e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_124 N_SE_c_140_p N_14_c_628_n 6.51345e-19 $X=0.258 $Y=0.135 $X2=0 $Y2=0
cc_125 VSS N_SE_c_85_n 2.40719e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.135
cc_126 VSS N_SE_c_87_n 5.30841e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.135
cc_127 VSS N_SE_c_104_p 9.86432e-19 $X=0.225 $Y=0.081 $X2=0.081 $Y2=0.135
cc_128 VSS N_SE_c_95_p 0.00129447f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_129 VSS N_SE_c_87_n 7.061e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_130 VSS N_SE_c_104_p 7.68051e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_131 VSS N_SE_c_85_n 8.44602e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.19
cc_132 VSS N_SE_c_87_n 5.36527e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.19
cc_133 VSS N_SE_c_88_n 0.00141783f $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.144
cc_134 VSS N_SE_c_88_n 2.35788e-19 $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.162
cc_135 VSS N_SE_c_87_n 6.93145e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.1785
cc_136 VSS N_SE_c_88_n 9.13621e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_137 VSS N_SE_c_88_n 4.6862e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_138 VSS N_SE_c_88_n 5.41611e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_139 VSS N_SE_c_88_n 8.51044e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_140 VSS N_SE_c_156_p 0.00129447f $X=0.279 $Y=0.135 $X2=0 $Y2=0
cc_141 VSS N_SE_c_87_n 3.48715e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_142 VSS N_SE_c_108_p 9.77595e-19 $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_143 VSS N_SE_c_88_n 2.40178e-19 $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.135
cc_144 VSS N_SE_c_88_n 6.42719e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_145 VSS N_SE_c_88_n 0.00110738f $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.162
cc_146 N_SE_c_92_p N_QN_c_676_n 8.29488e-19 $X=1.215 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_147 N_SE_c_88_n N_20_c_700_n 4.98441e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_148 N_6_M3_g N_D_M4_g 0.00304756f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_149 N_6_c_168_n N_D_c_236_n 9.71463e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_150 N_6_c_164_n D 3.33994e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_151 N_6_c_166_n D 0.00195518f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_152 N_6_c_178_n D 9.77589e-19 $X=0.351 $Y=0.126 $X2=0 $Y2=0
cc_153 N_6_M3_g N_SI_M5_g 2.48122e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_154 N_6_c_164_n SI 3.40688e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_155 N_6_c_186_p N_9_c_282_n 3.37164e-19 $X=0.936 $Y=0.081 $X2=0.891 $Y2=0.135
cc_156 N_6_c_164_n N_9_c_274_n 0.0011956f $X=0.9 $Y=0.081 $X2=0.817 $Y2=0.153
cc_157 N_6_c_164_n N_10_c_400_n 5.04077e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_158 N_6_c_164_n N_10_c_401_n 2.53924e-19 $X=0.9 $Y=0.081 $X2=0.056 $Y2=0.054
cc_159 N_6_c_164_n N_10_c_398_n 8.29294e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_160 N_6_c_164_n N_10_c_403_n 5.75824e-19 $X=0.9 $Y=0.081 $X2=0.018 $Y2=0.144
cc_161 N_6_c_164_n N_10_c_404_n 7.91051e-19 $X=0.9 $Y=0.081 $X2=0.047 $Y2=0.234
cc_162 N_6_c_164_n N_11_c_454_n 4.20387e-19 $X=0.9 $Y=0.081 $X2=0.018 $Y2=0.081
cc_163 N_6_c_164_n N_11_c_459_n 4.92006e-19 $X=0.9 $Y=0.081 $X2=0.054 $Y2=0.036
cc_164 N_6_c_164_n N_11_c_460_n 7.19039e-19 $X=0.9 $Y=0.081 $X2=0.054 $Y2=0.036
cc_165 N_6_c_169_n N_12_c_521_n 0.00124414f $X=1.19 $Y=0.0405 $X2=0.621
+ $Y2=0.135
cc_166 N_6_c_171_n N_12_c_521_n 2.40393e-19 $X=1.161 $Y=0.081 $X2=0.621
+ $Y2=0.135
cc_167 N_6_c_198_p N_12_c_523_n 5.25714e-19 $X=1.19 $Y=0.2295 $X2=0.891
+ $Y2=0.0405
cc_168 N_6_c_171_n N_12_c_515_n 9.95523e-19 $X=1.161 $Y=0.081 $X2=0.891
+ $Y2=0.135
cc_169 N_6_c_169_n N_12_c_516_n 3.43147e-19 $X=1.19 $Y=0.0405 $X2=0.071
+ $Y2=0.054
cc_170 N_6_c_174_n N_12_c_516_n 0.00251979f $X=1.161 $Y=0.049 $X2=0.071
+ $Y2=0.054
cc_171 N_6_c_202_p N_12_c_527_n 0.00251979f $X=1.17 $Y=0.234 $X2=0.018 $Y2=0.045
cc_172 N_6_c_171_n N_12_c_520_n 0.0012739f $X=1.161 $Y=0.081 $X2=0.018 $Y2=0.144
cc_173 N_6_c_204_p N_12_c_520_n 0.00251979f $X=1.161 $Y=0.2125 $X2=0.018
+ $Y2=0.144
cc_174 N_6_c_205_p N_12_c_530_n 0.00251979f $X=1.161 $Y=0.225 $X2=0.018
+ $Y2=0.081
cc_175 N_6_c_186_p N_13_c_557_n 6.23859e-19 $X=0.936 $Y=0.081 $X2=0.018
+ $Y2=0.225
cc_176 N_6_c_171_n N_13_c_560_n 3.66836e-19 $X=1.161 $Y=0.081 $X2=0.054
+ $Y2=0.036
cc_177 N_6_c_171_n N_13_c_568_n 5.24665e-19 $X=1.161 $Y=0.081 $X2=0.047
+ $Y2=0.036
cc_178 N_6_c_186_p N_13_c_569_n 3.12147e-19 $X=0.936 $Y=0.081 $X2=0.135
+ $Y2=0.153
cc_179 N_6_c_169_n N_13_c_551_n 2.50315e-19 $X=1.19 $Y=0.0405 $X2=0.891
+ $Y2=0.153
cc_180 N_6_c_211_p N_13_c_551_n 3.14624e-19 $X=1.179 $Y=0.234 $X2=0.891
+ $Y2=0.153
cc_181 N_6_c_171_n N_13_c_551_n 0.00815696f $X=1.161 $Y=0.081 $X2=0.891
+ $Y2=0.153
cc_182 N_6_c_174_n N_13_c_551_n 0.00110082f $X=1.161 $Y=0.049 $X2=0.891
+ $Y2=0.153
cc_183 N_6_c_198_p N_13_c_563_n 2.19627e-19 $X=1.19 $Y=0.2295 $X2=0.743
+ $Y2=0.153
cc_184 N_6_c_215_p N_13_c_563_n 3.14624e-19 $X=1.188 $Y=0.234 $X2=0.743
+ $Y2=0.153
cc_185 N_6_M3_g N_14_c_630_n 2.37298e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_186 VSS N_6_c_164_n 3.90811e-19 $X=0.9 $Y=0.081 $X2=0.621 $Y2=0.135
cc_187 VSS N_6_c_177_n 7.35661e-19 $X=0.351 $Y=0.099 $X2=0.621 $Y2=0.135
cc_188 VSS N_6_c_219_p 6.42252e-19 $X=0.351 $Y=0.081 $X2=0.621 $Y2=0.2295
cc_189 VSS N_6_c_219_p 0.00369658f $X=0.351 $Y=0.081 $X2=0.891 $Y2=0.135
cc_190 N_6_M3_g N_16_c_655_n 2.50526e-19 $X=0.351 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_191 N_6_c_166_n N_16_c_655_n 0.00110314f $X=0.351 $Y=0.135 $X2=0.891
+ $Y2=0.135
cc_192 VSS N_6_c_177_n 2.30452e-19 $X=0.351 $Y=0.099 $X2=0.135 $Y2=0.135
cc_193 VSS N_6_c_164_n 7.92007e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_194 VSS N_6_c_219_p 8.14481e-19 $X=0.351 $Y=0.081 $X2=0.891 $Y2=0.0405
cc_195 VSS N_6_c_164_n 2.67459e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_196 VSS N_6_c_164_n 3.16736e-19 $X=0.9 $Y=0.081 $X2=0.891 $Y2=0.135
cc_197 VSS N_6_c_164_n 2.43408e-19 $X=0.9 $Y=0.081 $X2=0.891 $Y2=0.135
cc_198 VSS N_6_c_164_n 5.19239e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_199 N_6_c_215_p N_QN_c_677_n 2.72644e-19 $X=1.188 $Y=0.234 $X2=0 $Y2=0
cc_200 N_6_c_186_p N_20_c_700_n 5.02041e-19 $X=0.936 $Y=0.081 $X2=0.621
+ $Y2=0.0675
cc_201 VSS N_6_c_219_p 2.73492e-19 $X=0.351 $Y=0.081 $X2=0.135 $Y2=0.054
cc_202 N_D_M4_g N_SI_M5_g 0.00348334f $X=0.405 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_203 D SI 7.00288e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_204 N_D_c_236_n N_SI_c_256_n 0.00109838f $X=0.405 $Y=0.135 $X2=0.621
+ $Y2=0.2295
cc_205 N_D_M4_g N_14_c_630_n 2.37298e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_206 VSS N_D_M4_g 3.08888e-19 $X=0.405 $Y=0.0675 $X2=0.891 $Y2=0.2295
cc_207 VSS D 5.77345e-19 $X=0.405 $Y=0.134 $X2=0.891 $Y2=0.2295
cc_208 N_D_M4_g N_16_c_657_n 2.43567e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_209 D N_16_c_657_n 0.00108212f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_210 D N_16_c_659_n 3.4434e-19 $X=0.405 $Y=0.134 $X2=0.071 $Y2=0.054
cc_211 VSS D 8.86227e-19 $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.135
cc_212 VSS D 0.00161923f $X=0.405 $Y=0.134 $X2=0.891 $Y2=0.0405
cc_213 N_SI_M5_g N_9_c_278_n 2.94371e-19 $X=0.459 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_214 N_SI_c_256_n N_9_c_278_n 5.18435e-19 $X=0.475 $Y=0.135 $X2=0.135
+ $Y2=0.054
cc_215 SI N_9_c_289_n 0.00114959f $X=0.473 $Y=0.135 $X2=0 $Y2=0
cc_216 SI N_9_c_314_n 0.00114959f $X=0.473 $Y=0.135 $X2=0.054 $Y2=0.234
cc_217 SI N_9_c_295_n 0.00239259f $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.153
cc_218 SI N_9_c_274_n 0.00167124f $X=0.473 $Y=0.135 $X2=0.817 $Y2=0.153
cc_219 SI N_14_c_626_n 0.00560919f $X=0.473 $Y=0.135 $X2=0.621 $Y2=0.2295
cc_220 SI N_14_c_633_n 0.00167456f $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.135
cc_221 N_SI_M5_g N_14_c_634_n 2.70361e-19 $X=0.459 $Y=0.0675 $X2=0.071 $Y2=0.054
cc_222 SI N_16_c_660_n 6.69571e-19 $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.0405
cc_223 VSS N_SI_M5_g 3.10987e-19 $X=0.459 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_224 VSS N_SI_c_256_n 2.08525e-19 $X=0.475 $Y=0.135 $X2=0.891 $Y2=0.135
cc_225 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.135
cc_226 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.2295
cc_227 VSS SI 0.00110314f $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.2295
cc_228 N_9_M7_g N_10_M8_g 0.00341068f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_229 N_9_M10_g N_10_M8_g 2.13359e-19 $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_230 N_9_c_282_n N_10_M8_g 0.00205997f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_231 N_9_c_298_n N_10_M8_g 3.19768e-19 $X=0.729 $Y=0.18 $X2=0.081 $Y2=0.054
cc_232 N_9_c_282_n N_10_c_397_n 5.52012e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_233 N_9_c_282_n N_10_c_410_n 2.12581e-19 $X=0.945 $Y=0.178 $X2=0.081
+ $Y2=0.144
cc_234 N_9_c_282_n N_10_M27_s 2.50995e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.167
cc_235 N_9_M10_g N_10_c_412_n 0.00200065f $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_236 N_9_c_282_n N_10_c_412_n 0.00322783f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_237 N_9_c_282_n N_10_c_394_n 3.41745e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_238 N_9_M10_g N_10_c_395_n 2.74825e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_239 N_9_M10_g N_10_c_396_n 2.10136e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_240 N_9_c_298_n N_10_c_417_n 6.73839e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_241 N_9_c_330_p N_10_c_418_n 0.00195059f $X=0.837 $Y=0.178 $X2=0 $Y2=0
cc_242 N_9_c_282_n N_10_c_418_n 0.00191847f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_243 N_9_M10_g N_10_c_404_n 3.61755e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_244 N_9_M7_g N_11_M9_g 2.13359e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_245 N_9_M10_g N_11_M9_g 0.00341068f $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_246 N_9_c_282_n N_11_M9_g 0.00302156f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_247 N_9_c_289_n N_11_c_444_n 7.70794e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_248 N_9_c_295_n N_11_c_444_n 0.001307f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_249 N_9_c_295_n N_11_c_466_n 0.00138499f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_250 N_9_c_274_n N_11_c_467_n 0.00160025f $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_251 N_9_M7_g N_11_c_453_n 4.38308e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_252 N_9_M7_g N_11_c_459_n 2.0845e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_253 N_9_M7_g N_11_c_460_n 2.27141e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_254 N_9_c_282_n N_11_c_449_n 0.0361494f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_255 N_9_c_282_n N_11_c_472_n 2.38252e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_256 N_9_c_298_n N_11_c_472_n 0.00386452f $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_257 N_9_c_346_p N_11_c_474_n 7.00743e-19 $X=0.675 $Y=0.178 $X2=0 $Y2=0
cc_258 N_9_c_282_n N_11_c_474_n 7.89771e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_259 N_9_c_274_n N_11_c_474_n 4.88732e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_260 N_9_M7_g N_11_c_477_n 2.5554e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_261 N_9_c_282_n N_11_c_477_n 3.47488e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_262 N_9_c_295_n N_11_c_477_n 2.13133e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_263 N_9_c_274_n N_11_c_477_n 4.32971e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_264 N_9_c_298_n N_11_c_477_n 2.60223e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_265 N_9_c_282_n N_11_c_482_n 4.26771e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_266 N_9_c_282_n N_11_c_451_n 4.41163e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_267 N_9_c_282_n N_11_c_452_n 3.33141e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_268 N_9_c_298_n N_11_c_452_n 9.1388e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_269 N_9_M7_g N_11_c_486_n 2.11651e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_270 N_9_c_282_n N_12_M12_g 0.00341068f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_271 N_9_c_282_n N_13_M13_g 2.13359e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_272 N_9_c_282_n N_13_c_555_n 8.27183e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_273 N_9_c_282_n N_13_M28_s 3.37661e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_274 N_9_c_282_n N_13_c_579_n 0.00145657f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_275 N_9_c_282_n N_13_c_568_n 3.13444e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_276 N_9_c_282_n N_13_c_581_n 2.6418e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_277 N_9_c_282_n N_13_c_582_n 0.00294656f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_278 N_9_c_282_n N_13_c_569_n 3.75802e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_279 N_9_c_282_n N_13_c_550_n 5.46321e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_280 N_9_c_288_n N_14_c_627_n 9.65806e-19 $X=0.16 $Y=0.216 $X2=0.081 $Y2=0.135
cc_281 N_9_c_274_n N_14_c_627_n 4.65646e-19 $X=0.729 $Y=0.189 $X2=0.081
+ $Y2=0.135
cc_282 N_9_c_300_n N_14_c_627_n 0.00109797f $X=0.189 $Y=0.164 $X2=0.081
+ $Y2=0.135
cc_283 N_9_c_289_n N_14_c_626_n 9.68946e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_284 N_9_c_274_n N_14_c_626_n 6.49405e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_285 N_9_c_374_p N_14_c_628_n 7.61293e-19 $X=0.189 $Y=0.234 $X2=0 $Y2=0
cc_286 N_9_c_274_n N_14_c_628_n 7.84624e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_287 N_9_c_274_n N_14_c_634_n 6.22262e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_288 VSS N_9_c_287_n 9.30745e-19 $X=0.16 $Y=0.054 $X2=0.081 $Y2=0.135
cc_289 N_9_c_274_n N_16_c_661_n 2.13751e-19 $X=0.729 $Y=0.189 $X2=0.081
+ $Y2=0.135
cc_290 N_9_c_274_n N_16_c_660_n 7.1298e-19 $X=0.729 $Y=0.189 $X2=0.081 $Y2=0.162
cc_291 N_9_c_274_n N_16_c_663_n 6.46208e-19 $X=0.729 $Y=0.189 $X2=0.081
+ $Y2=0.1785
cc_292 N_9_c_274_n N_16_c_655_n 4.50553e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_293 N_9_c_274_n N_16_c_665_n 4.86474e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_294 N_9_c_274_n N_16_c_666_n 4.60071e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_295 N_9_c_274_n N_16_c_657_n 4.38038e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_296 N_9_c_274_n N_16_c_659_n 2.31538e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_297 VSS N_9_c_278_n 3.33061e-19 $X=0.567 $Y=0.1355 $X2=0 $Y2=0
cc_298 VSS N_9_c_289_n 0.00110314f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_299 N_9_c_282_n N_19_M25_s 2.33161e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.216
cc_300 N_9_M7_g N_19_c_691_n 0.00248549f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_301 N_9_c_282_n N_19_c_691_n 0.00208457f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_302 N_9_c_274_n N_19_c_691_n 7.88525e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_303 N_9_c_282_n N_20_c_700_n 0.00250239f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_304 N_10_M8_g N_11_M9_g 0.00268443f $X=0.729 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_305 N_10_c_398_n N_11_M9_g 3.7702e-19 $X=0.792 $Y=0.09 $X2=0.135 $Y2=0.054
cc_306 N_10_c_399_n N_11_c_457_n 2.46574e-19 $X=0.81 $Y=0.054 $X2=0.027
+ $Y2=0.036
cc_307 N_10_c_400_n N_11_c_490_n 0.00360624f $X=0.747 $Y=0.09 $X2=0.054
+ $Y2=0.036
cc_308 N_10_c_401_n N_11_c_459_n 3.99428e-19 $X=0.747 $Y=0.09 $X2=0.054
+ $Y2=0.036
cc_309 N_10_c_396_n N_11_c_448_n 2.22221e-19 $X=0.837 $Y=0.165 $X2=0.054
+ $Y2=0.234
cc_310 N_10_c_427_p N_11_c_477_n 2.22221e-19 $X=0.837 $Y=0.225 $X2=0.0505
+ $Y2=0.234
cc_311 N_10_c_398_n N_11_c_482_n 0.00205899f $X=0.792 $Y=0.09 $X2=0.621
+ $Y2=0.135
cc_312 N_10_c_429_p N_11_c_482_n 7.38434e-19 $X=0.837 $Y=0.14 $X2=0.621
+ $Y2=0.135
cc_313 N_10_M8_g N_11_c_452_n 3.21351e-19 $X=0.729 $Y=0.0405 $X2=0.033 $Y2=0.153
cc_314 N_10_c_400_n N_11_c_452_n 0.00205899f $X=0.747 $Y=0.09 $X2=0.033
+ $Y2=0.153
cc_315 N_10_c_397_n N_13_c_555_n 0.00379158f $X=0.81 $Y=0.0405 $X2=0 $Y2=0
cc_316 N_10_c_399_n N_13_c_555_n 2.84891e-19 $X=0.81 $Y=0.054 $X2=0 $Y2=0
cc_317 N_10_c_404_n N_13_c_555_n 2.08929e-19 $X=0.837 $Y=0.09 $X2=0 $Y2=0
cc_318 N_10_c_412_n N_13_c_579_n 0.00222825f $X=0.866 $Y=0.2295 $X2=0 $Y2=0
cc_319 N_10_c_397_n N_13_c_557_n 3.41768e-19 $X=0.81 $Y=0.0405 $X2=0.018
+ $Y2=0.225
cc_320 N_10_c_404_n N_13_c_568_n 4.2911e-19 $X=0.837 $Y=0.09 $X2=0.047 $Y2=0.036
cc_321 N_10_c_418_n N_13_c_582_n 4.2911e-19 $X=0.837 $Y=0.207 $X2=0.054
+ $Y2=0.234
cc_322 N_10_c_412_n N_13_c_569_n 3.64454e-19 $X=0.866 $Y=0.2295 $X2=0.135
+ $Y2=0.153
cc_323 N_10_c_394_n N_13_c_569_n 4.86017e-19 $X=0.828 $Y=0.234 $X2=0.135
+ $Y2=0.153
cc_324 N_10_c_441_p N_13_c_550_n 4.2911e-19 $X=0.837 $Y=0.101 $X2=0.211
+ $Y2=0.153
cc_325 N_11_c_444_n N_14_c_626_n 0.00424458f $X=0.594 $Y=0.2025 $X2=0.621
+ $Y2=0.2295
cc_326 N_11_c_466_n N_14_c_626_n 4.3429e-19 $X=0.595 $Y=0.234 $X2=0.621
+ $Y2=0.2295
cc_327 N_11_c_466_n N_14_c_633_n 2.8677e-19 $X=0.595 $Y=0.234 $X2=0.891
+ $Y2=0.135
cc_328 VSS N_11_c_444_n 0.0016174f $X=0.594 $Y=0.2025 $X2=0.621 $Y2=0.0675
cc_329 VSS N_11_c_454_n 0.00414127f $X=0.648 $Y=0.036 $X2=0.621 $Y2=0.0675
cc_330 VSS N_11_c_455_n 3.30384e-19 $X=0.649 $Y=0.036 $X2=0.621 $Y2=0.0675
cc_331 VSS N_11_c_454_n 2.79363e-19 $X=0.648 $Y=0.036 $X2=0 $Y2=0
cc_332 VSS N_11_c_459_n 2.70508e-19 $X=0.693 $Y=0.081 $X2=0 $Y2=0
cc_333 N_11_c_444_n N_19_c_691_n 0.00167238f $X=0.594 $Y=0.2025 $X2=0.621
+ $Y2=0.0675
cc_334 N_11_c_507_p N_19_c_691_n 0.00315491f $X=0.684 $Y=0.234 $X2=0.621
+ $Y2=0.0675
cc_335 N_11_c_445_n N_19_c_691_n 0.00111131f $X=0.649 $Y=0.234 $X2=0.621
+ $Y2=0.0675
cc_336 N_11_c_454_n N_19_c_691_n 5.67227e-19 $X=0.648 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_337 N_11_c_510_p N_19_c_691_n 4.0515e-19 $X=0.693 $Y=0.225 $X2=0.621
+ $Y2=0.0675
cc_338 N_11_c_511_p N_19_c_691_n 0.0409693f $X=0.693 $Y=0.216 $X2=0.621
+ $Y2=0.0675
cc_339 N_11_c_453_n N_22_M8_s 2.44135e-19 $X=0.684 $Y=0.036 $X2=0.135 $Y2=0.054
cc_340 N_11_c_457_n N_22_M8_s 3.62465e-19 $X=0.693 $Y=0.062 $X2=0.135 $Y2=0.054
cc_341 N_12_M12_g N_13_M13_g 0.00268443f $X=0.999 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_342 N_12_c_519_n N_13_M13_g 3.55314e-19 $X=1.062 $Y=0.036 $X2=0.135 $Y2=0.054
cc_343 N_12_c_517_n N_13_c_556_n 0.00136796f $X=1.008 $Y=0.036 $X2=0.018
+ $Y2=0.045
cc_344 N_12_c_515_n N_13_c_560_n 0.00136796f $X=0.999 $Y=0.105 $X2=0.054
+ $Y2=0.036
cc_345 N_12_c_536_p N_13_c_568_n 3.34766e-19 $X=0.999 $Y=0.1055 $X2=0.047
+ $Y2=0.036
cc_346 N_12_c_515_n N_13_c_568_n 0.00136796f $X=0.999 $Y=0.105 $X2=0.047
+ $Y2=0.036
cc_347 N_12_c_527_n N_13_c_582_n 5.28703e-19 $X=1.107 $Y=0.225 $X2=0.054
+ $Y2=0.234
cc_348 N_12_M12_g N_13_c_602_n 6.35734e-19 $X=0.999 $Y=0.0405 $X2=0.0505
+ $Y2=0.234
cc_349 N_12_c_515_n N_13_c_602_n 7.99759e-19 $X=0.999 $Y=0.105 $X2=0.0505
+ $Y2=0.234
cc_350 N_12_c_519_n N_13_c_604_n 2.75024e-19 $X=1.062 $Y=0.036 $X2=0.621
+ $Y2=0.135
cc_351 N_12_c_530_n N_13_c_604_n 0.00266666f $X=1.107 $Y=0.171 $X2=0.621
+ $Y2=0.135
cc_352 N_12_c_523_n N_13_c_551_n 2.19627e-19 $X=1.078 $Y=0.2295 $X2=0.891
+ $Y2=0.153
cc_353 N_12_c_530_n N_13_c_551_n 0.00106087f $X=1.107 $Y=0.171 $X2=0.891
+ $Y2=0.153
cc_354 N_12_c_545_p N_13_c_551_n 5.80975e-19 $X=1.098 $Y=0.234 $X2=0.891
+ $Y2=0.153
cc_355 N_12_c_517_n N_20_c_700_n 5.06067e-19 $X=1.008 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_356 N_13_c_554_n N_QN_M16_d 3.7444e-19 $X=1.323 $Y=0.136 $X2=0.135 $Y2=0.054
cc_357 N_13_c_554_n N_QN_M33_d 3.85232e-19 $X=1.323 $Y=0.136 $X2=0.135 $Y2=0.216
cc_358 N_13_c_554_n N_QN_c_680_n 8.43851e-19 $X=1.323 $Y=0.136 $X2=0.621
+ $Y2=0.0675
cc_359 N_13_c_565_n N_QN_c_680_n 0.00132451f $X=1.269 $Y=0.136 $X2=0.621
+ $Y2=0.0675
cc_360 N_13_M16_g N_QN_c_676_n 4.61823e-19 $X=1.323 $Y=0.0675 $X2=0 $Y2=0
cc_361 N_13_c_554_n N_QN_c_676_n 5.30021e-19 $X=1.323 $Y=0.136 $X2=0 $Y2=0
cc_362 N_13_c_554_n N_QN_c_684_n 7.60428e-19 $X=1.323 $Y=0.136 $X2=0.621
+ $Y2=0.2295
cc_363 N_13_c_565_n N_QN_c_684_n 6.27401e-19 $X=1.269 $Y=0.136 $X2=0.621
+ $Y2=0.2295
cc_364 N_13_M16_g N_QN_c_677_n 4.56718e-19 $X=1.323 $Y=0.0675 $X2=0 $Y2=0
cc_365 N_13_c_554_n N_QN_c_677_n 5.38938e-19 $X=1.323 $Y=0.136 $X2=0 $Y2=0
cc_366 N_13_c_554_n N_QN_c_688_n 3.64608e-19 $X=1.323 $Y=0.136 $X2=0.056
+ $Y2=0.054
cc_367 N_13_c_565_n N_QN_c_688_n 0.00122416f $X=1.269 $Y=0.136 $X2=0.056
+ $Y2=0.054
cc_368 N_13_c_555_n N_20_c_700_n 0.00210698f $X=0.864 $Y=0.0405 $X2=0.621
+ $Y2=0.0675
cc_369 N_13_c_556_n N_20_c_700_n 0.00203632f $X=0.936 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_370 N_13_c_559_n N_20_c_700_n 0.00129774f $X=0.92 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_371 N_13_c_560_n N_20_c_700_n 0.00104094f $X=0.945 $Y=0.081 $X2=0.621
+ $Y2=0.0675
cc_372 N_13_c_625_p N_20_c_700_n 2.5109e-19 $X=0.99 $Y=0.162 $X2=0.621
+ $Y2=0.0675
cc_373 VSS N_14_c_627_n 0.00156967f $X=0.272 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_374 VSS N_14_c_626_n 0.00145555f $X=0.542 $Y=0.2025 $X2=0.891 $Y2=0.0405
cc_375 N_14_c_627_n N_16_c_669_n 0.003872f $X=0.272 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_376 N_14_c_630_n N_16_c_669_n 0.00248801f $X=0.447 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_377 N_14_c_626_n N_16_c_671_n 0.00434154f $X=0.542 $Y=0.2025 $X2=0.621
+ $Y2=0.0675
cc_378 N_14_c_630_n N_16_c_671_n 0.0025506f $X=0.447 $Y=0.234 $X2=0.621
+ $Y2=0.0675
cc_379 N_14_c_627_n N_16_c_661_n 3.19827e-19 $X=0.272 $Y=0.2025 $X2=0.621
+ $Y2=0.135
cc_380 N_14_c_630_n N_16_c_661_n 0.0113176f $X=0.447 $Y=0.234 $X2=0.621
+ $Y2=0.135
cc_381 VSS N_14_c_626_n 4.53012e-19 $X=0.542 $Y=0.2025 $X2=0 $Y2=0
cc_382 VSS N_16_c_671_n 0.00141703f $X=0.432 $Y=0.2025 $X2=0.135 $Y2=0.135

* END of "./SDFHx2_ASAP7_75t_SRAM.pex.sp.SDFHX2_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: SDFHx3_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 13:03:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "SDFHx3_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./SDFHx3_ASAP7_75t_SRAM.pex.sp.pex"
* File: SDFHx3_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 13:03:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_SDFHX3_ASAP7_75T_SRAM%CLK 2 5 7 11 16 18 19 20 VSS
c19 20 VSS 1.17072e-19 $X=0.081 $Y=0.1785
c20 19 VSS 3.55344e-20 $X=0.081 $Y=0.167
c21 18 VSS 9.34089e-20 $X=0.081 $Y=0.162
c22 16 VSS 0.00100628f $X=0.078 $Y=0.19
c23 11 VSS 0.00681069f $X=0.081 $Y=0.135
c24 5 VSS 0.00208806f $X=0.081 $Y=0.135
c25 2 VSS 0.0627545f $X=0.081 $Y=0.054
r26 19 20 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.167 $X2=0.081 $Y2=0.1785
r27 18 19 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.162 $X2=0.081 $Y2=0.167
r28 17 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.144 $X2=0.081 $Y2=0.162
r29 16 20 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.19 $X2=0.081 $Y2=0.1785
r30 11 17 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.144
r31 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r32 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r33 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%4 2 5 7 10 13 15 18 21 23 25 28 30 36 37 38 41 45
+ 52 59 64 71 72 73 74 75 77 79 80 84 92 VSS
c65 111 VSS 1.06551e-19 $X=0.03 $Y=0.153
c66 110 VSS 6.89947e-19 $X=0.027 $Y=0.153
c67 92 VSS 0.001222f $X=0.891 $Y=0.135
c68 84 VSS 0.00111816f $X=0.135 $Y=0.135
c69 80 VSS 0.00209834f $X=0.817 $Y=0.153
c70 79 VSS 0.00159119f $X=0.743 $Y=0.153
c71 77 VSS 0.00277988f $X=0.891 $Y=0.153
c72 75 VSS 0.0014306f $X=0.479 $Y=0.153
c73 74 VSS 0.00120845f $X=0.337 $Y=0.153
c74 73 VSS 9.39788e-19 $X=0.211 $Y=0.153
c75 72 VSS 0.00665478f $X=0.175 $Y=0.153
c76 71 VSS 9.40943e-19 $X=0.621 $Y=0.153
c77 64 VSS 6.72589e-19 $X=0.033 $Y=0.153
c78 59 VSS 5.26559e-19 $X=0.621 $Y=0.135
c79 55 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c80 54 VSS 0.00180216f $X=0.047 $Y=0.234
c81 52 VSS 0.00253483f $X=0.054 $Y=0.234
c82 50 VSS 0.00305101f $X=0.027 $Y=0.234
c83 48 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c84 47 VSS 0.00199699f $X=0.047 $Y=0.036
c85 45 VSS 0.00239525f $X=0.054 $Y=0.036
c86 43 VSS 0.00305101f $X=0.027 $Y=0.036
c87 42 VSS 5.16336e-19 $X=0.018 $Y=0.2125
c88 41 VSS 0.00180713f $X=0.018 $Y=0.2
c89 40 VSS 4.96914e-19 $X=0.018 $Y=0.225
c90 38 VSS 0.00159315f $X=0.018 $Y=0.1125
c91 37 VSS 0.00142827f $X=0.018 $Y=0.081
c92 36 VSS 0.00143809f $X=0.018 $Y=0.144
c93 33 VSS 0.0049466f $X=0.056 $Y=0.216
c94 30 VSS 2.98509e-19 $X=0.071 $Y=0.216
c95 28 VSS 0.00460164f $X=0.056 $Y=0.054
c96 25 VSS 2.98509e-19 $X=0.071 $Y=0.054
c97 21 VSS 0.00216055f $X=0.891 $Y=0.135
c98 18 VSS 0.0585656f $X=0.891 $Y=0.0405
c99 13 VSS 0.00201785f $X=0.621 $Y=0.135
c100 10 VSS 0.0601628f $X=0.621 $Y=0.0675
c101 5 VSS 0.00199564f $X=0.135 $Y=0.135
c102 2 VSS 0.0630095f $X=0.135 $Y=0.054
r103 110 111 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r104 107 110 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r105 79 80 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.743
+ $Y=0.153 $X2=0.817 $Y2=0.153
r106 77 80 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.817 $Y2=0.153
r107 77 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r108 74 75 9.64198 $w=1.8e-08 $l=1.42e-07 $layer=M2 $thickness=3.6e-08 $X=0.337
+ $Y=0.153 $X2=0.479 $Y2=0.153
r109 73 74 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.211
+ $Y=0.153 $X2=0.337 $Y2=0.153
r110 72 73 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.175
+ $Y=0.153 $X2=0.211 $Y2=0.153
r111 70 79 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.743 $Y2=0.153
r112 70 75 9.64198 $w=1.8e-08 $l=1.42e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.479 $Y2=0.153
r113 70 71 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.621 $Y=0.153 $X2=0.621
+ $Y2=0.153
r114 67 72 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.153 $X2=0.175 $Y2=0.153
r115 67 84 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.135 $Y=0.153 $X2=0.135
+ $Y2=0.153
r116 64 111 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r117 63 67 6.92593 $w=1.8e-08 $l=1.02e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.135 $Y2=0.153
r118 63 64 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r119 59 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.153
r120 54 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r121 52 55 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r122 50 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r123 47 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r124 45 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r125 43 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r126 41 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r127 40 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r128 40 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r129 39 107 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r130 39 41 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.2
r131 37 38 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.1125
r132 36 107 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r133 36 38 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1125
r134 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r135 35 37 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r136 33 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r137 30 33 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r138 28 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r139 25 28 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r140 21 92 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.135 $X2=0.891
+ $Y2=0.135
r141 21 23 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.135 $X2=0.891 $Y2=0.2295
r142 18 21 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.0405 $X2=0.891 $Y2=0.135
r143 13 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r144 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2295
r145 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r146 5 84 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r147 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r148 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%SE 2 5 7 10 13 15 19 22 23 24 31 33 41 44 45 46 47
+ 54 58 59 62 63 VSS
c79 63 VSS 2.09605e-19 $X=1.215 $Y=0.113
c80 62 VSS 0.00202057f $X=1.215 $Y=0.09
c81 59 VSS 2.63823e-19 $X=0.225 $Y=0.099
c82 58 VSS 5.90201e-19 $X=0.225 $Y=0.081
c83 54 VSS 0.00128643f $X=1.215 $Y=0.136
c84 47 VSS 0.0383019f $X=1.175 $Y=0.045
c85 46 VSS 0.00642311f $X=0.337 $Y=0.045
c86 45 VSS 0.00700571f $X=1.215 $Y=0.045
c87 44 VSS 0.00307515f $X=1.215 $Y=0.045
c88 41 VSS 0.00531f $X=0.225 $Y=0.045
c89 31 VSS 0.00110873f $X=0.225 $Y=0.126
c90 24 VSS 2.51525e-19 $X=0.279 $Y=0.135
c91 23 VSS 1.48251e-19 $X=0.261 $Y=0.135
c92 22 VSS 6.38823e-20 $X=0.258 $Y=0.135
c93 21 VSS 0.00134071f $X=0.255 $Y=0.135
c94 19 VSS 6.89032e-19 $X=0.297 $Y=0.135
c95 13 VSS 0.00244398f $X=1.215 $Y=0.136
c96 10 VSS 0.0611074f $X=1.215 $Y=0.0405
c97 5 VSS 0.00319967f $X=0.297 $Y=0.135
c98 2 VSS 0.063344f $X=0.297 $Y=0.0675
r99 62 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.09 $X2=1.215 $Y2=0.113
r100 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.081 $X2=0.225 $Y2=0.099
r101 54 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.136 $X2=1.215 $Y2=0.113
r102 46 47 56.9012 $w=1.8e-08 $l=8.38e-07 $layer=M2 $thickness=3.6e-08 $X=0.337
+ $Y=0.045 $X2=1.175 $Y2=0.045
r103 45 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.215 $Y2=0.09
r104 44 47 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.175 $Y2=0.045
r105 44 45 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.215 $Y=0.045 $X2=1.215
+ $Y2=0.045
r106 41 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.081
r107 40 46 7.60494 $w=1.8e-08 $l=1.12e-07 $layer=M2 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.337 $Y2=0.045
r108 40 41 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.225 $Y=0.045 $X2=0.225
+ $Y2=0.045
r109 31 59 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.099
r110 31 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r111 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.135 $X2=0.279 $Y2=0.135
r112 22 23 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.258
+ $Y=0.135 $X2=0.261 $Y2=0.135
r113 21 22 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.255
+ $Y=0.135 $X2=0.258 $Y2=0.135
r114 19 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.279 $Y2=0.135
r115 17 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.225 $Y2=0.135
r116 17 21 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.255 $Y2=0.135
r117 13 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.215 $Y=0.136 $X2=1.215
+ $Y2=0.136
r118 13 15 350.298 $w=2e-08 $l=9.35e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.136 $X2=1.215 $Y2=0.2295
r119 10 13 357.791 $w=2e-08 $l=9.55e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.0405 $X2=1.215 $Y2=0.136
r120 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r121 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r122 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%6 2 5 7 9 12 14 17 23 26 28 29 33 36 38 39 43 51
+ 57 58 65 VSS
c69 65 VSS 3.36547e-19 $X=1.161 $Y=0.2125
c70 58 VSS 5.45782e-19 $X=0.351 $Y=0.126
c71 57 VSS 8.0335e-19 $X=0.351 $Y=0.099
c72 51 VSS 0.00325146f $X=1.161 $Y=0.049
c73 43 VSS 3.66031e-19 $X=0.351 $Y=0.135
c74 39 VSS 9.89222e-19 $X=0.936 $Y=0.081
c75 38 VSS 0.00685031f $X=0.9 $Y=0.081
c76 36 VSS 0.00169093f $X=1.161 $Y=0.081
c77 33 VSS 8.10983e-19 $X=0.351 $Y=0.081
c78 29 VSS 7.48824e-19 $X=1.179 $Y=0.234
c79 28 VSS 0.00240687f $X=1.17 $Y=0.234
c80 26 VSS 0.00328115f $X=1.188 $Y=0.234
c81 23 VSS 9.88154e-20 $X=1.161 $Y=0.225
c82 17 VSS 0.00404882f $X=1.19 $Y=0.2295
c83 14 VSS 2.95772e-19 $X=1.205 $Y=0.2295
c84 12 VSS 0.060801f $X=1.19 $Y=0.0405
c85 9 VSS 3.14771e-19 $X=1.205 $Y=0.0405
c86 5 VSS 0.00125227f $X=0.351 $Y=0.135
c87 2 VSS 0.0585837f $X=0.351 $Y=0.0675
r88 64 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.2 $X2=1.161 $Y2=0.2125
r89 57 58 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.099 $X2=0.351 $Y2=0.126
r90 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.161 $Y=0.049 $X2=1.161
+ $Y2=0.049
r91 43 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.126
r92 38 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.9
+ $Y=0.081 $X2=0.936 $Y2=0.081
r93 37 64 8.08025 $w=1.8e-08 $l=1.19e-07 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.2
r94 37 51 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.049
r95 36 39 15.2778 $w=1.8e-08 $l=2.25e-07 $layer=M2 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=0.936 $Y2=0.081
r96 36 37 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.161 $Y=0.081 $X2=1.161
+ $Y2=0.081
r97 33 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.099
r98 32 38 37.2778 $w=1.8e-08 $l=5.49e-07 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.9 $Y2=0.081
r99 32 33 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.081 $X2=0.351
+ $Y2=0.081
r100 28 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.17
+ $Y=0.234 $X2=1.179 $Y2=0.234
r101 26 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.188
+ $Y=0.234 $X2=1.179 $Y2=0.234
r102 23 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.225 $X2=1.161 $Y2=0.2125
r103 22 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.17 $Y2=0.234
r104 22 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.161 $Y2=0.225
r105 17 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.188 $Y=0.234
+ $X2=1.188 $Y2=0.234
r106 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.2295 $X2=1.19 $Y2=0.2295
r107 12 50 16.2355 $w=3.7e-08 $l=2.9e-08 $layer=LISD $thickness=2.8e-08 $X=1.19
+ $Y=0.0455 $X2=1.161 $Y2=0.0455
r108 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.0405 $X2=1.19 $Y2=0.0405
r109 5 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r110 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r111 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%D 2 5 7 11 VSS
c18 11 VSS 0.00145113f $X=0.405 $Y=0.134
c19 5 VSS 0.00106786f $X=0.405 $Y=0.135
c20 2 VSS 0.0589243f $X=0.405 $Y=0.0675
r21 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%SI 2 7 11 14 VSS
c21 14 VSS 0.0032805f $X=0.475 $Y=0.135
c22 11 VSS 0.0035781f $X=0.473 $Y=0.135
c23 2 VSS 0.0640988f $X=0.459 $Y=0.0675
r24 11 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.475 $Y=0.135 $X2=0.475
+ $Y2=0.135
r25 5 14 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.475 $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%9 2 5 8 11 14 17 20 23 37 40 42 45 49 53 58 60 67
+ 69 74 78 80 96 101 102 103 104 106 VSS
c121 108 VSS 7.92414e-20 $X=0.189 $Y=0.207
c122 106 VSS 2.53862e-19 $X=0.189 $Y=0.178
c123 105 VSS 3.91706e-20 $X=0.189 $Y=0.167
c124 104 VSS 6.6467e-19 $X=0.189 $Y=0.164
c125 103 VSS 3.3761e-19 $X=0.189 $Y=0.144
c126 102 VSS 4.92067e-19 $X=0.189 $Y=0.121
c127 101 VSS 8.32677e-19 $X=0.189 $Y=0.099
c128 96 VSS 6.49238e-19 $X=0.729 $Y=0.18
c129 80 VSS 0.0152374f $X=0.729 $Y=0.189
c130 78 VSS 0.0013748f $X=0.567 $Y=0.189
c131 74 VSS 6.28429e-19 $X=0.189 $Y=0.189
c132 69 VSS 0.00386366f $X=0.18 $Y=0.234
c133 68 VSS 4.87314e-19 $X=0.189 $Y=0.225
c134 67 VSS 0.00199636f $X=0.189 $Y=0.234
c135 60 VSS 0.00373046f $X=0.18 $Y=0.036
c136 58 VSS 0.00194932f $X=0.189 $Y=0.036
c137 53 VSS 9.61695e-20 $X=0.567 $Y=0.18
c138 49 VSS 5.76385e-19 $X=0.567 $Y=0.135
c139 45 VSS 0.00566559f $X=0.16 $Y=0.216
c140 40 VSS 0.0055918f $X=0.16 $Y=0.054
c141 20 VSS 0.108836f $X=0.945 $Y=0.178
c142 17 VSS 1.08457e-19 $X=0.837 $Y=0.178
c143 14 VSS 0.0600244f $X=0.837 $Y=0.0405
c144 11 VSS 2.24613e-19 $X=0.675 $Y=0.178
c145 8 VSS 0.0602569f $X=0.675 $Y=0.0405
c146 2 VSS 0.0660345f $X=0.567 $Y=0.1355
r147 107 108 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.2 $X2=0.189 $Y2=0.207
r148 105 106 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.167 $X2=0.189 $Y2=0.178
r149 104 105 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.167
r150 103 104 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.164
r151 102 103 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.121 $X2=0.189 $Y2=0.144
r152 101 102 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.099 $X2=0.189 $Y2=0.121
r153 95 96 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.729 $Y=0.18 $X2=0.729
+ $Y2=0.18
r154 80 96 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.729 $Y=0.189 $X2=0.729
+ $Y2=0.189
r155 77 80 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.729 $Y2=0.189
r156 77 78 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.567 $Y=0.189 $X2=0.567
+ $Y2=0.189
r157 74 107 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.2
r158 74 106 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.178
r159 73 77 25.6667 $w=1.8e-08 $l=3.78e-07 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.567 $Y2=0.189
r160 73 74 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.189 $X2=0.189
+ $Y2=0.189
r161 69 70 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r162 68 108 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.207
r163 67 70 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r164 67 68 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.189 $Y2=0.225
r165 64 69 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r166 60 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r167 59 101 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.099
r168 58 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r169 58 59 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r170 55 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r171 53 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.18 $X2=0.567 $Y2=0.189
r172 52 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.171 $X2=0.567 $Y2=0.18
r173 49 52 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.171
r174 45 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r175 42 45 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r176 40 55 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r177 37 40 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r178 20 23 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.178 $X2=0.945 $Y2=0.2295
r179 17 20 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08 $X=0.837
+ $Y=0.178 $X2=0.945 $Y2=0.178
r180 17 95 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08 $X=0.837
+ $Y=0.178 $X2=0.729 $Y2=0.178
r181 14 17 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0405 $X2=0.837 $Y2=0.178
r182 11 95 43.022 $w=2.6e-08 $l=5.4e-08 $layer=LISD $thickness=2.8e-08 $X=0.675
+ $Y=0.178 $X2=0.729 $Y2=0.178
r183 8 11 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.178
r184 2 49 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r185 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1355 $X2=0.567 $Y2=0.2025
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%10 2 7 9 10 13 14 17 19 22 27 28 29 31 36 38 44 45
+ 46 47 48 49 50 54 VSS
c49 56 VSS 5.19568e-19 $X=0.828 $Y=0.09
c50 55 VSS 4.09996e-19 $X=0.819 $Y=0.09
c51 54 VSS 4.29e-19 $X=0.837 $Y=0.09
c52 50 VSS 5.92866e-19 $X=0.837 $Y=0.207
c53 49 VSS 1.19762e-19 $X=0.837 $Y=0.167
c54 48 VSS 1.59501e-19 $X=0.837 $Y=0.165
c55 47 VSS 3.13056e-19 $X=0.837 $Y=0.14
c56 46 VSS 5.61414e-19 $X=0.837 $Y=0.122
c57 45 VSS 1.91116e-19 $X=0.837 $Y=0.101
c58 44 VSS 4.02479e-19 $X=0.837 $Y=0.225
c59 42 VSS 3.58124e-20 $X=0.81 $Y=0.0715
c60 38 VSS 0.00112276f $X=0.81 $Y=0.054
c61 31 VSS 0.00670205f $X=0.828 $Y=0.234
c62 30 VSS 4.74851e-19 $X=0.7965 $Y=0.09
c63 29 VSS 0.00125276f $X=0.792 $Y=0.09
c64 28 VSS 0.00410211f $X=0.747 $Y=0.09
c65 27 VSS 4.49532e-19 $X=0.747 $Y=0.09
c66 24 VSS 1.65079e-19 $X=0.801 $Y=0.09
c67 22 VSS 0.0178177f $X=0.866 $Y=0.2295
c68 19 VSS 3.14771e-19 $X=0.881 $Y=0.2295
c69 17 VSS 2.67274e-19 $X=0.808 $Y=0.2295
c70 13 VSS 0.020153f $X=0.81 $Y=0.0405
c71 9 VSS 6.29543e-19 $X=0.827 $Y=0.0405
c72 2 VSS 0.0580179f $X=0.729 $Y=0.0405
r73 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.819
+ $Y=0.09 $X2=0.828 $Y2=0.09
r74 54 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.09 $X2=0.828 $Y2=0.09
r75 53 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.09 $X2=0.819 $Y2=0.09
r76 49 50 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.167 $X2=0.837 $Y2=0.207
r77 48 49 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.165 $X2=0.837 $Y2=0.167
r78 47 48 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.14 $X2=0.837 $Y2=0.165
r79 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.122 $X2=0.837 $Y2=0.14
r80 45 46 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.101 $X2=0.837 $Y2=0.122
r81 44 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.207
r82 43 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.09
r83 43 45 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.101
r84 41 42 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.062 $X2=0.81 $Y2=0.0715
r85 38 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.054 $X2=0.81 $Y2=0.062
r86 36 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.09
r87 36 42 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.0715
r88 31 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r89 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.81 $Y2=0.234
r90 29 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.09 $X2=0.7965 $Y2=0.09
r91 27 29 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.09 $X2=0.792 $Y2=0.09
r92 27 28 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.747 $Y=0.09 $X2=0.747
+ $Y2=0.09
r93 24 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.81 $Y2=0.09
r94 24 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.7965 $Y2=0.09
r95 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2295 $X2=0.866 $Y2=0.2295
r96 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.808
+ $Y=0.2295 $X2=0.866 $Y2=0.2295
r97 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.234 $X2=0.81
+ $Y2=0.234
r98 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2295 $X2=0.808 $Y2=0.2295
r99 13 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.054 $X2=0.81
+ $Y2=0.054
r100 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.0405 $X2=0.81 $Y2=0.0405
r101 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.0405 $X2=0.81 $Y2=0.0405
r102 5 28 16.3636 $w=2.2e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.09 $X2=0.747 $Y2=0.09
r103 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.09 $X2=0.729 $Y2=0.2295
r104 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0405 $X2=0.729 $Y2=0.09
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%11 2 5 7 9 14 17 21 22 25 30 31 33 34 37 39 40 43
+ 44 45 46 48 50 51 52 53 54 55 56 59 61 62 64 VSS
c72 64 VSS 1.00092e-19 $X=0.693 $Y=0.131
c73 61 VSS 9.09188e-19 $X=0.72 $Y=0.131
c74 59 VSS 6.42979e-19 $X=0.783 $Y=0.131
c75 56 VSS 1.82087e-19 $X=0.693 $Y=0.216
c76 55 VSS 1.40959e-19 $X=0.693 $Y=0.207
c77 54 VSS 1.07888e-19 $X=0.693 $Y=0.189
c78 53 VSS 1.66071e-19 $X=0.693 $Y=0.171
c79 52 VSS 2.71272e-19 $X=0.693 $Y=0.165
c80 51 VSS 3.53682e-19 $X=0.693 $Y=0.153
c81 50 VSS 2.11704e-19 $X=0.693 $Y=0.225
c82 48 VSS 4.15228e-19 $X=0.693 $Y=0.114
c83 47 VSS 2.7378e-19 $X=0.693 $Y=0.106
c84 46 VSS 5.46003e-20 $X=0.693 $Y=0.099
c85 45 VSS 5.96385e-20 $X=0.693 $Y=0.081
c86 43 VSS 1.65771e-19 $X=0.693 $Y=0.062
c87 42 VSS 2.30403e-19 $X=0.693 $Y=0.122
c88 40 VSS 0.00145015f $X=0.6665 $Y=0.036
c89 39 VSS 0.00201121f $X=0.649 $Y=0.036
c90 37 VSS 0.00303728f $X=0.648 $Y=0.036
c91 34 VSS 0.00412969f $X=0.684 $Y=0.036
c92 33 VSS 0.00297725f $X=0.649 $Y=0.234
c93 32 VSS 2.2805e-19 $X=0.612 $Y=0.234
c94 31 VSS 0.00126734f $X=0.609 $Y=0.234
c95 30 VSS 0.0016591f $X=0.595 $Y=0.234
c96 25 VSS 0.00558865f $X=0.684 $Y=0.234
c97 24 VSS 5.62656e-19 $X=0.594 $Y=0.2295
c98 21 VSS 0.00254121f $X=0.594 $Y=0.2025
c99 18 VSS 1.02475e-19 $X=0.5895 $Y=0.216
c100 16 VSS 5.70081e-19 $X=0.648 $Y=0.0405
c101 10 VSS 7.61325e-20 $X=0.6435 $Y=0.054
c102 5 VSS 0.00241128f $X=0.783 $Y=0.131
c103 2 VSS 0.0591782f $X=0.783 $Y=0.0405
r104 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.131 $X2=0.738 $Y2=0.131
r105 59 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.131 $X2=0.738 $Y2=0.131
r106 57 64 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.693 $Y2=0.131
r107 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.72 $Y2=0.131
r108 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.207 $X2=0.693 $Y2=0.216
r109 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.189 $X2=0.693 $Y2=0.207
r110 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.171 $X2=0.693 $Y2=0.189
r111 52 53 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.165 $X2=0.693 $Y2=0.171
r112 51 52 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.153 $X2=0.693 $Y2=0.165
r113 50 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.225 $X2=0.693 $Y2=0.216
r114 49 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.131
r115 49 51 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.153
r116 47 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.106 $X2=0.693 $Y2=0.114
r117 46 47 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.099 $X2=0.693 $Y2=0.106
r118 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.081 $X2=0.693 $Y2=0.099
r119 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.063 $X2=0.693 $Y2=0.081
r120 43 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.062 $X2=0.693 $Y2=0.063
r121 42 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.131
r122 42 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.114
r123 41 43 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.045 $X2=0.693 $Y2=0.062
r124 39 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.649
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r125 36 39 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.649 $Y2=0.036
r126 36 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r127 34 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.036 $X2=0.693 $Y2=0.045
r128 34 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r129 32 33 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.649 $Y2=0.234
r130 31 32 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.609
+ $Y=0.234 $X2=0.612 $Y2=0.234
r131 30 31 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.595
+ $Y=0.234 $X2=0.609 $Y2=0.234
r132 27 30 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.595 $Y2=0.234
r133 25 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.234 $X2=0.693 $Y2=0.225
r134 25 33 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.234 $X2=0.649 $Y2=0.234
r135 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2295 $X2=0.594 $Y2=0.2295
r136 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r137 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.594 $Y2=0.2295
r138 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.5895 $Y2=0.189
r139 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.189 $X2=0.5895 $Y2=0.189
r140 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r141 13 37 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r142 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.648 $Y2=0.0405
r143 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.6435 $Y2=0.081
r144 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.081 $X2=0.6435 $Y2=0.081
r145 5 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.131 $X2=0.783
+ $Y2=0.131
r146 5 7 369.03 $w=2e-08 $l=9.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.131 $X2=0.783 $Y2=0.2295
r147 2 5 339.058 $w=2e-08 $l=9.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.131
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%12 2 5 7 9 12 14 17 21 25 26 30 31 35 36 37 43 VSS
c33 43 VSS 0.00419842f $X=1.098 $Y=0.234
c34 42 VSS 0.00204425f $X=1.107 $Y=0.234
c35 37 VSS 0.00106194f $X=1.107 $Y=0.171
c36 36 VSS 0.00114954f $X=1.107 $Y=0.117
c37 35 VSS 0.00158518f $X=1.107 $Y=0.225
c38 33 VSS 7.70286e-19 $X=1.073 $Y=0.036
c39 32 VSS 4.41014e-19 $X=1.066 $Y=0.036
c40 31 VSS 0.00146362f $X=1.062 $Y=0.036
c41 30 VSS 0.00481311f $X=1.044 $Y=0.036
c42 26 VSS 0.00226308f $X=1.008 $Y=0.036
c43 25 VSS 0.00460331f $X=1.098 $Y=0.036
c44 21 VSS 7.16657e-19 $X=0.999 $Y=0.105
c45 17 VSS 0.00426839f $X=1.078 $Y=0.2295
c46 12 VSS 0.00485453f $X=1.078 $Y=0.0405
c47 5 VSS 0.00233254f $X=0.999 $Y=0.1055
c48 2 VSS 0.0590816f $X=0.999 $Y=0.0405
r49 43 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r50 42 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r51 39 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.098 $Y2=0.234
r52 36 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.117 $X2=1.107 $Y2=0.171
r53 35 42 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.234
r54 35 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.171
r55 34 36 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.045 $X2=1.107 $Y2=0.117
r56 32 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.066
+ $Y=0.036 $X2=1.073 $Y2=0.036
r57 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=1.062
+ $Y=0.036 $X2=1.066 $Y2=0.036
r58 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=1.062 $Y2=0.036
r59 28 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.036 $X2=1.073 $Y2=0.036
r60 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.008
+ $Y=0.036 $X2=1.044 $Y2=0.036
r61 25 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.098 $Y=0.036 $X2=1.107 $Y2=0.045
r62 25 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.036 $X2=1.08 $Y2=0.036
r63 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.999 $Y=0.045 $X2=1.008 $Y2=0.036
r64 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.045 $X2=0.999 $Y2=0.105
r65 17 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234 $X2=1.08
+ $Y2=0.234
r66 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2295 $X2=1.078 $Y2=0.2295
r67 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.036 $X2=1.08
+ $Y2=0.036
r68 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.0405 $X2=1.078 $Y2=0.0405
r69 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.105 $X2=0.999
+ $Y2=0.105
r70 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.1055 $X2=0.999 $Y2=0.2295
r71 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.0405 $X2=0.999 $Y2=0.1055
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%13 2 7 10 15 18 23 26 29 31 33 34 37 38 39 42 43
+ 48 49 51 54 55 56 57 59 62 63 66 76 81 84 86 87 94 VSS
c81 94 VSS 0.00327387f $X=1.269 $Y=0.136
c82 87 VSS 0.00160638f $X=1.229 $Y=0.153
c83 86 VSS 0.00791219f $X=1.175 $Y=0.153
c84 84 VSS 0.00437729f $X=1.269 $Y=0.153
c85 81 VSS 1.90597e-19 $X=0.945 $Y=0.153
c86 76 VSS 0.0033916f $X=0.936 $Y=0.234
c87 75 VSS 0.00253671f $X=0.945 $Y=0.234
c88 66 VSS 4.04001e-19 $X=1.053 $Y=0.14
c89 63 VSS 3.26354e-19 $X=1.008 $Y=0.162
c90 62 VSS 0.00199114f $X=0.99 $Y=0.162
c91 60 VSS 0.0023929f $X=1.044 $Y=0.162
c92 59 VSS 0.00104404f $X=0.945 $Y=0.225
c93 57 VSS 2.07499e-19 $X=0.945 $Y=0.136
c94 56 VSS 2.77769e-19 $X=0.945 $Y=0.119
c95 55 VSS 2.61356e-19 $X=0.945 $Y=0.101
c96 54 VSS 6.393e-19 $X=0.945 $Y=0.081
c97 53 VSS 3.04212e-19 $X=0.945 $Y=0.153
c98 51 VSS 0.00136569f $X=0.92 $Y=0.036
c99 50 VSS 4.8751e-19 $X=0.904 $Y=0.036
c100 49 VSS 0.00146362f $X=0.9 $Y=0.036
c101 48 VSS 0.00358427f $X=0.882 $Y=0.036
c102 43 VSS 0.00347893f $X=0.936 $Y=0.036
c103 42 VSS 0.00276615f $X=0.918 $Y=0.2295
c104 38 VSS 5.63046e-19 $X=0.935 $Y=0.2295
c105 37 VSS 0.0201056f $X=0.864 $Y=0.0405
c106 33 VSS 5.63046e-19 $X=0.881 $Y=0.0405
c107 29 VSS 0.0127604f $X=1.377 $Y=0.136
c108 26 VSS 0.0647964f $X=1.377 $Y=0.0675
c109 18 VSS 0.0615177f $X=1.323 $Y=0.0675
c110 10 VSS 0.0579453f $X=1.269 $Y=0.0675
c111 5 VSS 0.00302777f $X=1.053 $Y=0.14
c112 2 VSS 0.0627731f $X=1.053 $Y=0.0405
r113 86 87 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=1.175
+ $Y=0.153 $X2=1.229 $Y2=0.153
r114 84 87 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.269
+ $Y=0.153 $X2=1.229 $Y2=0.153
r115 84 94 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.269 $Y=0.153 $X2=1.269
+ $Y2=0.153
r116 80 86 15.6173 $w=1.8e-08 $l=2.3e-07 $layer=M2 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=1.175 $Y2=0.153
r117 80 81 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.945 $Y=0.153 $X2=0.945
+ $Y2=0.153
r118 76 77 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r119 75 77 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r120 72 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.234 $X2=0.936 $Y2=0.234
r121 64 66 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.153 $X2=1.053 $Y2=0.14
r122 62 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.99
+ $Y=0.162 $X2=1.008 $Y2=0.162
r123 61 81 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.945 $Y2=0.162
r124 61 62 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.99 $Y2=0.162
r125 60 64 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.162 $X2=1.053 $Y2=0.153
r126 60 63 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.162 $X2=1.008 $Y2=0.162
r127 59 75 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.234
r128 58 81 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.162
r129 58 59 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.225
r130 56 57 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.119 $X2=0.945 $Y2=0.136
r131 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.101 $X2=0.945 $Y2=0.119
r132 54 55 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.081 $X2=0.945 $Y2=0.101
r133 53 81 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.162
r134 53 57 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.136
r135 52 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.081
r136 50 51 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.904
+ $Y=0.036 $X2=0.92 $Y2=0.036
r137 49 50 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.036 $X2=0.904 $Y2=0.036
r138 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r139 45 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r140 43 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r141 43 51 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.92 $Y2=0.036
r142 42 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.234
+ $X2=0.918 $Y2=0.234
r143 39 42 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.2295 $X2=0.918 $Y2=0.2295
r144 38 42 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.935 $Y=0.2295 $X2=0.918 $Y2=0.2295
r145 37 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036
+ $X2=0.864 $Y2=0.036
r146 34 37 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.864 $Y2=0.0405
r147 33 37 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0405 $X2=0.864 $Y2=0.0405
r148 29 31 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.377 $Y=0.136 $X2=1.377 $Y2=0.2025
r149 26 29 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.377 $Y=0.0675 $X2=1.377 $Y2=0.136
r150 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.323
+ $Y=0.136 $X2=1.377 $Y2=0.136
r151 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.136 $X2=1.323 $Y2=0.2025
r152 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.0675 $X2=1.323 $Y2=0.136
r153 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.269
+ $Y=0.136 $X2=1.323 $Y2=0.136
r154 13 94 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.269 $Y=0.136 $X2=1.269
+ $Y2=0.136
r155 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.136 $X2=1.269 $Y2=0.2025
r156 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.0675 $X2=1.269 $Y2=0.136
r157 5 66 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.053 $Y=0.14 $X2=1.053
+ $Y2=0.14
r158 5 7 335.312 $w=2e-08 $l=8.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.14 $X2=1.053 $Y2=0.2295
r159 2 5 372.777 $w=2e-08 $l=9.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.0405 $X2=1.053 $Y2=0.14
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%14 1 4 6 11 14 21 23 24 25 VSS
c29 26 VSS 0.00225803f $X=0.485 $Y=0.234
c30 25 VSS 0.0014167f $X=0.461 $Y=0.234
c31 24 VSS 0.0134342f $X=0.447 $Y=0.234
c32 23 VSS 0.00523898f $X=0.309 $Y=0.234
c33 21 VSS 0.00168783f $X=0.486 $Y=0.234
c34 14 VSS 0.0195485f $X=0.542 $Y=0.2025
c35 11 VSS 3.25039e-19 $X=0.557 $Y=0.2025
c36 9 VSS 4.57278e-19 $X=0.484 $Y=0.2025
c37 4 VSS 0.00250857f $X=0.272 $Y=0.2025
c38 1 VSS 3.31752e-19 $X=0.287 $Y=0.2025
r39 25 26 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.461
+ $Y=0.234 $X2=0.485 $Y2=0.234
r40 24 25 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.234 $X2=0.461 $Y2=0.234
r41 23 24 9.37037 $w=1.8e-08 $l=1.38e-07 $layer=M1 $thickness=3.6e-08 $X=0.309
+ $Y=0.234 $X2=0.447 $Y2=0.234
r42 21 26 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.485 $Y2=0.234
r43 17 23 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.309 $Y2=0.234
r44 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.542 $Y2=0.2025
r45 9 14 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.484
+ $Y=0.2025 $X2=0.542 $Y2=0.2025
r46 9 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r47 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.2025 $X2=0.484 $Y2=0.2025
r48 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r49 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.272 $Y2=0.2025
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%16 1 2 5 6 7 10 12 18 20 21 22 23 24 25 VSS
c21 25 VSS 3.8923e-20 $X=0.423 $Y=0.198
c22 24 VSS 8.46035e-21 $X=0.414 $Y=0.198
c23 23 VSS 0.00116854f $X=0.396 $Y=0.198
c24 22 VSS 0.00134991f $X=0.379 $Y=0.198
c25 21 VSS 8.46035e-21 $X=0.36 $Y=0.198
c26 20 VSS 2.61077e-19 $X=0.342 $Y=0.198
c27 18 VSS 3.31089e-19 $X=0.432 $Y=0.198
c28 12 VSS 5.44897e-19 $X=0.324 $Y=0.198
c29 10 VSS 0.00631853f $X=0.432 $Y=0.2025
c30 6 VSS 5.67296e-19 $X=0.449 $Y=0.2025
c31 5 VSS 0.00790786f $X=0.324 $Y=0.2025
c32 1 VSS 6.05629e-19 $X=0.341 $Y=0.2025
r33 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.423 $Y2=0.198
r34 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.414 $Y2=0.198
r35 22 23 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.198 $X2=0.396 $Y2=0.198
r36 21 22 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.198 $X2=0.379 $Y2=0.198
r37 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r38 18 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.423 $Y2=0.198
r39 12 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.342 $Y2=0.198
r40 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r41 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r42 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r43 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198 $X2=0.324
+ $Y2=0.198
r44 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
r45 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%QN 1 2 6 11 12 15 16 21 24 29 40 42 VSS
c16 42 VSS 0.0054983f $X=1.431 $Y=0.2
c17 41 VSS 0.00201603f $X=1.431 $Y=0.09
c18 40 VSS 0.00112176f $X=1.433 $Y=0.223
c19 29 VSS 0.01957f $X=1.422 $Y=0.234
c20 28 VSS 0.00635401f $X=1.404 $Y=0.036
c21 24 VSS 0.0097085f $X=1.296 $Y=0.036
c22 21 VSS 0.0193971f $X=1.422 $Y=0.036
c23 19 VSS 0.00670088f $X=1.402 $Y=0.2025
c24 15 VSS 0.0101265f $X=1.296 $Y=0.2025
c25 11 VSS 5.72268e-19 $X=1.313 $Y=0.2025
c26 9 VSS 3.44349e-19 $X=1.402 $Y=0.0675
c27 1 VSS 5.72268e-19 $X=1.313 $Y=0.0675
r28 41 42 7.46914 $w=1.8e-08 $l=1.1e-07 $layer=M1 $thickness=3.6e-08 $X=1.431
+ $Y=0.09 $X2=1.431 $Y2=0.2
r29 40 42 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.431
+ $Y=0.223 $X2=1.431 $Y2=0.2
r30 38 40 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.431
+ $Y=0.225 $X2=1.431 $Y2=0.223
r31 37 41 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.431
+ $Y=0.045 $X2=1.431 $Y2=0.09
r32 31 35 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.234 $X2=1.404 $Y2=0.234
r33 29 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.422 $Y=0.234 $X2=1.431 $Y2=0.225
r34 29 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.422
+ $Y=0.234 $X2=1.404 $Y2=0.234
r35 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.404 $Y=0.036 $X2=1.404
+ $Y2=0.036
r36 23 27 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.036 $X2=1.404 $Y2=0.036
r37 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.036 $X2=1.296
+ $Y2=0.036
r38 21 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.422 $Y=0.036 $X2=1.431 $Y2=0.045
r39 21 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.422
+ $Y=0.036 $X2=1.404 $Y2=0.036
r40 19 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.404 $Y=0.234 $X2=1.404
+ $Y2=0.234
r41 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.387 $Y=0.2025 $X2=1.402 $Y2=0.2025
r42 15 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.234 $X2=1.296
+ $Y2=0.234
r43 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.279 $Y=0.2025 $X2=1.296 $Y2=0.2025
r44 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.313 $Y=0.2025 $X2=1.296 $Y2=0.2025
r45 9 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.404
+ $Y=0.0675 $X2=1.404 $Y2=0.036
r46 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.387
+ $Y=0.0675 $X2=1.402 $Y2=0.0675
r47 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.296
+ $Y=0.0675 $X2=1.296 $Y2=0.036
r48 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.279
+ $Y=0.0675 $X2=1.296 $Y2=0.0675
r49 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.313
+ $Y=0.0675 $X2=1.296 $Y2=0.0675
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%19 1 6 9 VSS
c10 9 VSS 0.0140217f $X=0.704 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.719 $Y=0.2295
c12 4 VSS 2.70811e-19 $X=0.646 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.646
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.631
+ $Y=0.2295 $X2=0.646 $Y2=0.2295
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%20 1 6 9 VSS
c9 9 VSS 0.0145746f $X=0.974 $Y=0.0405
c10 6 VSS 3.14771e-19 $X=0.989 $Y=0.0405
c11 4 VSS 2.65708e-19 $X=0.916 $Y=0.0405
r12 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r13 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.916
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r14 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.901
+ $Y=0.0405 $X2=0.916 $Y2=0.0405
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%22 1 2 VSS
c2 1 VSS 0.00203573f $X=0.719 $Y=0.0405
r3 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0405 $X2=0.685 $Y2=0.0405
.ends

.subckt PM_SDFHX3_ASAP7_75T_SRAM%23 1 2 VSS
c0 1 VSS 0.00214045f $X=0.989 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.2295 $X2=0.955 $Y2=0.2295
.ends


* END of "./SDFHx3_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt SDFHx3_ASAP7_75t_SRAM  VSS VDD CLK SE D SI QN
* 
* QN	QN
* SI	SI
* D	D
* SE	SE
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_9_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_SE_M2_g noxref_15 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 noxref_21 N_6_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 noxref_17 N_D_M4_g noxref_21 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 noxref_15 N_SI_M5_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 N_11_M6_d N_4_M6_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M7 N_22_M7_d N_9_M7_g N_11_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M8 VSS N_10_M8_g N_22_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.027
M9 N_10_M9_d N_11_M9_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_13_M10_d N_9_M10_g N_10_M10_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.827 $Y=0.027
M11 N_20_M11_d N_4_M11_g N_13_M11_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.027
M12 VSS N_12_M12_g N_20_M12_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.027
M13 N_12_M13_d N_13_M13_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.027
M14 VSS N_SE_M14_g N_6_M14_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.205
+ $Y=0.027
M15 N_QN_M15_d N_13_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M16 N_QN_M16_d N_13_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.027
M17 N_QN_M17_d N_13_M17_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.367
+ $Y=0.027
M18 VDD N_CLK_M18_g N_4_M18_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M19 N_9_M19_d N_4_M19_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M20 N_16_M20_d N_SE_M20_g N_14_M20_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M21 VDD N_6_M21_g N_16_M21_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M22 N_16_M22_d N_D_M22_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M23 N_14_M23_d N_SI_M23_g N_16_M23_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M24 N_11_M24_d N_9_M24_g N_14_M24_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M25 N_19_M25_d N_4_M25_g N_11_M25_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.611 $Y=0.216
M26 VDD N_10_M26_g N_19_M26_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.216
M27 N_10_M27_d N_11_M27_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M28 N_13_M28_d N_4_M28_g N_10_M28_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.216
M29 N_23_M29_d N_9_M29_g N_13_M29_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.935 $Y=0.216
M30 VDD N_12_M30_g N_23_M30_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.216
M31 N_12_M31_d N_13_M31_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.216
M32 VDD N_SE_M32_g N_6_M32_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.205
+ $Y=0.216
M33 N_QN_M33_d N_13_M33_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
M34 N_QN_M34_d N_13_M34_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.162
M35 N_QN_M35_d N_13_M35_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.367
+ $Y=0.162
*
* 
* .include "SDFHx3_ASAP7_75t_SRAM.pex.sp.SDFHX3_ASAP7_75T_SRAM.pxi"
* BEGIN of "./SDFHx3_ASAP7_75t_SRAM.pex.sp.SDFHX3_ASAP7_75T_SRAM.pxi"
* File: SDFHx3_ASAP7_75t_SRAM.pex.sp.SDFHX3_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 13:03:48 2017
* 
x_PM_SDFHX3_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M18_g N_CLK_c_3_p CLK
+ N_CLK_c_9_p N_CLK_c_7_p N_CLK_c_19_p VSS PM_SDFHX3_ASAP7_75T_SRAM%CLK
x_PM_SDFHX3_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_21_n N_4_M19_g N_4_M6_g N_4_c_41_p
+ N_4_M25_g N_4_M11_g N_4_c_45_p N_4_M28_g N_4_M0_s N_4_c_22_n N_4_M18_s
+ N_4_c_23_n N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_54_p N_4_c_35_p
+ N_4_c_28_n N_4_c_58_p N_4_c_29_n N_4_c_56_p N_4_c_32_p N_4_c_36_p N_4_c_46_p
+ N_4_c_34_p N_4_c_64_p N_4_c_31_n N_4_c_48_p VSS PM_SDFHX3_ASAP7_75T_SRAM%4
x_PM_SDFHX3_ASAP7_75T_SRAM%SE N_SE_M2_g N_SE_c_90_p N_SE_M20_g N_SE_M14_g
+ N_SE_c_126_p N_SE_M32_g N_SE_c_95_p N_SE_c_140_p N_SE_c_138_p N_SE_c_156_p
+ N_SE_c_86_n SE N_SE_c_85_n N_SE_c_91_p N_SE_c_92_p N_SE_c_87_n N_SE_c_88_n
+ N_SE_c_136_p N_SE_c_104_p N_SE_c_108_p N_SE_c_93_p N_SE_c_137_p VSS
+ PM_SDFHX3_ASAP7_75T_SRAM%SE
x_PM_SDFHX3_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_168_n N_6_M21_g N_6_M14_s N_6_c_169_n
+ N_6_M32_s N_6_c_198_p N_6_c_205_p N_6_c_215_p N_6_c_202_p N_6_c_211_p
+ N_6_c_219_p N_6_c_171_n N_6_c_164_n N_6_c_186_p N_6_c_166_n N_6_c_174_n
+ N_6_c_177_n N_6_c_178_n N_6_c_204_p VSS PM_SDFHX3_ASAP7_75T_SRAM%6
x_PM_SDFHX3_ASAP7_75T_SRAM%D N_D_M4_g N_D_c_236_n N_D_M22_g D VSS
+ PM_SDFHX3_ASAP7_75T_SRAM%D
x_PM_SDFHX3_ASAP7_75T_SRAM%SI N_SI_M5_g N_SI_M23_g SI N_SI_c_256_n VSS
+ PM_SDFHX3_ASAP7_75T_SRAM%SI
x_PM_SDFHX3_ASAP7_75T_SRAM%9 N_9_c_278_n N_9_M24_g N_9_M7_g N_9_c_346_p N_9_M10_g
+ N_9_c_330_p N_9_c_282_n N_9_M29_g N_9_M1_d N_9_c_287_n N_9_M19_d N_9_c_288_n
+ N_9_c_289_n N_9_c_314_n N_9_c_301_n N_9_c_272_n N_9_c_374_p N_9_c_292_n
+ N_9_c_273_n N_9_c_295_n N_9_c_274_n N_9_c_298_n N_9_c_275_n N_9_c_276_n
+ N_9_c_299_n N_9_c_300_n N_9_c_277_n VSS PM_SDFHX3_ASAP7_75T_SRAM%9
x_PM_SDFHX3_ASAP7_75T_SRAM%10 N_10_M8_g N_10_M26_g N_10_M10_s N_10_M9_d
+ N_10_c_397_n N_10_M27_d N_10_c_410_n N_10_M28_s N_10_c_412_n N_10_c_400_n
+ N_10_c_401_n N_10_c_398_n N_10_c_394_n N_10_c_403_n N_10_c_399_n N_10_c_427_p
+ N_10_c_441_p N_10_c_395_n N_10_c_429_p N_10_c_396_n N_10_c_417_n N_10_c_418_n
+ N_10_c_404_n VSS PM_SDFHX3_ASAP7_75T_SRAM%10
x_PM_SDFHX3_ASAP7_75T_SRAM%11 N_11_M9_g N_11_c_443_n N_11_M27_g N_11_M6_d N_11_M7_s
+ N_11_M24_d N_11_c_444_n N_11_M25_s N_11_c_507_p N_11_c_466_n N_11_c_467_n
+ N_11_c_445_n N_11_c_453_n N_11_c_454_n N_11_c_455_n N_11_c_456_n N_11_c_457_n
+ N_11_c_490_n N_11_c_459_n N_11_c_460_n N_11_c_447_n N_11_c_510_p N_11_c_448_n
+ N_11_c_449_n N_11_c_472_n N_11_c_474_n N_11_c_477_n N_11_c_511_p N_11_c_482_n
+ N_11_c_451_n N_11_c_452_n N_11_c_486_n VSS PM_SDFHX3_ASAP7_75T_SRAM%11
x_PM_SDFHX3_ASAP7_75T_SRAM%12 N_12_M12_g N_12_c_536_p N_12_M30_g N_12_M13_d
+ N_12_c_521_n N_12_M31_d N_12_c_523_n N_12_c_515_n N_12_c_516_n N_12_c_517_n
+ N_12_c_518_n N_12_c_519_n N_12_c_527_n N_12_c_520_n N_12_c_530_n N_12_c_545_p
+ VSS PM_SDFHX3_ASAP7_75T_SRAM%12
x_PM_SDFHX3_ASAP7_75T_SRAM%13 N_13_M13_g N_13_M31_g N_13_M15_g N_13_M33_g
+ N_13_M16_g N_13_M34_g N_13_M17_g N_13_c_554_n N_13_M35_g N_13_M11_s N_13_M10_d
+ N_13_c_555_n N_13_M29_s N_13_M28_d N_13_c_579_n N_13_c_556_n N_13_c_557_n
+ N_13_c_547_n N_13_c_559_n N_13_c_560_n N_13_c_568_n N_13_c_549_n N_13_c_581_n
+ N_13_c_582_n N_13_c_627_p N_13_c_602_n N_13_c_604_n N_13_c_569_n N_13_c_550_n
+ N_13_c_561_n N_13_c_551_n N_13_c_563_n N_13_c_565_n VSS
+ PM_SDFHX3_ASAP7_75T_SRAM%13
x_PM_SDFHX3_ASAP7_75T_SRAM%14 N_14_M20_s N_14_c_629_n N_14_M23_d N_14_M24_s
+ N_14_c_628_n N_14_c_635_n N_14_c_630_n N_14_c_632_n N_14_c_636_n VSS
+ PM_SDFHX3_ASAP7_75T_SRAM%14
x_PM_SDFHX3_ASAP7_75T_SRAM%16 N_16_M21_s N_16_M20_d N_16_c_671_n N_16_M23_s
+ N_16_M22_d N_16_c_673_n N_16_c_663_n N_16_c_662_n N_16_c_665_n N_16_c_657_n
+ N_16_c_667_n N_16_c_668_n N_16_c_659_n N_16_c_661_n VSS
+ PM_SDFHX3_ASAP7_75T_SRAM%16
x_PM_SDFHX3_ASAP7_75T_SRAM%QN N_QN_M16_d N_QN_M15_d N_QN_M17_d N_QN_M34_d
+ N_QN_M33_d N_QN_c_682_n N_QN_M35_d N_QN_c_678_n N_QN_c_687_n N_QN_c_679_n QN
+ N_QN_c_692_n VSS PM_SDFHX3_ASAP7_75T_SRAM%QN
x_PM_SDFHX3_ASAP7_75T_SRAM%19 N_19_M25_d N_19_M26_s N_19_c_695_n VSS
+ PM_SDFHX3_ASAP7_75T_SRAM%19
x_PM_SDFHX3_ASAP7_75T_SRAM%20 N_20_M11_d N_20_M12_s N_20_c_704_n VSS
+ PM_SDFHX3_ASAP7_75T_SRAM%20
x_PM_SDFHX3_ASAP7_75T_SRAM%22 N_22_M8_s N_22_M7_d VSS PM_SDFHX3_ASAP7_75T_SRAM%22
x_PM_SDFHX3_ASAP7_75T_SRAM%23 N_23_M30_s N_23_M29_d VSS PM_SDFHX3_ASAP7_75T_SRAM%23
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_CLK_c_2_p N_4_c_21_n 0.00105598f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_CLK_c_3_p N_4_c_22_n 2.66516e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.054
cc_4 N_CLK_c_3_p N_4_c_23_n 0.0012473f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.144
cc_5 N_CLK_c_3_p N_4_c_24_n 3.97017e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.081
cc_6 N_CLK_c_3_p N_4_c_25_n 0.0012473f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.1125
cc_7 N_CLK_c_7_p N_4_c_26_n 0.00140648f $X=0.081 $Y=0.167 $X2=0.018 $Y2=0.2
cc_8 N_CLK_c_3_p N_4_c_27_n 4.97741e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_9_p N_4_c_28_n 0.00123168f $X=0.081 $Y=0.162 $X2=0.033 $Y2=0.153
cc_10 N_CLK_c_3_p N_4_c_29_n 5.36602e-19 $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_11 N_CLK_c_9_p N_4_c_29_n 8.66987e-19 $X=0.081 $Y=0.162 $X2=0.175 $Y2=0.153
cc_12 N_CLK_c_3_p N_4_c_31_n 0.00203815f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_13 N_CLK_c_3_p N_SE_c_85_n 2.45198e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2
cc_14 N_CLK_c_3_p N_9_c_272_n 6.32319e-19 $X=0.081 $Y=0.135 $X2=0.621 $Y2=0.135
cc_15 CLK N_9_c_273_n 3.23206e-19 $X=0.078 $Y=0.19 $X2=0.337 $Y2=0.153
cc_16 CLK N_9_c_274_n 2.57347e-19 $X=0.078 $Y=0.19 $X2=0.817 $Y2=0.153
cc_17 N_CLK_c_3_p N_9_c_275_n 0.00114506f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_18 N_CLK_c_3_p N_9_c_276_n 3.05593e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_19 N_CLK_c_19_p N_9_c_277_n 3.05593e-19 $X=0.081 $Y=0.1785 $X2=0 $Y2=0
cc_20 N_4_c_32_p N_SE_c_86_n 8.13669e-19 $X=0.337 $Y=0.153 $X2=0 $Y2=0
cc_21 N_4_c_32_p N_SE_c_87_n 0.0022834f $X=0.337 $Y=0.153 $X2=0 $Y2=0
cc_22 N_4_c_34_p N_SE_c_88_n 0.0022834f $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_23 N_4_c_35_p N_6_c_164_n 3.98881e-19 $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_24 N_4_c_36_p N_6_c_164_n 0.0176158f $X=0.479 $Y=0.153 $X2=0 $Y2=0
cc_25 N_4_c_36_p N_6_c_166_n 0.00114531f $X=0.479 $Y=0.153 $X2=0 $Y2=0
cc_26 N_4_c_36_p D 0.00102191f $X=0.479 $Y=0.153 $X2=0.081 $Y2=0.135
cc_27 N_4_c_34_p SI 0.00113575f $X=0.743 $Y=0.153 $X2=0.081 $Y2=0.135
cc_28 N_4_M6_g N_9_c_278_n 0.00365763f $X=0.621 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_29 N_4_c_41_p N_9_c_278_n 9.97803e-19 $X=0.621 $Y=0.135 $X2=0.081 $Y2=0.054
cc_30 N_4_M6_g N_9_M7_g 0.00355599f $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_4_M11_g N_9_M10_g 0.00355599f $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_32 N_4_M11_g N_9_c_282_n 0.00605856f $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.1785
cc_33 N_4_c_45_p N_9_c_282_n 0.00180656f $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.1785
cc_34 N_4_c_46_p N_9_c_282_n 5.51712e-19 $X=0.891 $Y=0.153 $X2=0.081 $Y2=0.1785
cc_35 N_4_c_34_p N_9_c_282_n 0.00168667f $X=0.743 $Y=0.153 $X2=0.081 $Y2=0.1785
cc_36 N_4_c_48_p N_9_c_282_n 0.00123876f $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.1785
cc_37 N_4_c_29_n N_9_c_287_n 2.18034e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_38 N_4_c_29_n N_9_c_288_n 2.58357e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_35_p N_9_c_289_n 0.00279251f $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_34_p N_9_c_289_n 9.87747e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_41 N_4_c_29_n N_9_c_272_n 3.93085e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_42 N_4_c_54_p N_9_c_292_n 2.66501e-19 $X=0.054 $Y=0.234 $X2=0 $Y2=0
cc_43 N_4_c_29_n N_9_c_292_n 4.19323e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_44 N_4_c_56_p N_9_c_273_n 2.46239e-19 $X=0.211 $Y=0.153 $X2=0 $Y2=0
cc_45 N_4_c_34_p N_9_c_295_n 2.46239e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_46 N_4_c_58_p N_9_c_274_n 3.80004e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_56_p N_9_c_274_n 0.0471484f $X=0.211 $Y=0.153 $X2=0 $Y2=0
cc_48 N_4_c_34_p N_9_c_298_n 2.81643e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_49 N_4_c_31_n N_9_c_299_n 0.00218805f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_50 N_4_c_56_p N_9_c_300_n 0.00116576f $X=0.211 $Y=0.153 $X2=0 $Y2=0
cc_51 N_4_M6_g N_10_M8_g 2.82885e-19 $X=0.621 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_52 N_4_c_64_p N_10_c_394_n 5.29207e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_53 N_4_c_48_p N_10_c_395_n 0.00318254f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_54 N_4_c_46_p N_10_c_396_n 0.00128311f $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_55 N_4_M11_g N_11_M9_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_56 N_4_c_45_p N_11_c_443_n 2.98891e-19 $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.135
cc_57 N_4_c_58_p N_11_c_444_n 3.24488e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_58 N_4_M6_g N_11_c_445_n 3.41974e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_59 N_4_c_58_p N_11_c_445_n 0.00102727f $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_60 N_4_c_35_p N_11_c_447_n 0.00133841f $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_61 N_4_c_34_p N_11_c_448_n 7.726e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_62 N_4_c_58_p N_11_c_449_n 8.63476e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_63 N_4_c_34_p N_11_c_449_n 5.92766e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_64 N_4_c_34_p N_11_c_451_n 3.70527e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_65 N_4_c_64_p N_11_c_452_n 3.70527e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_66 N_4_M11_g N_12_M12_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_67 N_4_M11_g N_13_c_547_n 3.18506e-19 $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_68 N_4_c_48_p N_13_c_547_n 4.09234e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_69 N_4_c_48_p N_13_c_549_n 0.00320381f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_70 N_4_c_48_p N_13_c_550_n 3.56772e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_71 N_4_c_46_p N_13_c_551_n 9.47997e-19 $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_72 N_4_c_36_p N_14_c_628_n 4.23942e-19 $X=0.479 $Y=0.153 $X2=0 $Y2=0
cc_73 N_SE_M2_g N_6_M3_g 0.00304756f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_74 N_SE_c_90_p N_6_c_168_n 0.00126421f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_75 N_SE_c_91_p N_6_c_169_n 2.11282e-19 $X=1.215 $Y=0.045 $X2=0.081 $Y2=0.135
cc_76 N_SE_c_92_p N_6_c_169_n 8.20809e-19 $X=1.215 $Y=0.045 $X2=0.081 $Y2=0.135
cc_77 N_SE_c_93_p N_6_c_171_n 3.53759e-19 $X=1.215 $Y=0.09 $X2=0 $Y2=0
cc_78 N_SE_c_88_n N_6_c_164_n 0.0680793f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_79 N_SE_c_95_p N_6_c_166_n 8.79603e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_80 N_SE_c_92_p N_6_c_174_n 0.00733801f $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_81 N_SE_c_88_n N_6_c_174_n 0.00103045f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_82 N_SE_c_93_p N_6_c_174_n 3.73635e-19 $X=1.215 $Y=0.09 $X2=0 $Y2=0
cc_83 N_SE_c_88_n N_6_c_177_n 2.46239e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_84 N_SE_c_86_n N_6_c_178_n 3.24594e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_85 N_SE_M2_g N_D_M4_g 2.13359e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_86 N_SE_c_85_n N_9_c_301_n 0.00266639f $X=0.225 $Y=0.045 $X2=0 $Y2=0
cc_87 N_SE_c_87_n N_9_c_301_n 4.45368e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_88 N_SE_c_104_p N_9_c_301_n 2.64176e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_89 N_SE_c_86_n N_9_c_274_n 4.53301e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_90 N_SE_c_87_n N_9_c_274_n 3.907e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_91 N_SE_c_104_p N_9_c_275_n 0.00292661f $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_92 N_SE_c_108_p N_9_c_276_n 0.00266639f $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_93 N_SE_c_86_n N_9_c_299_n 0.00266639f $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_94 N_SE_c_88_n N_10_c_397_n 4.38905e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_95 N_SE_c_88_n N_10_c_398_n 3.00479e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_96 N_SE_c_88_n N_10_c_399_n 7.16568e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_97 N_SE_c_88_n N_11_c_453_n 0.00113636f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_98 N_SE_c_88_n N_11_c_454_n 2.78297e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_99 N_SE_c_88_n N_11_c_455_n 5.99401e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_100 N_SE_c_88_n N_11_c_456_n 4.8504e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_101 N_SE_c_88_n N_11_c_457_n 4.65038e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_102 N_SE_c_88_n N_12_c_515_n 5.48108e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_103 N_SE_c_88_n N_12_c_516_n 0.00109158f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_104 N_SE_c_88_n N_12_c_517_n 5.50727e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_105 N_SE_c_88_n N_12_c_518_n 9.11285e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_106 N_SE_c_88_n N_12_c_519_n 4.62125e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_107 N_SE_c_88_n N_12_c_520_n 5.48546e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_108 N_SE_M14_g N_13_M15_g 0.00268443f $X=1.215 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_109 N_SE_M14_g N_13_M16_g 2.13359e-19 $X=1.215 $Y=0.0405 $X2=0.081 $Y2=0.162
cc_110 N_SE_c_126_p N_13_c_554_n 0.00115475f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_111 N_SE_c_88_n N_13_c_555_n 2.30689e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_112 N_SE_c_88_n N_13_c_556_n 9.08574e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_113 N_SE_c_88_n N_13_c_557_n 0.00124317f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_114 N_SE_c_88_n N_13_c_547_n 4.54245e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_115 N_SE_c_88_n N_13_c_559_n 4.39544e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_116 N_SE_c_88_n N_13_c_560_n 5.37888e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_117 N_SE_c_92_p N_13_c_561_n 3.26078e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_118 N_SE_c_88_n N_13_c_551_n 9.36021e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_119 N_SE_c_91_p N_13_c_563_n 9.36021e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_120 N_SE_c_136_p N_13_c_563_n 0.00114818f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_121 N_SE_c_137_p N_13_c_565_n 0.00409386f $X=1.215 $Y=0.113 $X2=0 $Y2=0
cc_122 N_SE_c_138_p N_14_c_629_n 2.31793e-19 $X=0.261 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_123 N_SE_M2_g N_14_c_630_n 3.83731e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_124 N_SE_c_140_p N_14_c_630_n 6.51345e-19 $X=0.258 $Y=0.135 $X2=0 $Y2=0
cc_125 VSS N_SE_c_85_n 2.40719e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.135
cc_126 VSS N_SE_c_87_n 5.30841e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.135
cc_127 VSS N_SE_c_104_p 9.86432e-19 $X=0.225 $Y=0.081 $X2=0.081 $Y2=0.135
cc_128 VSS N_SE_c_95_p 0.00129447f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_129 VSS N_SE_c_87_n 7.061e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_130 VSS N_SE_c_104_p 7.68051e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_131 VSS N_SE_c_85_n 8.44602e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.19
cc_132 VSS N_SE_c_87_n 5.36527e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.19
cc_133 VSS N_SE_c_88_n 0.00141783f $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.144
cc_134 VSS N_SE_c_88_n 2.35788e-19 $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.162
cc_135 VSS N_SE_c_87_n 6.93145e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.1785
cc_136 VSS N_SE_c_88_n 9.13621e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_137 VSS N_SE_c_88_n 4.6862e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_138 VSS N_SE_c_88_n 5.41611e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_139 VSS N_SE_c_88_n 8.51044e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_140 VSS N_SE_c_156_p 0.00129447f $X=0.279 $Y=0.135 $X2=0 $Y2=0
cc_141 VSS N_SE_c_87_n 3.48715e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_142 VSS N_SE_c_108_p 9.77595e-19 $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_143 VSS N_SE_c_88_n 2.40178e-19 $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.135
cc_144 VSS N_SE_c_88_n 6.42719e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_145 VSS N_SE_c_88_n 0.00110738f $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.162
cc_146 N_SE_c_92_p N_QN_c_678_n 8.3796e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_147 N_SE_c_88_n N_20_c_704_n 4.98441e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_148 N_6_M3_g N_D_M4_g 0.00304756f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_149 N_6_c_168_n N_D_c_236_n 9.71463e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_150 N_6_c_164_n D 3.33994e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_151 N_6_c_166_n D 0.00195518f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_152 N_6_c_178_n D 9.77589e-19 $X=0.351 $Y=0.126 $X2=0 $Y2=0
cc_153 N_6_M3_g N_SI_M5_g 2.48122e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_154 N_6_c_164_n SI 3.40688e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_155 N_6_c_186_p N_9_c_282_n 3.37164e-19 $X=0.936 $Y=0.081 $X2=0.891 $Y2=0.135
cc_156 N_6_c_164_n N_9_c_274_n 0.0011956f $X=0.9 $Y=0.081 $X2=0.817 $Y2=0.153
cc_157 N_6_c_164_n N_10_c_400_n 5.04077e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_158 N_6_c_164_n N_10_c_401_n 2.53924e-19 $X=0.9 $Y=0.081 $X2=0.056 $Y2=0.054
cc_159 N_6_c_164_n N_10_c_398_n 8.29294e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_160 N_6_c_164_n N_10_c_403_n 5.75824e-19 $X=0.9 $Y=0.081 $X2=0.018 $Y2=0.144
cc_161 N_6_c_164_n N_10_c_404_n 7.91051e-19 $X=0.9 $Y=0.081 $X2=0.047 $Y2=0.234
cc_162 N_6_c_164_n N_11_c_454_n 4.20387e-19 $X=0.9 $Y=0.081 $X2=0.018 $Y2=0.081
cc_163 N_6_c_164_n N_11_c_459_n 4.92006e-19 $X=0.9 $Y=0.081 $X2=0.054 $Y2=0.036
cc_164 N_6_c_164_n N_11_c_460_n 7.19039e-19 $X=0.9 $Y=0.081 $X2=0.054 $Y2=0.036
cc_165 N_6_c_169_n N_12_c_521_n 0.00124414f $X=1.19 $Y=0.0405 $X2=0.621
+ $Y2=0.135
cc_166 N_6_c_171_n N_12_c_521_n 2.40393e-19 $X=1.161 $Y=0.081 $X2=0.621
+ $Y2=0.135
cc_167 N_6_c_198_p N_12_c_523_n 5.25714e-19 $X=1.19 $Y=0.2295 $X2=0.891
+ $Y2=0.0405
cc_168 N_6_c_171_n N_12_c_515_n 9.95523e-19 $X=1.161 $Y=0.081 $X2=0.891
+ $Y2=0.135
cc_169 N_6_c_169_n N_12_c_516_n 3.43147e-19 $X=1.19 $Y=0.0405 $X2=0.071
+ $Y2=0.054
cc_170 N_6_c_174_n N_12_c_516_n 0.00251979f $X=1.161 $Y=0.049 $X2=0.071
+ $Y2=0.054
cc_171 N_6_c_202_p N_12_c_527_n 0.00251979f $X=1.17 $Y=0.234 $X2=0.018 $Y2=0.045
cc_172 N_6_c_171_n N_12_c_520_n 0.0012739f $X=1.161 $Y=0.081 $X2=0.018 $Y2=0.144
cc_173 N_6_c_204_p N_12_c_520_n 0.00251979f $X=1.161 $Y=0.2125 $X2=0.018
+ $Y2=0.144
cc_174 N_6_c_205_p N_12_c_530_n 0.00251979f $X=1.161 $Y=0.225 $X2=0.018
+ $Y2=0.081
cc_175 N_6_c_186_p N_13_c_557_n 6.23859e-19 $X=0.936 $Y=0.081 $X2=0.0505
+ $Y2=0.036
cc_176 N_6_c_171_n N_13_c_560_n 3.66836e-19 $X=1.161 $Y=0.081 $X2=0.047
+ $Y2=0.234
cc_177 N_6_c_171_n N_13_c_568_n 5.24665e-19 $X=1.161 $Y=0.081 $X2=0.0505
+ $Y2=0.234
cc_178 N_6_c_186_p N_13_c_569_n 3.12147e-19 $X=0.936 $Y=0.081 $X2=0.891
+ $Y2=0.153
cc_179 N_6_c_169_n N_13_c_551_n 2.50315e-19 $X=1.19 $Y=0.0405 $X2=0 $Y2=0
cc_180 N_6_c_211_p N_13_c_551_n 3.14624e-19 $X=1.179 $Y=0.234 $X2=0 $Y2=0
cc_181 N_6_c_171_n N_13_c_551_n 0.00815696f $X=1.161 $Y=0.081 $X2=0 $Y2=0
cc_182 N_6_c_174_n N_13_c_551_n 0.00110082f $X=1.161 $Y=0.049 $X2=0 $Y2=0
cc_183 N_6_c_198_p N_13_c_563_n 2.19627e-19 $X=1.19 $Y=0.2295 $X2=0 $Y2=0
cc_184 N_6_c_215_p N_13_c_563_n 3.14624e-19 $X=1.188 $Y=0.234 $X2=0 $Y2=0
cc_185 N_6_M3_g N_14_c_632_n 2.37298e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_186 VSS N_6_c_164_n 3.90811e-19 $X=0.9 $Y=0.081 $X2=0.621 $Y2=0.135
cc_187 VSS N_6_c_177_n 7.35661e-19 $X=0.351 $Y=0.099 $X2=0.621 $Y2=0.135
cc_188 VSS N_6_c_219_p 6.42252e-19 $X=0.351 $Y=0.081 $X2=0.621 $Y2=0.2295
cc_189 VSS N_6_c_219_p 0.00369658f $X=0.351 $Y=0.081 $X2=0.891 $Y2=0.135
cc_190 N_6_M3_g N_16_c_657_n 2.50526e-19 $X=0.351 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_191 N_6_c_166_n N_16_c_657_n 0.00110314f $X=0.351 $Y=0.135 $X2=0.891
+ $Y2=0.135
cc_192 VSS N_6_c_177_n 2.30452e-19 $X=0.351 $Y=0.099 $X2=0.135 $Y2=0.135
cc_193 VSS N_6_c_164_n 7.92007e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_194 VSS N_6_c_219_p 8.14481e-19 $X=0.351 $Y=0.081 $X2=0.891 $Y2=0.0405
cc_195 VSS N_6_c_164_n 2.67459e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_196 VSS N_6_c_164_n 3.16736e-19 $X=0.9 $Y=0.081 $X2=0.891 $Y2=0.135
cc_197 VSS N_6_c_164_n 2.43408e-19 $X=0.9 $Y=0.081 $X2=0.891 $Y2=0.135
cc_198 VSS N_6_c_164_n 5.19239e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_199 N_6_c_215_p N_QN_c_679_n 2.75088e-19 $X=1.188 $Y=0.234 $X2=0 $Y2=0
cc_200 N_6_c_186_p N_20_c_704_n 5.02041e-19 $X=0.936 $Y=0.081 $X2=0.621
+ $Y2=0.0675
cc_201 VSS N_6_c_219_p 2.73492e-19 $X=0.351 $Y=0.081 $X2=0.135 $Y2=0.054
cc_202 N_D_M4_g N_SI_M5_g 0.00348334f $X=0.405 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_203 D SI 7.00288e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_204 N_D_c_236_n N_SI_c_256_n 0.00109838f $X=0.405 $Y=0.135 $X2=0.621
+ $Y2=0.2295
cc_205 N_D_M4_g N_14_c_632_n 2.37298e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_206 VSS N_D_M4_g 3.08888e-19 $X=0.405 $Y=0.0675 $X2=0.891 $Y2=0.2295
cc_207 VSS D 5.77345e-19 $X=0.405 $Y=0.134 $X2=0.891 $Y2=0.2295
cc_208 N_D_M4_g N_16_c_659_n 2.43567e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_209 D N_16_c_659_n 0.00108212f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_210 D N_16_c_661_n 3.4434e-19 $X=0.405 $Y=0.134 $X2=0.071 $Y2=0.054
cc_211 VSS D 8.86227e-19 $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.135
cc_212 VSS D 0.00161923f $X=0.405 $Y=0.134 $X2=0.891 $Y2=0.0405
cc_213 N_SI_M5_g N_9_c_278_n 2.94371e-19 $X=0.459 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_214 N_SI_c_256_n N_9_c_278_n 5.18435e-19 $X=0.475 $Y=0.135 $X2=0.135
+ $Y2=0.054
cc_215 SI N_9_c_289_n 0.00114959f $X=0.473 $Y=0.135 $X2=0 $Y2=0
cc_216 SI N_9_c_314_n 0.00114959f $X=0.473 $Y=0.135 $X2=0.054 $Y2=0.234
cc_217 SI N_9_c_295_n 0.00239259f $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.153
cc_218 SI N_9_c_274_n 0.00167124f $X=0.473 $Y=0.135 $X2=0.817 $Y2=0.153
cc_219 SI N_14_c_628_n 0.00560919f $X=0.473 $Y=0.135 $X2=0.621 $Y2=0.2295
cc_220 SI N_14_c_635_n 0.00167456f $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.135
cc_221 N_SI_M5_g N_14_c_636_n 2.70361e-19 $X=0.459 $Y=0.0675 $X2=0.071 $Y2=0.054
cc_222 SI N_16_c_662_n 6.69571e-19 $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.0405
cc_223 VSS N_SI_M5_g 3.10987e-19 $X=0.459 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_224 VSS N_SI_c_256_n 2.08525e-19 $X=0.475 $Y=0.135 $X2=0.891 $Y2=0.135
cc_225 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.135
cc_226 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.2295
cc_227 VSS SI 0.00110314f $X=0.473 $Y=0.135 $X2=0.891 $Y2=0.2295
cc_228 N_9_M7_g N_10_M8_g 0.00341068f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_229 N_9_M10_g N_10_M8_g 2.13359e-19 $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_230 N_9_c_282_n N_10_M8_g 0.00205997f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_231 N_9_c_298_n N_10_M8_g 3.19768e-19 $X=0.729 $Y=0.18 $X2=0.081 $Y2=0.054
cc_232 N_9_c_282_n N_10_c_397_n 5.52012e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_233 N_9_c_282_n N_10_c_410_n 2.12581e-19 $X=0.945 $Y=0.178 $X2=0.081
+ $Y2=0.144
cc_234 N_9_c_282_n N_10_M28_s 2.50995e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.167
cc_235 N_9_M10_g N_10_c_412_n 0.00200065f $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_236 N_9_c_282_n N_10_c_412_n 0.00322783f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_237 N_9_c_282_n N_10_c_394_n 3.41745e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_238 N_9_M10_g N_10_c_395_n 2.74825e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_239 N_9_M10_g N_10_c_396_n 2.10136e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_240 N_9_c_298_n N_10_c_417_n 6.73839e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_241 N_9_c_330_p N_10_c_418_n 0.00195059f $X=0.837 $Y=0.178 $X2=0 $Y2=0
cc_242 N_9_c_282_n N_10_c_418_n 0.00191847f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_243 N_9_M10_g N_10_c_404_n 3.61755e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_244 N_9_M7_g N_11_M9_g 2.13359e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_245 N_9_M10_g N_11_M9_g 0.00341068f $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_246 N_9_c_282_n N_11_M9_g 0.00302156f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_247 N_9_c_289_n N_11_c_444_n 7.70794e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_248 N_9_c_295_n N_11_c_444_n 0.001307f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_249 N_9_c_295_n N_11_c_466_n 0.00138499f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_250 N_9_c_274_n N_11_c_467_n 0.00160025f $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_251 N_9_M7_g N_11_c_453_n 4.38308e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_252 N_9_M7_g N_11_c_459_n 2.0845e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_253 N_9_M7_g N_11_c_460_n 2.27141e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_254 N_9_c_282_n N_11_c_449_n 0.0361494f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_255 N_9_c_282_n N_11_c_472_n 2.38252e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_256 N_9_c_298_n N_11_c_472_n 0.00386452f $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_257 N_9_c_346_p N_11_c_474_n 7.00743e-19 $X=0.675 $Y=0.178 $X2=0 $Y2=0
cc_258 N_9_c_282_n N_11_c_474_n 7.89771e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_259 N_9_c_274_n N_11_c_474_n 4.88732e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_260 N_9_M7_g N_11_c_477_n 2.5554e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_261 N_9_c_282_n N_11_c_477_n 3.47488e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_262 N_9_c_295_n N_11_c_477_n 2.13133e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_263 N_9_c_274_n N_11_c_477_n 4.32971e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_264 N_9_c_298_n N_11_c_477_n 2.60223e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_265 N_9_c_282_n N_11_c_482_n 4.26771e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_266 N_9_c_282_n N_11_c_451_n 4.41163e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_267 N_9_c_282_n N_11_c_452_n 3.33141e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_268 N_9_c_298_n N_11_c_452_n 9.1388e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_269 N_9_M7_g N_11_c_486_n 2.11651e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_270 N_9_c_282_n N_12_M12_g 0.00341068f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_271 N_9_c_282_n N_13_M13_g 2.13359e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_272 N_9_c_282_n N_13_c_555_n 8.27183e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_273 N_9_c_282_n N_13_M29_s 3.37661e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_274 N_9_c_282_n N_13_c_579_n 0.00145657f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_275 N_9_c_282_n N_13_c_568_n 3.13444e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_276 N_9_c_282_n N_13_c_581_n 2.6418e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_277 N_9_c_282_n N_13_c_582_n 0.00294656f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_278 N_9_c_282_n N_13_c_569_n 3.75802e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_279 N_9_c_282_n N_13_c_550_n 5.46321e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_280 N_9_c_288_n N_14_c_629_n 9.65806e-19 $X=0.16 $Y=0.216 $X2=0.081 $Y2=0.135
cc_281 N_9_c_274_n N_14_c_629_n 4.65646e-19 $X=0.729 $Y=0.189 $X2=0.081
+ $Y2=0.135
cc_282 N_9_c_300_n N_14_c_629_n 0.00109797f $X=0.189 $Y=0.164 $X2=0.081
+ $Y2=0.135
cc_283 N_9_c_289_n N_14_c_628_n 9.68946e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_284 N_9_c_274_n N_14_c_628_n 6.49405e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_285 N_9_c_374_p N_14_c_630_n 7.61293e-19 $X=0.189 $Y=0.234 $X2=0 $Y2=0
cc_286 N_9_c_274_n N_14_c_630_n 7.84624e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_287 N_9_c_274_n N_14_c_636_n 6.22262e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_288 VSS N_9_c_287_n 9.30745e-19 $X=0.16 $Y=0.054 $X2=0.081 $Y2=0.135
cc_289 N_9_c_274_n N_16_c_663_n 2.13751e-19 $X=0.729 $Y=0.189 $X2=0.081
+ $Y2=0.135
cc_290 N_9_c_274_n N_16_c_662_n 7.1298e-19 $X=0.729 $Y=0.189 $X2=0.081 $Y2=0.162
cc_291 N_9_c_274_n N_16_c_665_n 6.46208e-19 $X=0.729 $Y=0.189 $X2=0.081
+ $Y2=0.1785
cc_292 N_9_c_274_n N_16_c_657_n 4.50553e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_293 N_9_c_274_n N_16_c_667_n 4.86474e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_294 N_9_c_274_n N_16_c_668_n 4.60071e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_295 N_9_c_274_n N_16_c_659_n 4.38038e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_296 N_9_c_274_n N_16_c_661_n 2.31538e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_297 VSS N_9_c_278_n 3.33061e-19 $X=0.567 $Y=0.1355 $X2=0 $Y2=0
cc_298 VSS N_9_c_289_n 0.00110314f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_299 N_9_c_282_n N_19_M26_s 2.33161e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.216
cc_300 N_9_M7_g N_19_c_695_n 0.00248549f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_301 N_9_c_282_n N_19_c_695_n 0.00208457f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_302 N_9_c_274_n N_19_c_695_n 7.88525e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_303 N_9_c_282_n N_20_c_704_n 0.00250239f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_304 N_10_M8_g N_11_M9_g 0.00268443f $X=0.729 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_305 N_10_c_398_n N_11_M9_g 3.7702e-19 $X=0.792 $Y=0.09 $X2=0.135 $Y2=0.054
cc_306 N_10_c_399_n N_11_c_457_n 2.46574e-19 $X=0.81 $Y=0.054 $X2=0.027
+ $Y2=0.036
cc_307 N_10_c_400_n N_11_c_490_n 0.00360624f $X=0.747 $Y=0.09 $X2=0.054
+ $Y2=0.036
cc_308 N_10_c_401_n N_11_c_459_n 3.99428e-19 $X=0.747 $Y=0.09 $X2=0.054
+ $Y2=0.036
cc_309 N_10_c_396_n N_11_c_448_n 2.22221e-19 $X=0.837 $Y=0.165 $X2=0.054
+ $Y2=0.234
cc_310 N_10_c_427_p N_11_c_477_n 2.22221e-19 $X=0.837 $Y=0.225 $X2=0.0505
+ $Y2=0.234
cc_311 N_10_c_398_n N_11_c_482_n 0.00205899f $X=0.792 $Y=0.09 $X2=0.621
+ $Y2=0.135
cc_312 N_10_c_429_p N_11_c_482_n 7.38434e-19 $X=0.837 $Y=0.14 $X2=0.621
+ $Y2=0.135
cc_313 N_10_M8_g N_11_c_452_n 3.21351e-19 $X=0.729 $Y=0.0405 $X2=0.033 $Y2=0.153
cc_314 N_10_c_400_n N_11_c_452_n 0.00205899f $X=0.747 $Y=0.09 $X2=0.033
+ $Y2=0.153
cc_315 N_10_c_397_n N_13_c_555_n 0.00379158f $X=0.81 $Y=0.0405 $X2=0.018
+ $Y2=0.081
cc_316 N_10_c_399_n N_13_c_555_n 2.84891e-19 $X=0.81 $Y=0.054 $X2=0.018
+ $Y2=0.081
cc_317 N_10_c_404_n N_13_c_555_n 2.08929e-19 $X=0.837 $Y=0.09 $X2=0.018
+ $Y2=0.081
cc_318 N_10_c_412_n N_13_c_579_n 0.00222825f $X=0.866 $Y=0.2295 $X2=0.018
+ $Y2=0.2125
cc_319 N_10_c_397_n N_13_c_557_n 3.41768e-19 $X=0.81 $Y=0.0405 $X2=0.0505
+ $Y2=0.036
cc_320 N_10_c_404_n N_13_c_568_n 4.2911e-19 $X=0.837 $Y=0.09 $X2=0.0505
+ $Y2=0.234
cc_321 N_10_c_418_n N_13_c_582_n 4.2911e-19 $X=0.837 $Y=0.207 $X2=0.621
+ $Y2=0.135
cc_322 N_10_c_412_n N_13_c_569_n 3.64454e-19 $X=0.866 $Y=0.2295 $X2=0.891
+ $Y2=0.153
cc_323 N_10_c_394_n N_13_c_569_n 4.86017e-19 $X=0.828 $Y=0.234 $X2=0.891
+ $Y2=0.153
cc_324 N_10_c_441_p N_13_c_550_n 4.2911e-19 $X=0.837 $Y=0.101 $X2=0 $Y2=0
cc_325 N_11_c_444_n N_14_c_628_n 0.00424458f $X=0.594 $Y=0.2025 $X2=0.621
+ $Y2=0.2295
cc_326 N_11_c_466_n N_14_c_628_n 4.3429e-19 $X=0.595 $Y=0.234 $X2=0.621
+ $Y2=0.2295
cc_327 N_11_c_466_n N_14_c_635_n 2.8677e-19 $X=0.595 $Y=0.234 $X2=0.891
+ $Y2=0.135
cc_328 VSS N_11_c_444_n 0.0016174f $X=0.594 $Y=0.2025 $X2=0.621 $Y2=0.0675
cc_329 VSS N_11_c_454_n 0.00414127f $X=0.648 $Y=0.036 $X2=0.621 $Y2=0.0675
cc_330 VSS N_11_c_455_n 3.30384e-19 $X=0.649 $Y=0.036 $X2=0.621 $Y2=0.0675
cc_331 VSS N_11_c_454_n 2.79363e-19 $X=0.648 $Y=0.036 $X2=0 $Y2=0
cc_332 VSS N_11_c_459_n 2.70508e-19 $X=0.693 $Y=0.081 $X2=0 $Y2=0
cc_333 N_11_c_444_n N_19_c_695_n 0.00167238f $X=0.594 $Y=0.2025 $X2=0.621
+ $Y2=0.0675
cc_334 N_11_c_507_p N_19_c_695_n 0.00315491f $X=0.684 $Y=0.234 $X2=0.621
+ $Y2=0.0675
cc_335 N_11_c_445_n N_19_c_695_n 0.00111131f $X=0.649 $Y=0.234 $X2=0.621
+ $Y2=0.0675
cc_336 N_11_c_454_n N_19_c_695_n 5.67227e-19 $X=0.648 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_337 N_11_c_510_p N_19_c_695_n 4.0515e-19 $X=0.693 $Y=0.225 $X2=0.621
+ $Y2=0.0675
cc_338 N_11_c_511_p N_19_c_695_n 0.0409693f $X=0.693 $Y=0.216 $X2=0.621
+ $Y2=0.0675
cc_339 N_11_c_453_n N_22_M8_s 2.44135e-19 $X=0.684 $Y=0.036 $X2=0.135 $Y2=0.054
cc_340 N_11_c_457_n N_22_M8_s 3.62465e-19 $X=0.693 $Y=0.062 $X2=0.135 $Y2=0.054
cc_341 N_12_M12_g N_13_M13_g 0.00268443f $X=0.999 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_342 N_12_c_519_n N_13_M13_g 3.55314e-19 $X=1.062 $Y=0.036 $X2=0.135 $Y2=0.054
cc_343 N_12_c_517_n N_13_c_556_n 0.00136796f $X=1.008 $Y=0.036 $X2=0.027
+ $Y2=0.036
cc_344 N_12_c_515_n N_13_c_560_n 0.00136796f $X=0.999 $Y=0.105 $X2=0.047
+ $Y2=0.234
cc_345 N_12_c_536_p N_13_c_568_n 3.34766e-19 $X=0.999 $Y=0.1055 $X2=0.0505
+ $Y2=0.234
cc_346 N_12_c_515_n N_13_c_568_n 0.00136796f $X=0.999 $Y=0.105 $X2=0.0505
+ $Y2=0.234
cc_347 N_12_c_527_n N_13_c_582_n 5.28703e-19 $X=1.107 $Y=0.225 $X2=0.621
+ $Y2=0.135
cc_348 N_12_M12_g N_13_c_602_n 6.35734e-19 $X=0.999 $Y=0.0405 $X2=0.033
+ $Y2=0.153
cc_349 N_12_c_515_n N_13_c_602_n 7.99759e-19 $X=0.999 $Y=0.105 $X2=0.033
+ $Y2=0.153
cc_350 N_12_c_519_n N_13_c_604_n 2.75024e-19 $X=1.062 $Y=0.036 $X2=0.135
+ $Y2=0.153
cc_351 N_12_c_530_n N_13_c_604_n 0.00266666f $X=1.107 $Y=0.171 $X2=0.135
+ $Y2=0.153
cc_352 N_12_c_523_n N_13_c_551_n 2.19627e-19 $X=1.078 $Y=0.2295 $X2=0 $Y2=0
cc_353 N_12_c_530_n N_13_c_551_n 0.00106087f $X=1.107 $Y=0.171 $X2=0 $Y2=0
cc_354 N_12_c_545_p N_13_c_551_n 5.80975e-19 $X=1.098 $Y=0.234 $X2=0 $Y2=0
cc_355 N_12_c_517_n N_20_c_704_n 5.06067e-19 $X=1.008 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_356 N_13_c_554_n N_QN_M16_d 3.7444e-19 $X=1.377 $Y=0.136 $X2=0.135 $Y2=0.054
cc_357 N_13_c_554_n N_QN_M34_d 3.85232e-19 $X=1.377 $Y=0.136 $X2=0 $Y2=0
cc_358 N_13_c_554_n N_QN_c_682_n 8.43851e-19 $X=1.377 $Y=0.136 $X2=0.621
+ $Y2=0.2295
cc_359 N_13_c_565_n N_QN_c_682_n 0.00133574f $X=1.269 $Y=0.136 $X2=0.621
+ $Y2=0.2295
cc_360 N_13_M16_g N_QN_c_678_n 4.61823e-19 $X=1.323 $Y=0.0675 $X2=0.891
+ $Y2=0.135
cc_361 N_13_M17_g N_QN_c_678_n 4.61823e-19 $X=1.377 $Y=0.0675 $X2=0.891
+ $Y2=0.135
cc_362 N_13_c_554_n N_QN_c_678_n 0.00133259f $X=1.377 $Y=0.136 $X2=0.891
+ $Y2=0.135
cc_363 N_13_c_554_n N_QN_c_687_n 7.60428e-19 $X=1.377 $Y=0.136 $X2=0 $Y2=0
cc_364 N_13_c_565_n N_QN_c_687_n 6.32721e-19 $X=1.269 $Y=0.136 $X2=0 $Y2=0
cc_365 N_13_M16_g N_QN_c_679_n 4.56718e-19 $X=1.323 $Y=0.0675 $X2=0 $Y2=0
cc_366 N_13_M17_g N_QN_c_679_n 4.56718e-19 $X=1.377 $Y=0.0675 $X2=0 $Y2=0
cc_367 N_13_c_554_n N_QN_c_679_n 0.00135857f $X=1.377 $Y=0.136 $X2=0 $Y2=0
cc_368 N_13_c_554_n N_QN_c_692_n 3.72803e-19 $X=1.377 $Y=0.136 $X2=0.018
+ $Y2=0.2125
cc_369 N_13_c_565_n N_QN_c_692_n 5.78697e-19 $X=1.269 $Y=0.136 $X2=0.018
+ $Y2=0.2125
cc_370 N_13_c_555_n N_20_c_704_n 0.00210698f $X=0.864 $Y=0.0405 $X2=0.621
+ $Y2=0.0675
cc_371 N_13_c_556_n N_20_c_704_n 0.00203632f $X=0.936 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_372 N_13_c_559_n N_20_c_704_n 0.00129774f $X=0.92 $Y=0.036 $X2=0.621
+ $Y2=0.0675
cc_373 N_13_c_560_n N_20_c_704_n 0.00104094f $X=0.945 $Y=0.081 $X2=0.621
+ $Y2=0.0675
cc_374 N_13_c_627_p N_20_c_704_n 2.5109e-19 $X=0.99 $Y=0.162 $X2=0.621
+ $Y2=0.0675
cc_375 VSS N_14_c_629_n 0.00156967f $X=0.272 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_376 VSS N_14_c_628_n 0.00145555f $X=0.542 $Y=0.2025 $X2=0.891 $Y2=0.0405
cc_377 N_14_c_629_n N_16_c_671_n 0.003872f $X=0.272 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_378 N_14_c_632_n N_16_c_671_n 0.00248801f $X=0.447 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_379 N_14_c_628_n N_16_c_673_n 0.00434154f $X=0.542 $Y=0.2025 $X2=0.621
+ $Y2=0.0675
cc_380 N_14_c_632_n N_16_c_673_n 0.0025506f $X=0.447 $Y=0.234 $X2=0.621
+ $Y2=0.0675
cc_381 N_14_c_629_n N_16_c_663_n 3.19827e-19 $X=0.272 $Y=0.2025 $X2=0.621
+ $Y2=0.135
cc_382 N_14_c_632_n N_16_c_663_n 0.0113176f $X=0.447 $Y=0.234 $X2=0.621
+ $Y2=0.135
cc_383 VSS N_14_c_628_n 4.53012e-19 $X=0.542 $Y=0.2025 $X2=0 $Y2=0
cc_384 VSS N_16_c_673_n 0.00141703f $X=0.432 $Y=0.2025 $X2=0.135 $Y2=0.135

* END of "./SDFHx3_ASAP7_75t_SRAM.pex.sp.SDFHX3_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: SDFHx4_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 13:04:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "SDFHx4_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./SDFHx4_ASAP7_75t_SRAM.pex.sp.pex"
* File: SDFHx4_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 13:04:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_SDFHX4_ASAP7_75T_SRAM%CLK 2 5 7 11 VSS
c13 11 VSS 0.00547289f $X=0.081 $Y=0.1345
c14 5 VSS 0.00201135f $X=0.081 $Y=0.135
c15 2 VSS 0.0654663f $X=0.081 $Y=0.0675
r16 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%4 2 5 7 10 16 19 22 25 28 31 33 38 41 44 46 49 53
+ 54 62 69 77 78 86 88 89 93 99 100 104 109 114 VSS
c129 149 VSS 1.06551e-19 $X=0.03 $Y=0.153
c130 148 VSS 6.89947e-19 $X=0.027 $Y=0.153
c131 114 VSS 6.93139e-19 $X=1.161 $Y=0.135
c132 109 VSS 0.00122127f $X=1.053 $Y=0.135
c133 104 VSS 0.00139543f $X=0.837 $Y=0.135
c134 100 VSS 0.00122905f $X=0.693 $Y=0.135
c135 99 VSS 0.00304316f $X=0.693 $Y=0.135
c136 93 VSS 0.00227426f $X=0.135 $Y=0.135
c137 89 VSS 6.85269e-19 $X=1.141 $Y=0.153
c138 88 VSS 0.0136835f $X=1.121 $Y=0.153
c139 86 VSS 0.00121093f $X=1.161 $Y=0.153
c140 78 VSS 0.00841321f $X=0.434 $Y=0.153
c141 77 VSS 0.00707542f $X=0.175 $Y=0.153
c142 69 VSS 6.34103e-19 $X=0.033 $Y=0.153
c143 65 VSS 2.97869e-19 $X=0.0505 $Y=0.234
c144 64 VSS 0.00179897f $X=0.047 $Y=0.234
c145 62 VSS 0.00251086f $X=0.054 $Y=0.234
c146 60 VSS 0.00305101f $X=0.027 $Y=0.234
c147 56 VSS 2.97869e-19 $X=0.0505 $Y=0.036
c148 55 VSS 0.00199279f $X=0.047 $Y=0.036
c149 54 VSS 0.00633992f $X=0.054 $Y=0.036
c150 53 VSS 0.00448137f $X=0.054 $Y=0.036
c151 51 VSS 0.00306551f $X=0.027 $Y=0.036
c152 50 VSS 5.16336e-19 $X=0.018 $Y=0.2125
c153 49 VSS 0.00162011f $X=0.018 $Y=0.2
c154 48 VSS 4.96914e-19 $X=0.018 $Y=0.225
c155 46 VSS 0.00171312f $X=0.018 $Y=0.1035
c156 45 VSS 7.23544e-19 $X=0.018 $Y=0.063
c157 44 VSS 0.00176309f $X=0.018 $Y=0.144
c158 41 VSS 0.00628074f $X=0.056 $Y=0.2025
c159 38 VSS 3.02808e-19 $X=0.071 $Y=0.2025
c160 33 VSS 2.55988e-19 $X=0.071 $Y=0.0675
c161 31 VSS 8.78713e-19 $X=1.161 $Y=0.135
c162 28 VSS 0.0586114f $X=1.161 $Y=0.0675
c163 22 VSS 0.0642113f $X=1.053 $Y=0.135
c164 16 VSS 0.0600934f $X=0.837 $Y=0.135
c165 10 VSS 0.0644358f $X=0.675 $Y=0.0675
c166 5 VSS 0.00184301f $X=0.135 $Y=0.135
c167 2 VSS 0.0641982f $X=0.135 $Y=0.0675
r168 148 149 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r169 145 148 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r170 99 100 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.693 $Y=0.135
+ $X2=0.693 $Y2=0.135
r171 88 89 1.35802 $w=1.8e-08 $l=2e-08 $layer=M2 $thickness=3.6e-08 $X=1.121
+ $Y=0.153 $X2=1.141 $Y2=0.153
r172 86 89 1.35802 $w=1.8e-08 $l=2e-08 $layer=M2 $thickness=3.6e-08 $X=1.161
+ $Y=0.153 $X2=1.141 $Y2=0.153
r173 86 114 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.161 $Y=0.153 $X2=1.161
+ $Y2=0.153
r174 83 88 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=1.053
+ $Y=0.153 $X2=1.121 $Y2=0.153
r175 83 109 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.053 $Y=0.153 $X2=1.053
+ $Y2=0.153
r176 80 83 14.6667 $w=1.8e-08 $l=2.16e-07 $layer=M2 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=1.053 $Y2=0.153
r177 80 104 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.837 $Y=0.153 $X2=0.837
+ $Y2=0.153
r178 77 78 17.5864 $w=1.8e-08 $l=2.59e-07 $layer=M2 $thickness=3.6e-08 $X=0.175
+ $Y=0.153 $X2=0.434 $Y2=0.153
r179 75 80 9.77778 $w=1.8e-08 $l=1.44e-07 $layer=M2 $thickness=3.6e-08 $X=0.693
+ $Y=0.153 $X2=0.837 $Y2=0.153
r180 75 78 17.5864 $w=1.8e-08 $l=2.59e-07 $layer=M2 $thickness=3.6e-08 $X=0.693
+ $Y=0.153 $X2=0.434 $Y2=0.153
r181 75 100 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.693 $Y=0.153 $X2=0.693
+ $Y2=0.153
r182 72 77 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.153 $X2=0.175 $Y2=0.153
r183 72 93 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.135 $Y=0.153 $X2=0.135
+ $Y2=0.153
r184 69 149 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r185 68 72 6.92593 $w=1.8e-08 $l=1.02e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.135 $Y2=0.153
r186 68 69 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r187 64 65 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r188 62 65 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r189 60 64 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r190 55 56 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r191 53 56 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r192 53 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r193 51 55 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r194 49 50 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r195 48 60 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r196 48 50 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r197 47 145 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r198 47 49 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.2
r199 45 46 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.1035
r200 44 145 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r201 44 46 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1035
r202 43 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r203 43 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r204 41 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r205 38 41 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r206 36 54 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.054 $Y=0.0675 $X2=0.054 $Y2=0.036
r207 33 36 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r208 31 114 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.161 $Y=0.135
+ $X2=1.161 $Y2=0.135
r209 28 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.161 $Y=0.0675 $X2=1.161 $Y2=0.135
r210 22 109 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.053 $Y=0.135
+ $X2=1.053 $Y2=0.135
r211 22 25 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.135 $X2=1.053 $Y2=0.2025
r212 16 104 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.135
+ $X2=0.837 $Y2=0.135
r213 16 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.135 $X2=0.837 $Y2=0.2025
r214 13 99 16.3636 $w=2.2e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.693 $Y2=0.135
r215 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0675 $X2=0.675 $Y2=0.135
r216 5 93 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r217 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r218 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%SE 2 5 7 10 13 15 21 31 39 42 43 51 57 58 VSS
c56 58 VSS 6.15152e-20 $X=0.567 $Y=0.1205
c57 57 VSS 0.00112348f $X=0.567 $Y=0.106
c58 51 VSS 1.82947e-19 $X=0.567 $Y=0.135
c59 43 VSS 0.00116134f $X=0.567 $Y=0.081
c60 42 VSS 0.00971257f $X=0.567 $Y=0.081
c61 39 VSS 0.009659f $X=0.243 $Y=0.081
c62 31 VSS 0.0100986f $X=0.243 $Y=0.135
c63 23 VSS 1.33806e-20 $X=0.2745 $Y=0.135
c64 22 VSS 0.00149043f $X=0.271 $Y=0.135
c65 21 VSS 1.85952e-19 $X=0.278 $Y=0.1345
c66 13 VSS 0.00121878f $X=0.567 $Y=0.135
c67 10 VSS 0.0587511f $X=0.567 $Y=0.0675
c68 5 VSS 0.00645536f $X=0.297 $Y=0.135
c69 2 VSS 0.070241f $X=0.297 $Y=0.0675
r70 57 58 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.106 $X2=0.567 $Y2=0.1205
r71 51 58 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.1205
r72 43 57 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.567 $Y2=0.106
r73 42 43 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.567 $Y=0.081 $X2=0.567
+ $Y2=0.081
r74 38 42 22 $w=1.8e-08 $l=3.24e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.567 $Y2=0.081
r75 38 39 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.081 $X2=0.243
+ $Y2=0.081
r76 30 39 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.081
r77 30 31 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.135
r78 22 23 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.271
+ $Y=0.135 $X2=0.2745 $Y2=0.135
r79 21 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.28 $Y=0.135 $X2=0.28
+ $Y2=0.135
r80 21 23 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.278
+ $Y=0.135 $X2=0.2745 $Y2=0.135
r81 19 31 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.243 $Y2=0.135
r82 19 22 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.271 $Y2=0.135
r83 13 51 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r84 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r85 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r86 5 25 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.28 $Y2=0.135
r87 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r88 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%D 2 5 7 24 VSS
c24 24 VSS 0.0118434f $X=0.459 $Y=0.1345
c25 5 VSS 0.00185098f $X=0.459 $Y=0.135
c26 2 VSS 0.0629574f $X=0.459 $Y=0.0675
r27 5 24 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r28 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r29 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%7 2 5 7 9 14 17 20 22 23 24 25 26 27 29 30 31 32
+ 35 37 38 42 44 45 52 53 56 VSS
c54 56 VSS 1.61802e-19 $X=0.351 $Y=0.072
c55 53 VSS 0.00367986f $X=0.342 $Y=0.234
c56 52 VSS 0.00194932f $X=0.351 $Y=0.234
c57 45 VSS 0.0036746f $X=0.342 $Y=0.036
c58 44 VSS 0.00199758f $X=0.351 $Y=0.036
c59 42 VSS 0.00774698f $X=0.324 $Y=0.036
c60 38 VSS 2.76819e-19 $X=0.513 $Y=0.117
c61 37 VSS 4.68887e-19 $X=0.513 $Y=0.099
c62 35 VSS 2.69498e-19 $X=0.513 $Y=0.135
c63 32 VSS 4.17962e-19 $X=0.486 $Y=0.072
c64 31 VSS 3.38584e-20 $X=0.468 $Y=0.072
c65 30 VSS 0.00175333f $X=0.418 $Y=0.072
c66 29 VSS 8.4059e-19 $X=0.378 $Y=0.072
c67 27 VSS 6.46578e-19 $X=0.504 $Y=0.072
c68 26 VSS 5.547e-19 $X=0.351 $Y=0.1845
c69 25 VSS 1.96258e-19 $X=0.351 $Y=0.144
c70 24 VSS 5.10513e-19 $X=0.351 $Y=0.126
c71 23 VSS 3.64391e-19 $X=0.351 $Y=0.099
c72 22 VSS 5.81348e-19 $X=0.351 $Y=0.225
c73 20 VSS 4.51561e-19 $X=0.351 $Y=0.063
c74 17 VSS 0.00759509f $X=0.322 $Y=0.2025
c75 12 VSS 3.78024e-19 $X=0.322 $Y=0.0675
c76 5 VSS 0.00134234f $X=0.513 $Y=0.135
c77 2 VSS 0.0585448f $X=0.513 $Y=0.0675
r78 53 54 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.3465 $Y2=0.234
r79 52 54 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.234 $X2=0.3465 $Y2=0.234
r80 49 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.342 $Y2=0.234
r81 45 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.3465 $Y2=0.036
r82 44 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.036 $X2=0.3465 $Y2=0.036
r83 41 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r84 41 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r85 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.099 $X2=0.513 $Y2=0.117
r86 35 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.117
r87 33 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.081 $X2=0.513 $Y2=0.099
r88 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.072 $X2=0.486 $Y2=0.072
r89 30 31 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.072 $X2=0.468 $Y2=0.072
r90 29 30 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.418 $Y2=0.072
r91 28 56 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.072 $X2=0.351 $Y2=0.072
r92 28 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.072 $X2=0.378 $Y2=0.072
r93 27 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.072 $X2=0.513 $Y2=0.081
r94 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.072 $X2=0.486 $Y2=0.072
r95 25 26 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.144 $X2=0.351 $Y2=0.1845
r96 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.144
r97 23 24 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.099 $X2=0.351 $Y2=0.126
r98 22 52 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.234
r99 22 26 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.1845
r100 21 56 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.072
r101 21 23 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.099
r102 20 56 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.063 $X2=0.351 $Y2=0.072
r103 19 44 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.036
r104 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.063
r105 17 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r106 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.322 $Y2=0.2025
r107 12 42 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r108 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.322 $Y2=0.0675
r109 5 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r110 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r111 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%SI 2 5 7 11 VSS
c25 11 VSS 0.0106807f $X=0.621 $Y=0.1345
c26 5 VSS 0.00120269f $X=0.621 $Y=0.135
c27 2 VSS 0.0596457f $X=0.621 $Y=0.0675
r28 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r29 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r30 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%9 2 5 7 10 13 15 17 22 25 27 29 30 39 40 46 50 51
+ 52 54 55 75 76 77 78 VSS
c78 80 VSS 1.0884e-19 $X=0.189 $Y=0.2125
c79 78 VSS 6.27945e-20 $X=0.189 $Y=0.1115
c80 77 VSS 5.52069e-19 $X=0.189 $Y=0.106
c81 76 VSS 2.10509e-19 $X=0.189 $Y=0.081
c82 75 VSS 1.53051e-19 $X=0.189 $Y=0.063
c83 55 VSS 0.00125248f $X=1.107 $Y=0.117
c84 54 VSS 0.0141151f $X=1.107 $Y=0.117
c85 52 VSS 0.00253771f $X=0.581 $Y=0.117
c86 51 VSS 0.00193299f $X=0.229 $Y=0.117
c87 50 VSS 7.51069e-19 $X=0.783 $Y=0.117
c88 46 VSS 0.00140427f $X=0.189 $Y=0.117
c89 40 VSS 0.00383164f $X=0.18 $Y=0.234
c90 39 VSS 4.95331e-19 $X=0.189 $Y=0.225
c91 38 VSS 0.00196236f $X=0.189 $Y=0.234
c92 30 VSS 0.00842362f $X=0.162 $Y=0.036
c93 29 VSS 0.00322168f $X=0.162 $Y=0.036
c94 27 VSS 0.00535983f $X=0.18 $Y=0.036
c95 25 VSS 0.00868282f $X=0.16 $Y=0.2025
c96 20 VSS 2.55988e-19 $X=0.16 $Y=0.0675
c97 13 VSS 0.001261f $X=1.107 $Y=0.135
c98 10 VSS 0.0599455f $X=1.107 $Y=0.0675
c99 5 VSS 0.00144009f $X=0.783 $Y=0.135
c100 2 VSS 0.0633669f $X=0.783 $Y=0.0675
r101 79 80 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.2 $X2=0.189 $Y2=0.2125
r102 77 78 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.106 $X2=0.189 $Y2=0.1115
r103 76 77 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.081 $X2=0.189 $Y2=0.106
r104 75 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.063 $X2=0.189 $Y2=0.081
r105 54 55 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.107 $Y=0.117 $X2=1.107
+ $Y2=0.117
r106 51 52 23.9012 $w=1.8e-08 $l=3.52e-07 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.117 $X2=0.581 $Y2=0.117
r107 49 54 22 $w=1.8e-08 $l=3.24e-07 $layer=M2 $thickness=3.6e-08 $X=0.783
+ $Y=0.117 $X2=1.107 $Y2=0.117
r108 49 52 13.716 $w=1.8e-08 $l=2.02e-07 $layer=M2 $thickness=3.6e-08 $X=0.783
+ $Y=0.117 $X2=0.581 $Y2=0.117
r109 49 50 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.783 $Y=0.117 $X2=0.783
+ $Y2=0.117
r110 46 79 5.6358 $w=1.8e-08 $l=8.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.117 $X2=0.189 $Y2=0.2
r111 46 78 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.117 $X2=0.189 $Y2=0.1115
r112 45 51 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.117 $X2=0.229 $Y2=0.117
r113 45 46 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.117 $X2=0.189
+ $Y2=0.117
r114 43 75 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r115 40 41 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r116 39 80 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.2125
r117 38 41 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r118 38 39 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.189 $Y2=0.225
r119 35 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r120 29 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r121 27 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r122 27 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.162 $Y2=0.036
r123 25 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r124 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.16 $Y2=0.2025
r125 20 30 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.162 $Y=0.0675 $X2=0.162 $Y2=0.036
r126 17 20 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.16 $Y2=0.0675
r127 13 55 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.107 $Y=0.135 $X2=1.107
+ $Y2=0.135
r128 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.135 $X2=1.107 $Y2=0.2025
r129 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.0675 $X2=1.107 $Y2=0.135
r130 5 50 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.135 $X2=0.783
+ $Y2=0.135
r131 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.135 $X2=0.783 $Y2=0.2025
r132 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0675 $X2=0.783 $Y2=0.135
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%10 4 7 9 11 16 19 21 26 29 33 36 38 40 42 43 49
+ VSS
c36 49 VSS 0.0362427f $X=0.999 $Y=0.162
c37 43 VSS 5.31938e-19 $X=0.954 $Y=0.072
c38 42 VSS 0.00378458f $X=0.936 $Y=0.072
c39 40 VSS 0.001558f $X=0.972 $Y=0.072
c40 38 VSS 8.97194e-19 $X=0.9 $Y=0.072
c41 36 VSS 6.15152e-20 $X=0.891 $Y=0.1205
c42 35 VSS 0.00121732f $X=0.891 $Y=0.106
c43 33 VSS 2.4766e-19 $X=0.891 $Y=0.135
c44 29 VSS 0.0227313f $X=1.028 $Y=0.2025
c45 26 VSS 3.25039e-19 $X=1.043 $Y=0.2025
c46 19 VSS 0.0555224f $X=1.082 $Y=0.0675
c47 16 VSS 3.25039e-19 $X=1.097 $Y=0.0675
c48 14 VSS 3.34937e-19 $X=0.97 $Y=0.0675
c49 7 VSS 0.00125164f $X=0.891 $Y=0.135
c50 4 VSS 0.0584835f $X=0.891 $Y=0.0675
r51 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.072 $X2=0.954 $Y2=0.072
r52 40 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.072 $X2=0.954 $Y2=0.072
r53 38 42 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.072 $X2=0.936 $Y2=0.072
r54 35 36 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.106 $X2=0.891 $Y2=0.1205
r55 33 36 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.135 $X2=0.891 $Y2=0.1205
r56 31 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.891 $Y=0.081 $X2=0.9 $Y2=0.072
r57 31 35 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.081 $X2=0.891 $Y2=0.106
r58 29 49 14.4321 $w=7.8e-08 $l=4.05e-08 $layer=LISD $thickness=2.8e-08 $X=0.999
+ $Y=0.2025 $X2=0.999 $Y2=0.162
r59 26 29 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.043 $Y=0.2025 $X2=1.028 $Y2=0.2025
r60 21 29 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.2025 $X2=0.97 $Y2=0.2025
r61 19 53 21.3536 $w=8.1e-08 $l=8.35e-08 $layer=LISD $thickness=2.8e-08 $X=1.082
+ $Y=0.0675 $X2=0.9985 $Y2=0.0675
r62 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.097 $Y=0.0675 $X2=1.082 $Y2=0.0675
r63 14 53 7.28836 $w=8.1e-08 $l=2.85e-08 $layer=LISD $thickness=2.8e-08 $X=0.97
+ $Y=0.0675 $X2=0.9985 $Y2=0.0675
r64 14 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.072 $X2=0.972
+ $Y2=0.072
r65 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.0675 $X2=0.97 $Y2=0.0675
r66 7 33 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.135 $X2=0.891
+ $Y2=0.135
r67 7 9 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.135 $X2=0.891 $Y2=0.2025
r68 4 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.0675 $X2=0.891 $Y2=0.135
r69 1 53 7.09296 $w=8.1e-08 $l=4.05e-08 $layer=LISD $thickness=2.8e-08 $X=0.9985
+ $Y=0.108 $X2=0.9985 $Y2=0.0675
r70 1 49 24.8571 $w=4.5e-08 $l=5.4e-08 $layer=LISD $thickness=2.8e-08 $X=0.9985
+ $Y=0.108 $X2=0.9985 $Y2=0.162
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%11 2 5 7 9 14 17 19 20 23 24 26 32 33 34 35 36 37
+ 38 40 46 47 49 50 51 54 59 VSS
c59 60 VSS 4.719e-19 $X=0.945 $Y=0.2
c60 59 VSS 0.00101748f $X=0.945 $Y=0.189
c61 58 VSS 1.67924e-19 $X=0.945 $Y=0.167
c62 54 VSS 2.26463e-19 $X=0.945 $Y=0.135
c63 52 VSS 0.00105105f $X=0.945 $Y=0.225
c64 51 VSS 0.00146362f $X=0.9 $Y=0.234
c65 50 VSS 0.00353771f $X=0.882 $Y=0.234
c66 49 VSS 0.0014995f $X=0.846 $Y=0.234
c67 48 VSS 0.00101201f $X=0.828 $Y=0.234
c68 47 VSS 0.0020447f $X=0.819 $Y=0.234
c69 46 VSS 0.00834642f $X=0.936 $Y=0.234
c70 44 VSS 1.03629e-19 $X=0.81 $Y=0.216
c71 40 VSS 5.31938e-19 $X=0.792 $Y=0.198
c72 39 VSS 2.07422e-19 $X=0.774 $Y=0.198
c73 38 VSS 4.09554e-20 $X=0.77 $Y=0.198
c74 37 VSS 8.20366e-20 $X=0.767 $Y=0.198
c75 36 VSS 6.34818e-19 $X=0.756 $Y=0.198
c76 35 VSS 7.00738e-19 $X=0.801 $Y=0.198
c77 34 VSS 2.66851e-19 $X=0.747 $Y=0.178
c78 33 VSS 1.28225e-19 $X=0.747 $Y=0.167
c79 32 VSS 9.95178e-19 $X=0.747 $Y=0.164
c80 26 VSS 4.68208e-19 $X=0.747 $Y=0.09
c81 24 VSS 2.54721e-19 $X=0.747 $Y=0.189
c82 23 VSS 0.00458934f $X=0.81 $Y=0.2025
c83 19 VSS 6.04398e-19 $X=0.827 $Y=0.2025
c84 17 VSS 0.0144192f $X=0.758 $Y=0.0675
c85 14 VSS 3.25039e-19 $X=0.773 $Y=0.0675
c86 12 VSS 6.23621e-19 $X=0.7 $Y=0.0675
c87 5 VSS 0.0014001f $X=0.945 $Y=0.135
c88 2 VSS 0.0619707f $X=0.945 $Y=0.0675
r89 59 60 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.189 $X2=0.945 $Y2=0.2
r90 58 59 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.167 $X2=0.945 $Y2=0.189
r91 57 58 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.164 $X2=0.945 $Y2=0.167
r92 54 57 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.135 $X2=0.945 $Y2=0.164
r93 52 60 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.2
r94 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.234 $X2=0.9 $Y2=0.234
r95 49 50 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.234 $X2=0.882 $Y2=0.234
r96 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.846 $Y2=0.234
r97 47 48 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.819
+ $Y=0.234 $X2=0.828 $Y2=0.234
r98 46 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r99 46 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.9 $Y2=0.234
r100 42 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.81 $Y=0.225 $X2=0.819 $Y2=0.234
r101 42 44 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.225 $X2=0.81 $Y2=0.216
r102 41 44 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.207 $X2=0.81 $Y2=0.216
r103 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.198 $X2=0.792 $Y2=0.198
r104 38 39 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.77
+ $Y=0.198 $X2=0.774 $Y2=0.198
r105 37 38 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.767
+ $Y=0.198 $X2=0.77 $Y2=0.198
r106 36 37 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.198 $X2=0.767 $Y2=0.198
r107 35 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.801 $Y=0.198 $X2=0.81 $Y2=0.207
r108 35 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.198 $X2=0.792 $Y2=0.198
r109 33 34 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.167 $X2=0.747 $Y2=0.178
r110 32 33 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.164 $X2=0.747 $Y2=0.167
r111 31 32 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.121 $X2=0.747 $Y2=0.164
r112 26 31 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.09 $X2=0.747 $Y2=0.121
r113 24 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.747 $Y=0.189 $X2=0.756 $Y2=0.198
r114 24 34 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.189 $X2=0.747 $Y2=0.178
r115 23 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.216 $X2=0.81
+ $Y2=0.216
r116 20 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2025 $X2=0.81 $Y2=0.2025
r117 19 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.2025 $X2=0.81 $Y2=0.2025
r118 17 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.747 $Y=0.09 $X2=0.747
+ $Y2=0.09
r119 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.758 $Y2=0.0675
r120 12 17 12.0194 $w=8.1e-08 $l=4.7e-08 $layer=LISD $thickness=2.8e-08 $X=0.7
+ $Y=0.0675 $X2=0.747 $Y2=0.0675
r121 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.0675 $X2=0.7 $Y2=0.0675
r122 5 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.945 $Y=0.135 $X2=0.945
+ $Y2=0.135
r123 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.945
+ $Y=0.135 $X2=0.945 $Y2=0.2025
r124 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.945
+ $Y=0.0675 $X2=0.945 $Y2=0.135
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%12 2 5 7 9 12 14 17 19 21 25 27 32 36 37 38 43 44
+ VSS
c31 44 VSS 2.89087e-19 $X=1.314 $Y=0.09
c32 43 VSS 1.16913e-19 $X=1.323 $Y=0.09
c33 38 VSS 1.92014e-19 $X=1.323 $Y=0.144
c34 37 VSS 2.83021e-19 $X=1.323 $Y=0.126
c35 36 VSS 4.65462e-19 $X=1.323 $Y=0.182
c36 34 VSS 1.81242e-20 $X=1.2915 $Y=0.191
c37 33 VSS 2.15286e-20 $X=1.287 $Y=0.191
c38 32 VSS 0.00127461f $X=1.283 $Y=0.191
c39 31 VSS 7.15474e-19 $X=1.242 $Y=0.191
c40 27 VSS 5.27395e-20 $X=1.224 $Y=0.191
c41 26 VSS 3.73006e-19 $X=1.314 $Y=0.191
c42 25 VSS 2.89178e-19 $X=1.215 $Y=0.163
c43 21 VSS 1.79849e-19 $X=1.215 $Y=0.135
c44 19 VSS 7.49026e-19 $X=1.215 $Y=0.182
c45 17 VSS 0.00885042f $X=1.294 $Y=0.2025
c46 12 VSS 0.0205477f $X=1.294 $Y=0.0675
c47 5 VSS 0.00122128f $X=1.215 $Y=0.135
c48 2 VSS 0.0583406f $X=1.215 $Y=0.0675
r49 44 45 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.314
+ $Y=0.09 $X2=1.3185 $Y2=0.09
r50 43 45 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.09 $X2=1.3185 $Y2=0.09
r51 40 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.09 $X2=1.314 $Y2=0.09
r52 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.126 $X2=1.323 $Y2=0.144
r53 36 38 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.182 $X2=1.323 $Y2=0.144
r54 35 43 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.099 $X2=1.323 $Y2=0.09
r55 35 37 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.099 $X2=1.323 $Y2=0.126
r56 33 34 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.287
+ $Y=0.191 $X2=1.2915 $Y2=0.191
r57 32 33 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=1.283
+ $Y=0.191 $X2=1.287 $Y2=0.191
r58 31 32 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.242
+ $Y=0.191 $X2=1.283 $Y2=0.191
r59 29 34 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.191 $X2=1.2915 $Y2=0.191
r60 27 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.224
+ $Y=0.191 $X2=1.242 $Y2=0.191
r61 26 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.314 $Y=0.191 $X2=1.323 $Y2=0.182
r62 26 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.314
+ $Y=0.191 $X2=1.296 $Y2=0.191
r63 24 25 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.144 $X2=1.215 $Y2=0.163
r64 21 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.135 $X2=1.215 $Y2=0.144
r65 19 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.215 $Y=0.182 $X2=1.224 $Y2=0.191
r66 19 25 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.182 $X2=1.215 $Y2=0.163
r67 17 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.191 $X2=1.296
+ $Y2=0.191
r68 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.279 $Y=0.2025 $X2=1.294 $Y2=0.2025
r69 12 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.09 $X2=1.296
+ $Y2=0.09
r70 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.279 $Y=0.0675 $X2=1.294 $Y2=0.0675
r71 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.215 $Y=0.135 $X2=1.215
+ $Y2=0.135
r72 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.215
+ $Y=0.135 $X2=1.215 $Y2=0.2025
r73 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.215
+ $Y=0.0675 $X2=1.215 $Y2=0.135
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%13 2 5 7 10 15 18 23 26 31 34 37 39 41 42 46 47 50
+ 51 53 59 60 61 62 63 66 67 72 73 74 77 80 81 82 83 86 87 90 91 92 94 105 107
+ 110 VSS
c67 110 VSS 2.79962e-19 $X=1.377 $Y=0.135
c68 108 VSS 4.98311e-20 $X=1.2645 $Y=0.135
c69 107 VSS 3.49116e-19 $X=1.26 $Y=0.135
c70 105 VSS 5.14517e-19 $X=1.269 $Y=0.135
c71 101 VSS 0.00253921f $X=1.251 $Y=0.036
c72 97 VSS 0.00331528f $X=1.431 $Y=0.135
c73 94 VSS 0.00474203f $X=1.377 $Y=0.225
c74 92 VSS 0.00144937f $X=1.377 $Y=0.1035
c75 91 VSS 0.00219086f $X=1.377 $Y=0.081
c76 90 VSS 0.00103511f $X=1.377 $Y=0.126
c77 88 VSS 0.00208651f $X=1.35 $Y=0.036
c78 87 VSS 0.00350381f $X=1.332 $Y=0.036
c79 86 VSS 3.87876e-19 $X=1.287 $Y=0.036
c80 85 VSS 0.00192765f $X=1.283 $Y=0.036
c81 83 VSS 0.00526264f $X=1.368 $Y=0.036
c82 82 VSS 4.91035e-19 $X=1.251 $Y=0.116
c83 81 VSS 2.41096e-19 $X=1.251 $Y=0.106
c84 80 VSS 7.80213e-19 $X=1.251 $Y=0.099
c85 79 VSS 4.80483e-19 $X=1.251 $Y=0.081
c86 78 VSS 4.9709e-19 $X=1.251 $Y=0.07
c87 77 VSS 0.00124273f $X=1.251 $Y=0.063
c88 76 VSS 1.26074e-19 $X=1.251 $Y=0.126
c89 74 VSS 0.00146362f $X=1.224 $Y=0.036
c90 73 VSS 0.00333697f $X=1.206 $Y=0.036
c91 72 VSS 0.00146362f $X=1.17 $Y=0.036
c92 71 VSS 0.00251494f $X=1.152 $Y=0.036
c93 67 VSS 0.0045992f $X=1.134 $Y=0.036
c94 66 VSS 0.00224226f $X=1.134 $Y=0.036
c95 64 VSS 0.00328022f $X=1.242 $Y=0.036
c96 63 VSS 0.0129562f $X=1.332 $Y=0.234
c97 62 VSS 0.00350786f $X=1.206 $Y=0.234
c98 61 VSS 0.00141253f $X=1.17 $Y=0.234
c99 60 VSS 0.00310297f $X=1.152 $Y=0.234
c100 59 VSS 0.00146362f $X=1.116 $Y=0.234
c101 58 VSS 0.00245593f $X=1.098 $Y=0.234
c102 53 VSS 0.00215392f $X=1.08 $Y=0.234
c103 51 VSS 0.00775972f $X=1.368 $Y=0.234
c104 50 VSS 0.00362692f $X=1.08 $Y=0.2025
c105 46 VSS 5.38922e-19 $X=1.097 $Y=0.2025
c106 41 VSS 5.38922e-19 $X=1.151 $Y=0.0675
c107 37 VSS 0.0148754f $X=1.593 $Y=0.135
c108 34 VSS 0.0645347f $X=1.593 $Y=0.0675
c109 26 VSS 0.0644226f $X=1.539 $Y=0.0675
c110 18 VSS 0.0644226f $X=1.485 $Y=0.0675
c111 10 VSS 0.0650932f $X=1.431 $Y=0.0675
c112 5 VSS 0.00193244f $X=1.269 $Y=0.135
c113 2 VSS 0.0615704f $X=1.269 $Y=0.0675
r114 107 108 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.26
+ $Y=0.135 $X2=1.2645 $Y2=0.135
r115 105 108 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.269 $Y=0.135 $X2=1.2645 $Y2=0.135
r116 102 107 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.135 $X2=1.26 $Y2=0.135
r117 95 110 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.386
+ $Y=0.135 $X2=1.377 $Y2=0.135
r118 95 97 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.386
+ $Y=0.135 $X2=1.431 $Y2=0.135
r119 93 110 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.144 $X2=1.377 $Y2=0.135
r120 93 94 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.144 $X2=1.377 $Y2=0.225
r121 91 92 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.081 $X2=1.377 $Y2=0.1035
r122 90 110 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.126 $X2=1.377 $Y2=0.135
r123 90 92 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.126 $X2=1.377 $Y2=0.1035
r124 89 91 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.045 $X2=1.377 $Y2=0.081
r125 87 88 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.332
+ $Y=0.036 $X2=1.35 $Y2=0.036
r126 86 87 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.287
+ $Y=0.036 $X2=1.332 $Y2=0.036
r127 85 86 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=1.283
+ $Y=0.036 $X2=1.287 $Y2=0.036
r128 84 101 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.26
+ $Y=0.036 $X2=1.251 $Y2=0.036
r129 84 85 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.26
+ $Y=0.036 $X2=1.283 $Y2=0.036
r130 83 89 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.368 $Y=0.036 $X2=1.377 $Y2=0.045
r131 83 88 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.368
+ $Y=0.036 $X2=1.35 $Y2=0.036
r132 81 82 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.106 $X2=1.251 $Y2=0.116
r133 80 81 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.099 $X2=1.251 $Y2=0.106
r134 79 80 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.081 $X2=1.251 $Y2=0.099
r135 78 79 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.07 $X2=1.251 $Y2=0.081
r136 77 78 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.063 $X2=1.251 $Y2=0.07
r137 76 102 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.126 $X2=1.251 $Y2=0.135
r138 76 82 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.126 $X2=1.251 $Y2=0.116
r139 75 101 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.045 $X2=1.251 $Y2=0.036
r140 75 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.045 $X2=1.251 $Y2=0.063
r141 73 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.206
+ $Y=0.036 $X2=1.224 $Y2=0.036
r142 72 73 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.17
+ $Y=0.036 $X2=1.206 $Y2=0.036
r143 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.152
+ $Y=0.036 $X2=1.17 $Y2=0.036
r144 66 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.036 $X2=1.152 $Y2=0.036
r145 66 67 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.134 $Y=0.036
+ $X2=1.134 $Y2=0.036
r146 64 101 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.242
+ $Y=0.036 $X2=1.251 $Y2=0.036
r147 64 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.242
+ $Y=0.036 $X2=1.224 $Y2=0.036
r148 62 63 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M1 $thickness=3.6e-08 $X=1.206
+ $Y=0.234 $X2=1.332 $Y2=0.234
r149 61 62 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.17
+ $Y=0.234 $X2=1.206 $Y2=0.234
r150 60 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.152
+ $Y=0.234 $X2=1.17 $Y2=0.234
r151 59 60 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.116
+ $Y=0.234 $X2=1.152 $Y2=0.234
r152 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.234 $X2=1.116 $Y2=0.234
r153 53 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.098 $Y2=0.234
r154 51 94 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.368 $Y=0.234 $X2=1.377 $Y2=0.225
r155 51 63 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.368
+ $Y=0.234 $X2=1.332 $Y2=0.234
r156 50 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234 $X2=1.08
+ $Y2=0.234
r157 47 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2025 $X2=1.08 $Y2=0.2025
r158 46 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.097 $Y=0.2025 $X2=1.08 $Y2=0.2025
r159 45 67 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=1.134 $Y=0.0675 $X2=1.134 $Y2=0.036
r160 42 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.117 $Y=0.0675 $X2=1.134 $Y2=0.0675
r161 41 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.151 $Y=0.0675 $X2=1.134 $Y2=0.0675
r162 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.593 $Y=0.135 $X2=1.593 $Y2=0.2025
r163 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.593 $Y=0.0675 $X2=1.593 $Y2=0.135
r164 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.539
+ $Y=0.135 $X2=1.593 $Y2=0.135
r165 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.539 $Y=0.135 $X2=1.539 $Y2=0.2025
r166 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.539 $Y=0.0675 $X2=1.539 $Y2=0.135
r167 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.485
+ $Y=0.135 $X2=1.539 $Y2=0.135
r168 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.485 $Y=0.135 $X2=1.485 $Y2=0.2025
r169 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.485 $Y=0.0675 $X2=1.485 $Y2=0.135
r170 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.431
+ $Y=0.135 $X2=1.485 $Y2=0.135
r171 13 97 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.431 $Y=0.135 $X2=1.431
+ $Y2=0.135
r172 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.431 $Y=0.135 $X2=1.431 $Y2=0.2025
r173 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.431 $Y=0.0675 $X2=1.431 $Y2=0.135
r174 5 105 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.269 $Y=0.135 $X2=1.269
+ $Y2=0.135
r175 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.269
+ $Y=0.135 $X2=1.269 $Y2=0.2025
r176 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.269
+ $Y=0.0675 $X2=1.269 $Y2=0.135
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%15 1 4 6 7 10 11 14 23 24 26 27 28 30 33 34 35 36
+ 37 VSS
c32 37 VSS 8.46035e-21 $X=0.63 $Y=0.198
c33 36 VSS 1.62375e-19 $X=0.612 $Y=0.198
c34 35 VSS 9.14524e-20 $X=0.599 $Y=0.198
c35 34 VSS 3.12342e-19 $X=0.58 $Y=0.198
c36 33 VSS 5.31938e-19 $X=0.576 $Y=0.198
c37 32 VSS 0.00134307f $X=0.558 $Y=0.198
c38 30 VSS 5.86427e-19 $X=0.648 $Y=0.198
c39 28 VSS 3.95078e-19 $X=0.531 $Y=0.198
c40 27 VSS 5.17397e-19 $X=0.522 $Y=0.198
c41 26 VSS 0.00400558f $X=0.504 $Y=0.198
c42 25 VSS 4.26131e-19 $X=0.468 $Y=0.198
c43 24 VSS 1.4604e-19 $X=0.459 $Y=0.198
c44 23 VSS 5.61374e-19 $X=0.45 $Y=0.198
c45 14 VSS 0.00375596f $X=0.646 $Y=0.2025
c46 10 VSS 0.00555436f $X=0.54 $Y=0.2025
c47 6 VSS 6.69874e-19 $X=0.557 $Y=0.2025
c48 4 VSS 0.00689207f $X=0.434 $Y=0.2025
c49 1 VSS 2.69461e-19 $X=0.449 $Y=0.2025
r50 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.198 $X2=0.63 $Y2=0.198
r51 35 36 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.599
+ $Y=0.198 $X2=0.612 $Y2=0.198
r52 34 35 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.58
+ $Y=0.198 $X2=0.599 $Y2=0.198
r53 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.198 $X2=0.58 $Y2=0.198
r54 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.198 $X2=0.576 $Y2=0.198
r55 30 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.198 $X2=0.63 $Y2=0.198
r56 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.198 $X2=0.531 $Y2=0.198
r57 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.198 $X2=0.522 $Y2=0.198
r58 25 26 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.198 $X2=0.504 $Y2=0.198
r59 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.198 $X2=0.468 $Y2=0.198
r60 23 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.198 $X2=0.459 $Y2=0.198
r61 21 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.198 $X2=0.558 $Y2=0.198
r62 21 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.198 $X2=0.531 $Y2=0.198
r63 17 23 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.45 $Y2=0.198
r64 14 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.198 $X2=0.648
+ $Y2=0.198
r65 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.646 $Y2=0.2025
r66 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.198 $X2=0.54
+ $Y2=0.198
r67 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r68 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r69 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r70 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.449
+ $Y=0.2025 $X2=0.434 $Y2=0.2025
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%16 1 2 5 6 9 16 18 19 20 21 23 VSS
c26 23 VSS 7.00634e-19 $X=0.747 $Y=0.234
c27 22 VSS 0.00298267f $X=0.738 $Y=0.234
c28 21 VSS 0.00103868f $X=0.711 $Y=0.234
c29 20 VSS 0.00157473f $X=0.702 $Y=0.234
c30 19 VSS 0.00206804f $X=0.684 $Y=0.234
c31 18 VSS 0.00706733f $X=0.662 $Y=0.234
c32 16 VSS 0.00225063f $X=0.756 $Y=0.234
c33 9 VSS 0.00363839f $X=0.758 $Y=0.2025
c34 6 VSS 7.37037e-19 $X=0.773 $Y=0.2025
c35 5 VSS 0.00358468f $X=0.594 $Y=0.2025
c36 1 VSS 6.32999e-19 $X=0.611 $Y=0.2025
r37 22 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.234 $X2=0.747 $Y2=0.234
r38 21 22 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.711
+ $Y=0.234 $X2=0.738 $Y2=0.234
r39 20 21 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.234 $X2=0.711 $Y2=0.234
r40 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.234 $X2=0.702 $Y2=0.234
r41 18 19 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.662
+ $Y=0.234 $X2=0.684 $Y2=0.234
r42 16 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.747 $Y2=0.234
r43 12 18 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.662 $Y2=0.234
r44 9 16 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234 $X2=0.756
+ $Y2=0.234
r45 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2025 $X2=0.758 $Y2=0.2025
r46 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r47 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.577
+ $Y=0.2025 $X2=0.594 $Y2=0.2025
r48 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.611
+ $Y=0.2025 $X2=0.594 $Y2=0.2025
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%QN 1 2 6 7 11 12 15 16 17 20 21 23 24 30 31 33 44
+ 45 VSS
c19 48 VSS 0.00300284f $X=1.6465 $Y=0.1845
c20 46 VSS 2.62283e-19 $X=1.6465 $Y=0.13025
c21 45 VSS 0.00548083f $X=1.6465 $Y=0.126
c22 44 VSS 6.00307e-19 $X=1.646 $Y=0.1345
c23 42 VSS 0.00247012f $X=1.6465 $Y=0.225
c24 33 VSS 0.00155282f $X=1.458 $Y=0.234
c25 31 VSS 0.0249971f $X=1.637 $Y=0.234
c26 30 VSS 0.00929647f $X=1.566 $Y=0.036
c27 24 VSS 0.00904424f $X=1.458 $Y=0.036
c28 23 VSS 0.00155282f $X=1.458 $Y=0.036
c29 21 VSS 0.0249971f $X=1.637 $Y=0.036
c30 20 VSS 0.00929647f $X=1.566 $Y=0.2025
c31 16 VSS 5.38922e-19 $X=1.583 $Y=0.2025
c32 15 VSS 0.00918054f $X=1.458 $Y=0.2025
c33 11 VSS 5.72268e-19 $X=1.475 $Y=0.2025
c34 6 VSS 5.38922e-19 $X=1.583 $Y=0.0675
c35 1 VSS 5.72268e-19 $X=1.475 $Y=0.0675
r36 47 48 2.57237 $w=1.9e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.144 $X2=1.6465 $Y2=0.1845
r37 45 46 0.26994 $w=1.9e-08 $l=4.25e-09 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.126 $X2=1.6465 $Y2=0.13025
r38 44 47 0.603395 $w=1.9e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.1345 $X2=1.6465 $Y2=0.144
r39 44 46 0.26994 $w=1.9e-08 $l=4.25e-09 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.1345 $X2=1.6465 $Y2=0.13025
r40 42 48 2.57237 $w=1.9e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.225 $X2=1.6465 $Y2=0.1845
r41 41 45 5.14474 $w=1.9e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.045 $X2=1.6465 $Y2=0.126
r42 33 39 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.458
+ $Y=0.234 $X2=1.566 $Y2=0.234
r43 31 42 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.637 $Y=0.234 $X2=1.6465 $Y2=0.225
r44 31 39 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.637
+ $Y=0.234 $X2=1.566 $Y2=0.234
r45 29 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.566 $Y=0.036 $X2=1.566
+ $Y2=0.036
r46 23 29 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.458
+ $Y=0.036 $X2=1.566 $Y2=0.036
r47 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.458 $Y=0.036 $X2=1.458
+ $Y2=0.036
r48 21 41 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.637 $Y=0.036 $X2=1.6465 $Y2=0.045
r49 21 29 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.637
+ $Y=0.036 $X2=1.566 $Y2=0.036
r50 20 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.566 $Y=0.234 $X2=1.566
+ $Y2=0.234
r51 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.549 $Y=0.2025 $X2=1.566 $Y2=0.2025
r52 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.583 $Y=0.2025 $X2=1.566 $Y2=0.2025
r53 15 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.458 $Y=0.234 $X2=1.458
+ $Y2=0.234
r54 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.441 $Y=0.2025 $X2=1.458 $Y2=0.2025
r55 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.475 $Y=0.2025 $X2=1.458 $Y2=0.2025
r56 10 30 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.566
+ $Y=0.0675 $X2=1.566 $Y2=0.036
r57 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.549 $Y=0.0675 $X2=1.566 $Y2=0.0675
r58 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.583 $Y=0.0675 $X2=1.566 $Y2=0.0675
r59 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.458
+ $Y=0.0675 $X2=1.458 $Y2=0.036
r60 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.441
+ $Y=0.0675 $X2=1.458 $Y2=0.0675
r61 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.475
+ $Y=0.0675 $X2=1.458 $Y2=0.0675
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%18 1 6 9 VSS
c11 9 VSS 0.0193928f $X=0.866 $Y=0.0675
c12 6 VSS 3.25039e-19 $X=0.881 $Y=0.0675
c13 4 VSS 3.25039e-19 $X=0.808 $Y=0.0675
r14 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.881
+ $Y=0.0675 $X2=0.866 $Y2=0.0675
r15 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.808
+ $Y=0.0675 $X2=0.866 $Y2=0.0675
r16 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.793
+ $Y=0.0675 $X2=0.808 $Y2=0.0675
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%19 1 6 9 VSS
c13 9 VSS 0.0132338f $X=1.19 $Y=0.2025
c14 6 VSS 3.22787e-19 $X=1.205 $Y=0.2025
c15 4 VSS 3.14547e-19 $X=1.132 $Y=0.2025
r16 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=1.205
+ $Y=0.2025 $X2=1.19 $Y2=0.2025
r17 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=1.132
+ $Y=0.2025 $X2=1.19 $Y2=0.2025
r18 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=1.117
+ $Y=0.2025 $X2=1.132 $Y2=0.2025
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%22 1 2 VSS
c1 1 VSS 0.00183233f $X=1.205 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=1.205
+ $Y=0.0675 $X2=1.171 $Y2=0.0675
.ends

.subckt PM_SDFHX4_ASAP7_75T_SRAM%23 1 2 VSS
c1 1 VSS 0.00183233f $X=0.881 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.881
+ $Y=0.2025 $X2=0.847 $Y2=0.2025
.ends


* END of "./SDFHx4_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt SDFHx4_ASAP7_75t_SRAM  VSS VDD CLK SE D SI QN
* 
* QN	QN
* SI	SI
* D	D
* SE	SE
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_9_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_7_M2_d N_SE_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 noxref_20 N_D_M3_g noxref_14 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M4 VSS N_7_M4_g noxref_20 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M5 noxref_21 N_SE_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M6 noxref_14 N_SI_M6_g noxref_21 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M7 N_11_M7_d N_4_M7_g noxref_14 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M8 N_18_M8_d N_9_M8_g N_11_M8_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.027
M9 VSS N_10_M9_g N_18_M9_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.027
M10 N_10_M10_d N_11_M10_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.027
M11 N_13_M11_d N_9_M11_g N_10_M11_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=1.097 $Y=0.027
M12 N_22_M12_d N_4_M12_g N_13_M12_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=1.151 $Y=0.027
M13 VSS N_12_M13_g N_22_M13_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.027
M14 N_12_M14_d N_13_M14_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M15 N_QN_M15_d N_13_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.421
+ $Y=0.027
M16 N_QN_M16_d N_13_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.475
+ $Y=0.027
M17 N_QN_M17_d N_13_M17_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.529
+ $Y=0.027
M18 N_QN_M18_d N_13_M18_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.583
+ $Y=0.027
M19 VDD N_CLK_M19_g N_4_M19_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M20 N_9_M20_d N_4_M20_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M21 N_7_M21_d N_SE_M21_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M22 VDD N_D_M22_g N_15_M22_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M23 N_15_M23_d N_7_M23_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M24 N_16_M24_d N_SE_M24_g N_15_M24_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M25 N_15_M25_d N_SI_M25_g N_16_M25_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.611 $Y=0.162
M26 N_11_M26_d N_9_M26_g N_16_M26_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.773 $Y=0.162
M27 N_23_M27_d N_4_M27_g N_11_M27_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.827 $Y=0.162
M28 VDD N_10_M28_g N_23_M28_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.162
M29 N_10_M29_d N_11_M29_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.162
M30 N_13_M30_d N_4_M30_g N_10_M30_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=1.043 $Y=0.162
M31 N_19_M31_d N_9_M31_g N_13_M31_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=1.097 $Y=0.162
M32 VDD N_12_M32_g N_19_M32_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.162
M33 N_12_M33_d N_13_M33_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
M34 N_QN_M34_d N_13_M34_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.421
+ $Y=0.162
M35 N_QN_M35_d N_13_M35_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.475
+ $Y=0.162
M36 N_QN_M36_d N_13_M36_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.529
+ $Y=0.162
M37 N_QN_M37_d N_13_M37_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.583
+ $Y=0.162
*
* 
* .include "SDFHx4_ASAP7_75t_SRAM.pex.sp.SDFHX4_ASAP7_75T_SRAM.pxi"
* BEGIN of "./SDFHx4_ASAP7_75t_SRAM.pex.sp.SDFHX4_ASAP7_75T_SRAM.pxi"
* File: SDFHx4_ASAP7_75t_SRAM.pex.sp.SDFHX4_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 13:04:10 2017
* 
x_PM_SDFHX4_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M19_g CLK VSS
+ PM_SDFHX4_ASAP7_75T_SRAM%CLK
x_PM_SDFHX4_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_15_n N_4_M20_g N_4_M7_g N_4_c_45_p
+ N_4_M27_g N_4_c_48_p N_4_M30_g N_4_M12_g N_4_c_51_p N_4_M0_s N_4_M19_s
+ N_4_c_16_n N_4_c_17_n N_4_c_18_n N_4_c_19_n N_4_c_20_n N_4_c_22_n N_4_c_60_p
+ N_4_c_23_n N_4_c_24_n N_4_c_27_p N_4_c_112_p N_4_c_31_p N_4_c_120_p N_4_c_25_n
+ N_4_c_39_p N_4_c_43_p N_4_c_65_p N_4_c_72_p N_4_c_73_p VSS
+ PM_SDFHX4_ASAP7_75T_SRAM%4
x_PM_SDFHX4_ASAP7_75T_SRAM%SE N_SE_M2_g N_SE_c_143_n N_SE_M21_g N_SE_M5_g
+ N_SE_c_153_p N_SE_M24_g SE N_SE_c_146_n N_SE_c_154_p N_SE_c_147_n N_SE_c_159_p
+ N_SE_c_148_n N_SE_c_166_p N_SE_c_167_p VSS PM_SDFHX4_ASAP7_75T_SRAM%SE
x_PM_SDFHX4_ASAP7_75T_SRAM%D N_D_M3_g N_D_c_202_n N_D_M22_g D VSS
+ PM_SDFHX4_ASAP7_75T_SRAM%D
x_PM_SDFHX4_ASAP7_75T_SRAM%7 N_7_M4_g N_7_c_228_n N_7_M23_g N_7_M2_d N_7_M21_d
+ N_7_c_223_n N_7_c_229_n N_7_c_250_n N_7_c_230_n N_7_c_251_n N_7_c_231_n
+ N_7_c_224_n N_7_c_233_n N_7_c_235_n N_7_c_236_n N_7_c_237_n N_7_c_238_n
+ N_7_c_225_n N_7_c_240_n N_7_c_242_n N_7_c_243_n N_7_c_273_p N_7_c_244_n
+ N_7_c_259_n N_7_c_226_n N_7_c_247_n VSS PM_SDFHX4_ASAP7_75T_SRAM%7
x_PM_SDFHX4_ASAP7_75T_SRAM%SI N_SI_M6_g N_SI_c_278_n N_SI_M25_g SI VSS
+ PM_SDFHX4_ASAP7_75T_SRAM%SI
x_PM_SDFHX4_ASAP7_75T_SRAM%9 N_9_M8_g N_9_c_305_n N_9_M26_g N_9_M11_g N_9_c_309_n
+ N_9_M31_g N_9_M1_d N_9_M20_d N_9_c_311_n N_9_c_337_n N_9_c_314_n N_9_c_317_n
+ N_9_c_338_n N_9_c_319_n N_9_c_321_n N_9_c_323_n N_9_c_325_n N_9_c_327_n
+ N_9_c_328_n N_9_c_333_n N_9_c_347_n N_9_c_302_n N_9_c_349_n N_9_c_336_n VSS
+ PM_SDFHX4_ASAP7_75T_SRAM%9
x_PM_SDFHX4_ASAP7_75T_SRAM%10 N_10_M9_g N_10_c_381_n N_10_M28_g N_10_M10_d
+ N_10_M11_s N_10_c_382_n N_10_M29_d N_10_M30_s N_10_c_385_n N_10_c_387_n
+ N_10_c_395_n N_10_c_388_n N_10_c_396_n N_10_c_397_n N_10_c_400_p N_10_c_389_n
+ VSS PM_SDFHX4_ASAP7_75T_SRAM%10
x_PM_SDFHX4_ASAP7_75T_SRAM%11 N_11_M10_g N_11_c_418_n N_11_M29_g N_11_M7_d
+ N_11_M8_s N_11_c_419_n N_11_M27_s N_11_M26_d N_11_c_422_n N_11_c_461_p
+ N_11_c_436_n N_11_c_423_n N_11_c_425_n N_11_c_457_p N_11_c_426_n N_11_c_458_p
+ N_11_c_427_n N_11_c_466_p N_11_c_443_n N_11_c_428_n N_11_c_469_p N_11_c_429_n
+ N_11_c_431_n N_11_c_449_n N_11_c_432_n N_11_c_434_n VSS
+ PM_SDFHX4_ASAP7_75T_SRAM%11
x_PM_SDFHX4_ASAP7_75T_SRAM%12 N_12_M13_g N_12_c_476_n N_12_M32_g N_12_M14_d
+ N_12_c_487_p N_12_M33_d N_12_c_485_p N_12_c_477_n N_12_c_478_n N_12_c_479_n
+ N_12_c_486_p N_12_c_482_p N_12_c_500_p N_12_c_492_p N_12_c_501_p N_12_c_499_p
+ N_12_c_491_p VSS PM_SDFHX4_ASAP7_75T_SRAM%12
x_PM_SDFHX4_ASAP7_75T_SRAM%13 N_13_M14_g N_13_c_526_n N_13_M33_g N_13_M15_g
+ N_13_M34_g N_13_M16_g N_13_M35_g N_13_M17_g N_13_M36_g N_13_M18_g N_13_c_547_p
+ N_13_M37_g N_13_M12_s N_13_M11_d N_13_M31_s N_13_M30_d N_13_c_507_n
+ N_13_c_564_p N_13_c_509_n N_13_c_516_n N_13_c_511_n N_13_c_512_n N_13_c_569_p
+ N_13_c_527_n N_13_c_522_n N_13_c_513_n N_13_c_514_n N_13_c_571_p N_13_c_531_n
+ N_13_c_533_n N_13_c_534_n N_13_c_535_n N_13_c_536_n N_13_c_557_p N_13_c_537_n
+ N_13_c_538_n N_13_c_540_n N_13_c_541_n N_13_c_542_n N_13_c_543_n N_13_c_544_n
+ N_13_c_545_n N_13_c_546_n VSS PM_SDFHX4_ASAP7_75T_SRAM%13
x_PM_SDFHX4_ASAP7_75T_SRAM%15 N_15_M22_s N_15_c_573_n N_15_M24_s N_15_M23_d
+ N_15_c_574_n N_15_M25_d N_15_c_575_n N_15_c_576_n N_15_c_586_n N_15_c_577_n
+ N_15_c_588_n N_15_c_578_n N_15_c_579_n N_15_c_581_n N_15_c_580_n N_15_c_599_p
+ N_15_c_600_p N_15_c_591_n VSS PM_SDFHX4_ASAP7_75T_SRAM%15
x_PM_SDFHX4_ASAP7_75T_SRAM%16 N_16_M25_s N_16_M24_d N_16_c_605_n N_16_M26_s
+ N_16_c_611_n N_16_c_619_n N_16_c_610_n N_16_c_606_n N_16_c_608_n N_16_c_609_n
+ N_16_c_622_n VSS PM_SDFHX4_ASAP7_75T_SRAM%16
x_PM_SDFHX4_ASAP7_75T_SRAM%QN N_QN_M16_d N_QN_M15_d N_QN_M18_d N_QN_M17_d
+ N_QN_M35_d N_QN_M34_d N_QN_c_634_n N_QN_M37_d N_QN_M36_d N_QN_c_636_n
+ N_QN_c_637_n N_QN_c_640_n N_QN_c_642_n N_QN_c_643_n N_QN_c_644_n N_QN_c_647_n
+ QN N_QN_c_649_n VSS PM_SDFHX4_ASAP7_75T_SRAM%QN
x_PM_SDFHX4_ASAP7_75T_SRAM%18 N_18_M8_d N_18_M9_s N_18_c_650_n VSS
+ PM_SDFHX4_ASAP7_75T_SRAM%18
x_PM_SDFHX4_ASAP7_75T_SRAM%19 N_19_M31_d N_19_M32_s N_19_c_661_n VSS
+ PM_SDFHX4_ASAP7_75T_SRAM%19
x_PM_SDFHX4_ASAP7_75T_SRAM%22 N_22_M13_s N_22_M12_d VSS PM_SDFHX4_ASAP7_75T_SRAM%22
x_PM_SDFHX4_ASAP7_75T_SRAM%23 N_23_M28_s N_23_M27_d VSS PM_SDFHX4_ASAP7_75T_SRAM%23
cc_1 N_CLK_M0_g N_4_M1_g 0.00287079f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_CLK_c_2_p N_4_c_15_n 0.00101351f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 CLK N_4_c_16_n 0.00120883f $X=0.081 $Y=0.1345 $X2=0.056 $Y2=0.2025
cc_4 CLK N_4_c_17_n 0.00119149f $X=0.081 $Y=0.1345 $X2=0.018 $Y2=0.144
cc_5 CLK N_4_c_18_n 0.00119149f $X=0.081 $Y=0.1345 $X2=0.018 $Y2=0.1035
cc_6 CLK N_4_c_19_n 9.60838e-19 $X=0.081 $Y=0.1345 $X2=0.018 $Y2=0.2
cc_7 N_CLK_M0_g N_4_c_20_n 2.42213e-19 $X=0.081 $Y=0.0675 $X2=0.054 $Y2=0.036
cc_8 CLK N_4_c_20_n 0.00198701f $X=0.081 $Y=0.1345 $X2=0.054 $Y2=0.036
cc_9 CLK N_4_c_22_n 9.57337e-19 $X=0.081 $Y=0.1345 $X2=0.054 $Y2=0.036
cc_10 CLK N_4_c_23_n 0.00123168f $X=0.081 $Y=0.1345 $X2=0.033 $Y2=0.153
cc_11 CLK N_4_c_24_n 0.0011151f $X=0.081 $Y=0.1345 $X2=0.175 $Y2=0.153
cc_12 CLK N_4_c_25_n 0.00362754f $X=0.081 $Y=0.1345 $X2=0.135 $Y2=0.135
cc_13 CLK N_9_c_302_n 2.03179e-19 $X=0.081 $Y=0.1345 $X2=0.693 $Y2=0.153
cc_14 N_4_c_15_n N_SE_c_143_n 2.02054e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 N_4_c_27_p N_SE_c_143_n 2.65253e-19 $X=0.434 $Y=0.153 $X2=0.081 $Y2=0.135
cc_16 N_4_M7_g N_SE_M5_g 2.88628e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_17 N_4_c_27_p N_SE_c_146_n 8.88734e-19 $X=0.434 $Y=0.153 $X2=0 $Y2=0
cc_18 N_4_c_27_p N_SE_c_147_n 0.00161831f $X=0.434 $Y=0.153 $X2=0 $Y2=0
cc_19 N_4_c_31_p N_SE_c_148_n 8.13099e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_20 N_4_c_27_p D 0.00130673f $X=0.434 $Y=0.153 $X2=0 $Y2=0
cc_21 N_4_c_31_p D 8.67096e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_22 N_4_c_27_p N_7_c_223_n 3.0124e-19 $X=0.434 $Y=0.153 $X2=0 $Y2=0
cc_23 N_4_c_27_p N_7_c_224_n 9.75625e-19 $X=0.434 $Y=0.153 $X2=0 $Y2=0
cc_24 N_4_c_31_p N_7_c_225_n 8.02031e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_25 N_4_c_27_p N_7_c_226_n 3.70293e-19 $X=0.434 $Y=0.153 $X2=0 $Y2=0
cc_26 N_4_M7_g N_SI_M6_g 0.00360681f $X=0.675 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_27 N_4_c_39_p N_SI_c_278_n 0.00113912f $X=0.693 $Y=0.135 $X2=0.081 $Y2=0.135
cc_28 N_4_M7_g SI 4.66746e-19 $X=0.675 $Y=0.0675 $X2=0.081 $Y2=0.1345
cc_29 N_4_c_31_p SI 8.81805e-19 $X=1.121 $Y=0.153 $X2=0.081 $Y2=0.1345
cc_30 N_4_c_39_p SI 2.88916e-19 $X=0.693 $Y=0.135 $X2=0.081 $Y2=0.1345
cc_31 N_4_c_43_p SI 0.00176948f $X=0.693 $Y=0.135 $X2=0.081 $Y2=0.1345
cc_32 N_4_M7_g N_9_M8_g 2.94371e-19 $X=0.675 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_33 N_4_c_45_p N_9_M8_g 0.00355599f $X=0.837 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_34 N_4_c_45_p N_9_c_305_n 0.00105615f $X=0.837 $Y=0.135 $X2=0.081 $Y2=0.135
cc_35 N_4_c_39_p N_9_c_305_n 4.70423e-19 $X=0.693 $Y=0.135 $X2=0.081 $Y2=0.135
cc_36 N_4_c_48_p N_9_M11_g 0.00365763f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_M12_g N_9_M11_g 0.00355599f $X=1.161 $Y=0.0675 $X2=0 $Y2=0
cc_38 N_4_c_48_p N_9_c_309_n 0.00104184f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_39 N_4_c_51_p N_9_c_309_n 9.99654e-19 $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_16_n N_9_c_311_n 2.58009e-19 $X=0.056 $Y=0.2025 $X2=0 $Y2=0
cc_41 N_4_c_24_n N_9_c_311_n 3.0124e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_42 N_4_c_25_n N_9_c_311_n 0.00114532f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_43 N_4_M1_g N_9_c_314_n 3.59377e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_4_c_20_n N_9_c_314_n 6.34683e-19 $X=0.054 $Y=0.036 $X2=0 $Y2=0
cc_45 N_4_c_25_n N_9_c_314_n 5.18786e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_22_n N_9_c_317_n 2.56213e-19 $X=0.054 $Y=0.036 $X2=0 $Y2=0
cc_47 N_4_c_24_n N_9_c_317_n 2.54113e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_48 N_4_c_60_p N_9_c_319_n 2.66501e-19 $X=0.054 $Y=0.234 $X2=0 $Y2=0
cc_49 N_4_c_24_n N_9_c_319_n 3.67164e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_50 N_4_c_27_p N_9_c_321_n 0.00116045f $X=0.434 $Y=0.153 $X2=0 $Y2=0
cc_51 N_4_c_25_n N_9_c_321_n 2.80227e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_52 N_4_c_31_p N_9_c_323_n 9.64586e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_53 N_4_c_65_p N_9_c_323_n 0.00403694f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_54 N_4_c_27_p N_9_c_325_n 0.0392002f $X=0.434 $Y=0.153 $X2=0 $Y2=0
cc_55 N_4_c_25_n N_9_c_325_n 3.53776e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_56 N_4_c_31_p N_9_c_327_n 0.0392002f $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_57 N_4_c_39_p N_9_c_328_n 2.05876e-19 $X=0.693 $Y=0.135 $X2=0 $Y2=0
cc_58 N_4_c_43_p N_9_c_328_n 2.46239e-19 $X=0.693 $Y=0.135 $X2=0 $Y2=0
cc_59 N_4_c_65_p N_9_c_328_n 0.00115955f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_60 N_4_c_72_p N_9_c_328_n 0.00124223f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_61 N_4_c_73_p N_9_c_328_n 3.53776e-19 $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_62 N_4_c_31_p N_9_c_333_n 0.00107275f $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_63 N_4_c_72_p N_9_c_333_n 0.00262191f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_64 N_4_c_73_p N_9_c_333_n 0.00260528f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_65 N_4_c_25_n N_9_c_336_n 0.00362295f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_66 N_4_c_45_p N_10_M9_g 0.00341068f $X=0.837 $Y=0.135 $X2=0.081 $Y2=0.135
cc_67 N_4_c_45_p N_10_c_381_n 0.00105614f $X=0.837 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_68 N_4_c_48_p N_10_c_382_n 0.00639681f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_69 N_4_c_31_p N_10_c_382_n 2.84796e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_70 N_4_c_72_p N_10_c_382_n 0.00138138f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_71 N_4_c_31_p N_10_c_385_n 7.48953e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_72 N_4_c_72_p N_10_c_385_n 0.00132074f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_73 N_4_c_31_p N_10_c_387_n 8.26567e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_74 N_4_c_65_p N_10_c_388_n 0.00384331f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_75 N_4_c_31_p N_10_c_389_n 4.07109e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_76 N_4_c_72_p N_10_c_389_n 0.00113688f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_77 N_4_c_45_p N_11_M10_g 2.13359e-19 $X=0.837 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_78 N_4_c_48_p N_11_M10_g 2.82885e-19 $X=1.053 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_79 N_4_c_48_p N_11_c_418_n 5.25211e-19 $X=1.053 $Y=0.135 $X2=0.081 $Y2=0.135
cc_80 N_4_c_31_p N_11_c_419_n 3.09707e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_81 N_4_c_39_p N_11_c_419_n 0.0010746f $X=0.693 $Y=0.135 $X2=0 $Y2=0
cc_82 N_4_c_43_p N_11_c_419_n 3.92611e-19 $X=0.693 $Y=0.135 $X2=0 $Y2=0
cc_83 N_4_c_31_p N_11_c_422_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_84 N_4_c_31_p N_11_c_423_n 8.09198e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_85 N_4_c_43_p N_11_c_423_n 0.00106879f $X=0.693 $Y=0.135 $X2=0 $Y2=0
cc_86 N_4_c_43_p N_11_c_425_n 0.00106879f $X=0.693 $Y=0.135 $X2=0 $Y2=0
cc_87 N_4_c_31_p N_11_c_426_n 3.46508e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_88 N_4_c_31_p N_11_c_427_n 2.42614e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_89 N_4_c_31_p N_11_c_428_n 4.07711e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_90 N_4_c_45_p N_11_c_429_n 3.51501e-19 $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_91 N_4_c_65_p N_11_c_429_n 5.11397e-19 $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_92 N_4_c_31_p N_11_c_431_n 7.80087e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_93 N_4_c_31_p N_11_c_432_n 0.00107683f $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_94 N_4_c_72_p N_11_c_432_n 4.32979e-19 $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_95 N_4_c_72_p N_11_c_434_n 4.15367e-19 $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_96 N_4_M12_g N_12_M13_g 0.00341068f $X=1.161 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_97 N_4_c_51_p N_12_c_476_n 9.22047e-19 $X=1.161 $Y=0.135 $X2=0.081 $Y2=0.135
cc_98 N_4_c_73_p N_12_c_477_n 0.00206054f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_99 N_4_c_73_p N_12_c_478_n 0.00206054f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_100 N_4_c_112_p N_12_c_479_n 3.54035e-19 $X=1.161 $Y=0.153 $X2=0 $Y2=0
cc_101 N_4_M12_g N_13_M14_g 2.13359e-19 $X=1.161 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_102 N_4_c_31_p N_13_c_507_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_103 N_4_c_72_p N_13_c_507_n 0.00130837f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_104 N_4_c_48_p N_13_c_509_n 2.20599e-19 $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_105 N_4_c_31_p N_13_c_509_n 5.75548e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_106 N_4_c_31_p N_13_c_511_n 3.8246e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_107 N_4_c_73_p N_13_c_512_n 0.00102938f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_108 N_4_c_120_p N_13_c_513_n 2.51466e-19 $X=1.141 $Y=0.153 $X2=0 $Y2=0
cc_109 N_4_M12_g N_13_c_514_n 3.57114e-19 $X=1.161 $Y=0.0675 $X2=0 $Y2=0
cc_110 N_4_c_73_p N_13_c_514_n 5.22021e-19 $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_111 N_4_c_27_p N_15_c_573_n 2.98103e-19 $X=0.434 $Y=0.153 $X2=0.081 $Y2=0.135
cc_112 N_4_c_31_p N_15_c_574_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_113 N_4_c_31_p N_15_c_575_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0.081 $Y2=0.135
cc_114 N_4_c_27_p N_15_c_576_n 3.08895e-19 $X=0.434 $Y=0.153 $X2=0 $Y2=0
cc_115 N_4_c_31_p N_15_c_577_n 4.72621e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_116 N_4_c_31_p N_15_c_578_n 4.8224e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_117 N_4_c_31_p N_15_c_579_n 3.65983e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_118 N_4_c_31_p N_15_c_580_n 4.66683e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_119 N_4_c_31_p N_16_c_605_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0.081 $Y2=0.135
cc_120 N_4_M7_g N_16_c_606_n 4.39425e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_121 N_4_c_31_p N_16_c_606_n 3.48349e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_122 N_4_c_43_p N_16_c_608_n 5.53288e-19 $X=0.693 $Y=0.135 $X2=0 $Y2=0
cc_123 N_4_c_31_p N_16_c_609_n 6.02073e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_124 N_4_c_45_p N_18_c_650_n 0.00639681f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_125 N_4_c_31_p N_18_c_650_n 3.30527e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_126 N_4_c_65_p N_18_c_650_n 0.00372445f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_127 N_4_M12_g N_19_c_661_n 0.00382563f $X=1.161 $Y=0.0675 $X2=0 $Y2=0
cc_128 N_4_c_51_p N_19_c_661_n 0.0019701f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_129 N_4_c_120_p N_19_c_661_n 4.50035e-19 $X=1.141 $Y=0.153 $X2=0 $Y2=0
cc_130 N_4_c_73_p N_19_c_661_n 0.00376163f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_131 N_SE_M5_g N_D_M3_g 2.13359e-19 $X=0.567 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_132 N_SE_c_143_n N_D_c_202_n 2.39808e-19 $X=0.297 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_133 N_SE_c_147_n D 3.54801e-19 $X=0.567 $Y=0.081 $X2=1.053 $Y2=0.2025
cc_134 N_SE_M5_g N_7_M4_g 0.00304756f $X=0.567 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_135 N_SE_c_153_p N_7_c_228_n 0.00105615f $X=0.567 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_136 N_SE_c_154_p N_7_c_229_n 6.84024e-19 $X=0.243 $Y=0.081 $X2=0 $Y2=0
cc_137 N_SE_c_147_n N_7_c_230_n 6.55402e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_138 SE N_7_c_231_n 4.48296e-19 $X=0.278 $Y=0.1345 $X2=1.053 $Y2=0.2025
cc_139 N_SE_c_146_n N_7_c_224_n 6.16983e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_140 N_SE_c_147_n N_7_c_233_n 9.88868e-19 $X=0.567 $Y=0.081 $X2=1.161
+ $Y2=0.0675
cc_141 N_SE_c_159_p N_7_c_233_n 0.00105704f $X=0.567 $Y=0.081 $X2=1.161
+ $Y2=0.0675
cc_142 N_SE_c_147_n N_7_c_235_n 4.38038e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_143 N_SE_c_147_n N_7_c_236_n 0.00100123f $X=0.567 $Y=0.081 $X2=1.161
+ $Y2=0.135
cc_144 N_SE_c_147_n N_7_c_237_n 0.00123902f $X=0.567 $Y=0.081 $X2=1.161
+ $Y2=0.135
cc_145 N_SE_c_147_n N_7_c_238_n 4.81197e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_146 N_SE_c_148_n N_7_c_225_n 0.00105704f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_147 N_SE_c_147_n N_7_c_240_n 5.77999e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_148 N_SE_c_166_p N_7_c_240_n 0.00115045f $X=0.567 $Y=0.106 $X2=0 $Y2=0
cc_149 N_SE_c_167_p N_7_c_242_n 0.00105704f $X=0.567 $Y=0.1205 $X2=0.071
+ $Y2=0.2025
cc_150 N_SE_c_147_n N_7_c_243_n 3.53821e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_151 N_SE_c_154_p N_7_c_244_n 6.58915e-19 $X=0.243 $Y=0.081 $X2=0.018
+ $Y2=0.063
cc_152 N_SE_c_147_n N_7_c_244_n 4.3742e-19 $X=0.567 $Y=0.081 $X2=0.018 $Y2=0.063
cc_153 N_SE_c_146_n N_7_c_226_n 6.58915e-19 $X=0.243 $Y=0.135 $X2=0.054
+ $Y2=0.036
cc_154 N_SE_c_147_n N_7_c_247_n 3.89571e-19 $X=0.567 $Y=0.081 $X2=0.0505
+ $Y2=0.036
cc_155 N_SE_M5_g N_SI_M6_g 0.00348334f $X=0.567 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_156 N_SE_c_153_p N_SI_c_278_n 0.00105615f $X=0.567 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_157 N_SE_c_159_p SI 7.03144e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_158 N_SE_c_148_n SI 0.00123983f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_159 N_SE_c_166_p SI 5.30073e-19 $X=0.567 $Y=0.106 $X2=0 $Y2=0
cc_160 N_SE_c_167_p SI 0.00123983f $X=0.567 $Y=0.1205 $X2=0 $Y2=0
cc_161 N_SE_c_154_p N_9_c_337_n 0.00211968f $X=0.243 $Y=0.081 $X2=1.161
+ $Y2=0.0675
cc_162 N_SE_c_146_n N_9_c_338_n 0.00211968f $X=0.243 $Y=0.135 $X2=0.056
+ $Y2=0.2025
cc_163 N_SE_c_146_n N_9_c_321_n 0.00211968f $X=0.243 $Y=0.135 $X2=0.018
+ $Y2=0.1035
cc_164 N_SE_c_143_n N_9_c_327_n 2.61615e-19 $X=0.297 $Y=0.135 $X2=0.054
+ $Y2=0.036
cc_165 N_SE_c_154_p N_9_c_327_n 0.00115508f $X=0.243 $Y=0.081 $X2=0.054
+ $Y2=0.036
cc_166 N_SE_c_147_n N_9_c_327_n 0.0291996f $X=0.567 $Y=0.081 $X2=0.054 $Y2=0.036
cc_167 N_SE_c_148_n N_9_c_327_n 3.29785e-19 $X=0.567 $Y=0.135 $X2=0.054
+ $Y2=0.036
cc_168 N_SE_c_166_p N_9_c_327_n 2.46239e-19 $X=0.567 $Y=0.106 $X2=0.054
+ $Y2=0.036
cc_169 N_SE_c_167_p N_9_c_327_n 5.96604e-19 $X=0.567 $Y=0.1205 $X2=0.054
+ $Y2=0.036
cc_170 N_SE_c_159_p N_9_c_328_n 3.45641e-19 $X=0.567 $Y=0.081 $X2=0.054
+ $Y2=0.036
cc_171 N_SE_c_154_p N_9_c_347_n 0.00211968f $X=0.243 $Y=0.081 $X2=0.693
+ $Y2=0.153
cc_172 N_SE_c_147_n N_9_c_302_n 3.51588e-19 $X=0.567 $Y=0.081 $X2=0.693
+ $Y2=0.153
cc_173 N_SE_c_146_n N_9_c_349_n 0.00211968f $X=0.243 $Y=0.135 $X2=0.175
+ $Y2=0.153
cc_174 VSS N_SE_c_147_n 2.01433e-19 $X=0.567 $Y=0.081 $X2=0.675 $Y2=0.135
cc_175 VSS N_SE_c_147_n 4.83825e-19 $X=0.567 $Y=0.081 $X2=0.837 $Y2=0.2025
cc_176 VSS N_SE_M5_g 2.34002e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_177 VSS N_SE_c_159_p 0.00426739f $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_178 N_SE_M5_g N_15_c_581_n 3.61002e-19 $X=0.567 $Y=0.0675 $X2=0.071
+ $Y2=0.0675
cc_179 N_SE_c_148_n N_15_c_581_n 0.00117826f $X=0.567 $Y=0.135 $X2=0.071
+ $Y2=0.0675
cc_180 VSS N_SE_c_159_p 3.06453e-19 $X=0.567 $Y=0.081 $X2=0.135 $Y2=0.0675
cc_181 N_D_M3_g N_7_M4_g 0.00304756f $X=0.459 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_182 N_D_c_202_n N_7_c_228_n 0.00105595f $X=0.459 $Y=0.135 $X2=0.135 $Y2=0.135
cc_183 D N_7_c_250_n 0.00251305f $X=0.459 $Y=0.1345 $X2=1.053 $Y2=0.135
cc_184 D N_7_c_251_n 0.00251305f $X=0.459 $Y=0.1345 $X2=1.053 $Y2=0.2025
cc_185 D N_7_c_231_n 0.00251305f $X=0.459 $Y=0.1345 $X2=1.053 $Y2=0.2025
cc_186 D N_7_c_224_n 0.00251305f $X=0.459 $Y=0.1345 $X2=0 $Y2=0
cc_187 D N_7_c_236_n 0.00388774f $X=0.459 $Y=0.1345 $X2=1.161 $Y2=0.135
cc_188 N_D_M3_g N_7_c_237_n 2.16728e-19 $X=0.459 $Y=0.0675 $X2=1.161 $Y2=0.135
cc_189 D N_7_c_237_n 0.00388774f $X=0.459 $Y=0.1345 $X2=1.161 $Y2=0.135
cc_190 D N_7_c_225_n 0.00141867f $X=0.459 $Y=0.1345 $X2=0 $Y2=0
cc_191 D N_7_c_242_n 0.00141867f $X=0.459 $Y=0.1345 $X2=0.071 $Y2=0.2025
cc_192 D N_7_c_259_n 0.00251305f $X=0.459 $Y=0.1345 $X2=0.054 $Y2=0.036
cc_193 D N_9_c_327_n 0.0013631f $X=0.459 $Y=0.1345 $X2=0.054 $Y2=0.036
cc_194 VSS D 0.00172965f $X=0.459 $Y=0.1345 $X2=0.675 $Y2=0.135
cc_195 VSS N_D_M3_g 2.37298e-19 $X=0.459 $Y=0.0675 $X2=0.837 $Y2=0.2025
cc_196 D N_15_M22_s 3.13248e-19 $X=0.459 $Y=0.1345 $X2=0.135 $Y2=0.0675
cc_197 D N_15_c_573_n 0.00310236f $X=0.459 $Y=0.1345 $X2=0.135 $Y2=0.135
cc_198 D N_15_c_576_n 0.00415606f $X=0.459 $Y=0.1345 $X2=0 $Y2=0
cc_199 D N_15_c_586_n 0.00115405f $X=0.459 $Y=0.1345 $X2=1.053 $Y2=0.2025
cc_200 N_7_M4_g N_SI_M6_g 2.48122e-19 $X=0.513 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_201 N_7_c_223_n N_9_c_311_n 2.28803e-19 $X=0.322 $Y=0.2025 $X2=1.053
+ $Y2=0.2025
cc_202 N_7_c_251_n N_9_c_327_n 9.86944e-19 $X=0.351 $Y=0.126 $X2=0.054 $Y2=0.036
cc_203 N_7_c_225_n N_9_c_327_n 4.55831e-19 $X=0.513 $Y=0.135 $X2=0.054 $Y2=0.036
cc_204 N_7_c_242_n N_9_c_327_n 4.65024e-19 $X=0.513 $Y=0.117 $X2=0.054 $Y2=0.036
cc_205 VSS N_7_c_237_n 3.22316e-19 $X=0.468 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_206 VSS N_7_c_229_n 2.68628e-19 $X=0.351 $Y=0.063 $X2=0.675 $Y2=0.135
cc_207 VSS N_7_c_230_n 2.08206e-19 $X=0.351 $Y=0.099 $X2=0.675 $Y2=0.135
cc_208 VSS N_7_c_237_n 0.00291153f $X=0.468 $Y=0.072 $X2=0.675 $Y2=0.135
cc_209 VSS N_7_c_240_n 2.08206e-19 $X=0.513 $Y=0.099 $X2=0.675 $Y2=0.135
cc_210 VSS N_7_c_243_n 0.00133246f $X=0.324 $Y=0.036 $X2=0.675 $Y2=0.135
cc_211 VSS N_7_M4_g 2.34002e-19 $X=0.513 $Y=0.0675 $X2=0.837 $Y2=0.2025
cc_212 VSS N_7_c_237_n 0.00904478f $X=0.468 $Y=0.072 $X2=0.837 $Y2=0.2025
cc_213 VSS N_7_c_273_p 6.34674e-19 $X=0.351 $Y=0.036 $X2=0.837 $Y2=0.2025
cc_214 N_7_c_223_n N_15_c_573_n 0.00134514f $X=0.322 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_215 N_7_M4_g N_15_c_588_n 3.50974e-19 $X=0.513 $Y=0.0675 $X2=1.161 $Y2=0.0675
cc_216 N_7_c_225_n N_15_c_588_n 0.00116301f $X=0.513 $Y=0.135 $X2=1.161
+ $Y2=0.0675
cc_217 SI N_9_c_328_n 0.00204819f $X=0.621 $Y=0.1345 $X2=0.054 $Y2=0.036
cc_218 SI N_11_c_419_n 0.0083394f $X=0.621 $Y=0.1345 $X2=0 $Y2=0
cc_219 SI N_11_c_436_n 0.00227527f $X=0.621 $Y=0.1345 $X2=0 $Y2=0
cc_220 VSS SI 0.00196285f $X=0.621 $Y=0.1345 $X2=0.837 $Y2=0.135
cc_221 VSS SI 0.00389367f $X=0.621 $Y=0.1345 $X2=0 $Y2=0
cc_222 VSS N_SI_M6_g 3.5204e-19 $X=0.621 $Y=0.0675 $X2=1.053 $Y2=0.135
cc_223 VSS SI 6.77952e-19 $X=0.621 $Y=0.1345 $X2=1.053 $Y2=0.135
cc_224 VSS SI 0.0010238f $X=0.621 $Y=0.1345 $X2=0 $Y2=0
cc_225 SI N_15_c_579_n 4.77922e-19 $X=0.621 $Y=0.1345 $X2=1.161 $Y2=0.135
cc_226 N_SI_M6_g N_15_c_591_n 2.75159e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_227 SI N_15_c_591_n 0.00116629f $X=0.621 $Y=0.1345 $X2=0 $Y2=0
cc_228 N_SI_M6_g N_16_c_610_n 2.38237e-19 $X=0.621 $Y=0.0675 $X2=0.837
+ $Y2=0.2025
cc_229 N_9_M8_g N_10_M9_g 2.82885e-19 $X=0.783 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_230 N_9_c_328_n N_10_c_382_n 0.00134228f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_231 N_9_c_333_n N_10_c_382_n 0.00127195f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_232 N_9_c_328_n N_10_c_387_n 3.31762e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_233 N_9_c_328_n N_10_c_395_n 5.67404e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_234 N_9_c_328_n N_10_c_396_n 3.4734e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_235 N_9_c_328_n N_10_c_397_n 4.8206e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_236 N_9_c_328_n N_10_c_389_n 4.09721e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_237 N_9_c_323_n N_11_c_419_n 4.91424e-19 $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_238 N_9_c_328_n N_11_c_419_n 8.86983e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_239 N_9_c_323_n N_11_c_436_n 0.00811029f $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_240 N_9_c_328_n N_11_c_436_n 5.82789e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_241 N_9_c_323_n N_11_c_423_n 2.60223e-19 $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_242 N_9_c_328_n N_11_c_423_n 3.09845e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_243 N_9_M8_g N_11_c_443_n 3.61002e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_244 N_9_c_323_n N_11_c_443_n 0.001177f $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_245 N_9_c_328_n N_11_c_432_n 9.67845e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_246 N_9_M11_g N_12_M13_g 2.82885e-19 $X=1.107 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_247 N_9_M11_g N_13_c_516_n 3.47081e-19 $X=1.107 $Y=0.0675 $X2=0 $Y2=0
cc_248 N_9_c_333_n N_13_c_516_n 4.94366e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_249 N_9_c_333_n N_13_c_513_n 0.00130997f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_250 VSS N_9_c_328_n 2.05877e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_251 N_9_c_323_n N_18_c_650_n 0.00102036f $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_252 N_9_c_328_n N_18_c_650_n 0.00124591f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_253 N_10_M9_g N_11_M10_g 0.00268443f $X=0.891 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_254 N_10_c_400_p N_11_M10_g 3.61002e-19 $X=0.954 $Y=0.072 $X2=0.135
+ $Y2=0.0675
cc_255 N_10_c_381_n N_11_c_418_n 0.00105598f $X=0.891 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_256 N_10_M9_g N_11_c_449_n 3.56998e-19 $X=0.891 $Y=0.0675 $X2=0.027 $Y2=0.036
cc_257 N_10_c_387_n N_11_c_449_n 4.80589e-19 $X=0.891 $Y=0.135 $X2=0.027
+ $Y2=0.036
cc_258 N_10_c_385_n N_11_c_432_n 0.00242354f $X=1.028 $Y=0.2025 $X2=0.054
+ $Y2=0.036
cc_259 N_10_c_395_n N_11_c_432_n 0.0021413f $X=0.891 $Y=0.1205 $X2=0.054
+ $Y2=0.036
cc_260 N_10_c_400_p N_11_c_432_n 0.00118287f $X=0.954 $Y=0.072 $X2=0.054
+ $Y2=0.036
cc_261 N_10_c_389_n N_11_c_432_n 0.00115834f $X=0.999 $Y=0.162 $X2=0.054
+ $Y2=0.036
cc_262 N_10_c_382_n N_13_c_507_n 0.00122411f $X=1.082 $Y=0.0675 $X2=0.018
+ $Y2=0.2125
cc_263 N_10_c_385_n N_13_c_507_n 0.00270924f $X=1.028 $Y=0.2025 $X2=0.018
+ $Y2=0.2125
cc_264 N_10_c_385_n N_13_c_509_n 5.74875e-19 $X=1.028 $Y=0.2025 $X2=0.054
+ $Y2=0.036
cc_265 N_10_c_382_n N_13_c_522_n 3.1278e-19 $X=1.082 $Y=0.0675 $X2=0 $Y2=0
cc_266 N_10_c_382_n N_13_c_513_n 0.00278091f $X=1.082 $Y=0.0675 $X2=0.033
+ $Y2=0.153
cc_267 N_10_c_382_n N_18_c_650_n 3.26365e-19 $X=1.082 $Y=0.0675 $X2=0.675
+ $Y2=0.0675
cc_268 N_10_c_388_n N_18_c_650_n 0.00127189f $X=0.9 $Y=0.072 $X2=0.675
+ $Y2=0.0675
cc_269 N_10_c_385_n N_19_c_661_n 3.11986e-19 $X=1.028 $Y=0.2025 $X2=0.675
+ $Y2=0.0675
cc_270 VSS N_11_c_419_n 2.62157e-19 $X=0.758 $Y=0.0675 $X2=0.837 $Y2=0.135
cc_271 VSS N_11_c_419_n 0.004062f $X=0.758 $Y=0.0675 $X2=0 $Y2=0
cc_272 N_11_c_457_p N_15_c_575_n 2.93059e-19 $X=0.747 $Y=0.178 $X2=0 $Y2=0
cc_273 N_11_c_458_p N_15_c_579_n 6.37567e-19 $X=0.756 $Y=0.198 $X2=1.161
+ $Y2=0.135
cc_274 N_11_c_419_n N_16_c_611_n 0.00114234f $X=0.758 $Y=0.0675 $X2=0.675
+ $Y2=0.0675
cc_275 N_11_c_422_n N_16_c_611_n 0.00380633f $X=0.81 $Y=0.2025 $X2=0.675
+ $Y2=0.0675
cc_276 N_11_c_461_p N_16_c_611_n 3.87816e-19 $X=0.747 $Y=0.189 $X2=0.675
+ $Y2=0.0675
cc_277 N_11_c_423_n N_16_c_611_n 4.18661e-19 $X=0.747 $Y=0.164 $X2=0.675
+ $Y2=0.0675
cc_278 N_11_c_457_p N_16_c_611_n 4.06284e-19 $X=0.747 $Y=0.178 $X2=0.675
+ $Y2=0.0675
cc_279 N_11_c_458_p N_16_c_611_n 6.70593e-19 $X=0.756 $Y=0.198 $X2=0.675
+ $Y2=0.0675
cc_280 N_11_c_427_n N_16_c_611_n 7.05929e-19 $X=0.767 $Y=0.198 $X2=0.675
+ $Y2=0.0675
cc_281 N_11_c_466_p N_16_c_611_n 4.19603e-19 $X=0.77 $Y=0.198 $X2=0.675
+ $Y2=0.0675
cc_282 N_11_c_422_n N_16_c_619_n 2.42261e-19 $X=0.81 $Y=0.2025 $X2=0.837
+ $Y2=0.135
cc_283 N_11_c_427_n N_16_c_619_n 0.00137625f $X=0.767 $Y=0.198 $X2=0.837
+ $Y2=0.135
cc_284 N_11_c_469_p N_16_c_619_n 9.77254e-19 $X=0.819 $Y=0.234 $X2=0.837
+ $Y2=0.135
cc_285 N_11_c_458_p N_16_c_622_n 0.00137625f $X=0.756 $Y=0.198 $X2=0 $Y2=0
cc_286 N_11_c_419_n N_18_c_650_n 0.00479956f $X=0.758 $Y=0.0675 $X2=0.675
+ $Y2=0.0675
cc_287 N_11_c_422_n N_18_c_650_n 0.00138279f $X=0.81 $Y=0.2025 $X2=0.675
+ $Y2=0.0675
cc_288 N_11_c_431_n N_18_c_650_n 4.23207e-19 $X=0.882 $Y=0.234 $X2=0.675
+ $Y2=0.0675
cc_289 N_11_c_431_n N_23_M28_s 5.02871e-19 $X=0.882 $Y=0.234 $X2=0.135
+ $Y2=0.0675
cc_290 N_12_M13_g N_13_M14_g 0.00268443f $X=1.215 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_291 N_12_c_482_p N_13_M14_g 3.29607e-19 $X=1.283 $Y=0.191 $X2=0.135
+ $Y2=0.0675
cc_292 N_12_c_476_n N_13_c_526_n 0.00108446f $X=1.215 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_293 N_12_M13_g N_13_c_527_n 2.64276e-19 $X=1.215 $Y=0.0675 $X2=0.054
+ $Y2=0.234
cc_294 N_12_c_485_p N_13_c_527_n 0.00321328f $X=1.294 $Y=0.2025 $X2=0.054
+ $Y2=0.234
cc_295 N_12_c_486_p N_13_c_527_n 0.00838811f $X=1.224 $Y=0.191 $X2=0.054
+ $Y2=0.234
cc_296 N_12_c_487_p N_13_c_513_n 2.02397e-19 $X=1.294 $Y=0.0675 $X2=0.033
+ $Y2=0.153
cc_297 N_12_M13_g N_13_c_531_n 3.57119e-19 $X=1.215 $Y=0.0675 $X2=0.693
+ $Y2=0.153
cc_298 N_12_c_478_n N_13_c_531_n 5.37372e-19 $X=1.215 $Y=0.135 $X2=0.693
+ $Y2=0.153
cc_299 N_12_c_487_p N_13_c_533_n 0.00115323f $X=1.294 $Y=0.0675 $X2=0.175
+ $Y2=0.153
cc_300 N_12_c_491_p N_13_c_534_n 9.36593e-19 $X=1.314 $Y=0.09 $X2=0.837
+ $Y2=0.153
cc_301 N_12_c_492_p N_13_c_535_n 7.6566e-19 $X=1.323 $Y=0.126 $X2=0.837
+ $Y2=0.153
cc_302 N_12_c_478_n N_13_c_536_n 0.0030621f $X=1.215 $Y=0.135 $X2=1.053
+ $Y2=0.153
cc_303 N_12_c_487_p N_13_c_537_n 6.1907e-19 $X=1.294 $Y=0.0675 $X2=1.161
+ $Y2=0.153
cc_304 N_12_c_487_p N_13_c_538_n 0.003475f $X=1.294 $Y=0.0675 $X2=1.161
+ $Y2=0.153
cc_305 N_12_c_491_p N_13_c_538_n 0.00207793f $X=1.314 $Y=0.09 $X2=1.161
+ $Y2=0.153
cc_306 N_12_c_492_p N_13_c_540_n 0.00149664f $X=1.323 $Y=0.126 $X2=0 $Y2=0
cc_307 N_12_c_487_p N_13_c_541_n 3.63761e-19 $X=1.294 $Y=0.0675 $X2=0 $Y2=0
cc_308 N_12_c_499_p N_13_c_542_n 0.00149664f $X=1.323 $Y=0.09 $X2=0.135
+ $Y2=0.135
cc_309 N_12_c_500_p N_13_c_543_n 0.00149664f $X=1.323 $Y=0.182 $X2=0 $Y2=0
cc_310 N_12_c_501_p N_13_c_544_n 9.53904e-19 $X=1.323 $Y=0.144 $X2=0 $Y2=0
cc_311 N_12_c_482_p N_13_c_545_n 0.00190954f $X=1.283 $Y=0.191 $X2=0 $Y2=0
cc_312 N_12_c_501_p N_13_c_546_n 0.00149664f $X=1.323 $Y=0.144 $X2=0 $Y2=0
cc_313 N_12_c_485_p N_19_c_661_n 2.83378e-19 $X=1.294 $Y=0.2025 $X2=0.675
+ $Y2=0.0675
cc_314 N_12_c_479_n N_19_c_661_n 0.00102083f $X=1.215 $Y=0.163 $X2=0.675
+ $Y2=0.0675
cc_315 N_13_c_547_p N_QN_M16_d 3.8044e-19 $X=1.593 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_316 N_13_c_547_p N_QN_M18_d 3.80663e-19 $X=1.593 $Y=0.135 $X2=0.135
+ $Y2=0.2025
cc_317 N_13_c_547_p N_QN_M35_d 3.8044e-19 $X=1.593 $Y=0.135 $X2=0 $Y2=0
cc_318 N_13_c_547_p N_QN_c_634_n 7.78051e-19 $X=1.593 $Y=0.135 $X2=0.837
+ $Y2=0.135
cc_319 N_13_c_547_p N_QN_M37_d 3.80663e-19 $X=1.593 $Y=0.135 $X2=0.837 $Y2=0.135
cc_320 N_13_c_547_p N_QN_c_636_n 8.00061e-19 $X=1.593 $Y=0.135 $X2=0 $Y2=0
cc_321 N_13_M16_g N_QN_c_637_n 4.59284e-19 $X=1.485 $Y=0.0675 $X2=1.053
+ $Y2=0.135
cc_322 N_13_M17_g N_QN_c_637_n 4.59284e-19 $X=1.539 $Y=0.0675 $X2=1.053
+ $Y2=0.135
cc_323 N_13_M18_g N_QN_c_637_n 4.59284e-19 $X=1.593 $Y=0.0675 $X2=1.053
+ $Y2=0.135
cc_324 N_13_c_547_p N_QN_c_640_n 0.00187443f $X=1.593 $Y=0.135 $X2=0 $Y2=0
cc_325 N_13_c_557_p N_QN_c_640_n 4.23911e-19 $X=1.368 $Y=0.036 $X2=0 $Y2=0
cc_326 N_13_c_547_p N_QN_c_642_n 7.78051e-19 $X=1.593 $Y=0.135 $X2=1.053
+ $Y2=0.2025
cc_327 N_13_c_547_p N_QN_c_643_n 8.00061e-19 $X=1.593 $Y=0.135 $X2=1.161
+ $Y2=0.135
cc_328 N_13_M16_g N_QN_c_644_n 4.59284e-19 $X=1.485 $Y=0.0675 $X2=1.161
+ $Y2=0.135
cc_329 N_13_M17_g N_QN_c_644_n 4.59284e-19 $X=1.539 $Y=0.0675 $X2=1.161
+ $Y2=0.135
cc_330 N_13_M18_g N_QN_c_644_n 4.59284e-19 $X=1.593 $Y=0.0675 $X2=1.161
+ $Y2=0.135
cc_331 N_13_c_547_p N_QN_c_647_n 0.00187443f $X=1.593 $Y=0.135 $X2=0.071
+ $Y2=0.0675
cc_332 N_13_c_564_p N_QN_c_647_n 4.26942e-19 $X=1.368 $Y=0.234 $X2=0.071
+ $Y2=0.0675
cc_333 N_13_c_547_p N_QN_c_649_n 5.09179e-19 $X=1.593 $Y=0.135 $X2=0.018
+ $Y2=0.063
cc_334 N_13_c_507_n N_19_c_661_n 0.00412407f $X=1.08 $Y=0.2025 $X2=0.675
+ $Y2=0.0675
cc_335 N_13_c_511_n N_19_c_661_n 0.00284013f $X=1.152 $Y=0.234 $X2=0.675
+ $Y2=0.0675
cc_336 N_13_c_512_n N_19_c_661_n 0.00111255f $X=1.17 $Y=0.234 $X2=0.675
+ $Y2=0.0675
cc_337 N_13_c_569_p N_19_c_661_n 0.00302676f $X=1.206 $Y=0.234 $X2=0.675
+ $Y2=0.0675
cc_338 N_13_c_513_n N_19_c_661_n 0.00114658f $X=1.134 $Y=0.036 $X2=0.675
+ $Y2=0.0675
cc_339 N_13_c_571_p N_19_c_661_n 2.10553e-19 $X=1.206 $Y=0.036 $X2=0.675
+ $Y2=0.0675
cc_340 N_13_c_571_p N_22_M13_s 4.40115e-19 $X=1.206 $Y=0.036 $X2=0.135
+ $Y2=0.0675
cc_341 VSS N_15_c_573_n 0.0012476f $X=0.432 $Y=0.036 $X2=0.135 $Y2=0.135
cc_342 VSS N_15_c_575_n 0.0012783f $X=0.648 $Y=0.036 $X2=0 $Y2=0
cc_343 VSS N_18_c_650_n 3.09059e-19 $X=0.648 $Y=0.036 $X2=0.675 $Y2=0.0675
cc_344 N_15_c_574_n N_16_c_605_n 0.00323532f $X=0.54 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_345 N_15_c_575_n N_16_c_605_n 0.00352176f $X=0.646 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_346 N_15_c_599_p N_16_c_605_n 0.00145268f $X=0.599 $Y=0.198 $X2=0.135
+ $Y2=0.135
cc_347 N_15_c_600_p N_16_c_605_n 8.58362e-19 $X=0.612 $Y=0.198 $X2=0.135
+ $Y2=0.135
cc_348 N_15_c_575_n N_16_c_611_n 0.00122215f $X=0.646 $Y=0.2025 $X2=0.675
+ $Y2=0.0675
cc_349 N_15_c_574_n N_16_c_610_n 5.00576e-19 $X=0.54 $Y=0.2025 $X2=0.837
+ $Y2=0.2025
cc_350 N_15_c_575_n N_16_c_610_n 0.0030897f $X=0.646 $Y=0.2025 $X2=0.837
+ $Y2=0.2025
cc_351 N_15_c_599_p N_16_c_610_n 0.00701208f $X=0.599 $Y=0.198 $X2=0.837
+ $Y2=0.2025

* END of "./SDFHx4_ASAP7_75t_SRAM.pex.sp.SDFHX4_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: SDFLx1_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 13:04:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "SDFLx1_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./SDFLx1_ASAP7_75t_SRAM.pex.sp.pex"
* File: SDFLx1_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 13:04:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_SDFLX1_ASAP7_75T_SRAM%CLK 2 5 7 11 16 VSS
c12 11 VSS 0.00713456f $X=0.081 $Y=0.135
c13 5 VSS 0.00188964f $X=0.081 $Y=0.135
c14 2 VSS 0.0628473f $X=0.081 $Y=0.054
r15 11 16 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.15
r16 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%4 2 5 7 10 13 16 19 22 25 28 31 45 48 50 57 58 65
+ 72 79 83 86 90 97 100 101 102 104 123 VSS
c121 134 VSS 7.0154e-20 $X=0.03 $Y=0.189
c122 133 VSS 5.9624e-19 $X=0.027 $Y=0.189
c123 123 VSS 6.49238e-19 $X=0.729 $Y=0.18
c124 104 VSS 0.00976003f $X=0.729 $Y=0.189
c125 102 VSS 0.00542037f $X=0.371 $Y=0.189
c126 101 VSS 0.00609885f $X=0.175 $Y=0.189
c127 100 VSS 0.0013748f $X=0.567 $Y=0.189
c128 97 VSS 0.00291011f $X=0.135 $Y=0.189
c129 93 VSS 5.52785e-19 $X=0.033 $Y=0.189
c130 90 VSS 9.61695e-20 $X=0.567 $Y=0.18
c131 86 VSS 5.76385e-19 $X=0.567 $Y=0.135
c132 83 VSS 1.05495e-19 $X=0.135 $Y=0.18
c133 79 VSS 6.50523e-19 $X=0.135 $Y=0.135
c134 75 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c135 74 VSS 0.00169428f $X=0.047 $Y=0.234
c136 72 VSS 0.0024557f $X=0.054 $Y=0.234
c137 70 VSS 0.00306385f $X=0.027 $Y=0.234
c138 68 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c139 67 VSS 0.00205521f $X=0.047 $Y=0.036
c140 65 VSS 0.00239525f $X=0.054 $Y=0.036
c141 63 VSS 0.00305101f $X=0.027 $Y=0.036
c142 62 VSS 3.84318e-19 $X=0.018 $Y=0.216
c143 61 VSS 3.30259e-19 $X=0.018 $Y=0.207
c144 60 VSS 3.64183e-19 $X=0.018 $Y=0.225
c145 58 VSS 0.0039492f $X=0.018 $Y=0.164
c146 57 VSS 0.00142827f $X=0.018 $Y=0.081
c147 56 VSS 8.21418e-19 $X=0.018 $Y=0.18
c148 53 VSS 0.00514186f $X=0.056 $Y=0.216
c149 50 VSS 2.98509e-19 $X=0.071 $Y=0.216
c150 48 VSS 0.00458629f $X=0.056 $Y=0.054
c151 45 VSS 2.98509e-19 $X=0.071 $Y=0.054
c152 28 VSS 0.108004f $X=0.945 $Y=0.178
c153 25 VSS 1.08457e-19 $X=0.837 $Y=0.178
c154 22 VSS 0.060017f $X=0.837 $Y=0.0405
c155 19 VSS 2.24613e-19 $X=0.675 $Y=0.178
c156 16 VSS 0.0602569f $X=0.675 $Y=0.0405
c157 10 VSS 0.0660345f $X=0.567 $Y=0.1355
c158 5 VSS 0.00179729f $X=0.135 $Y=0.135
c159 2 VSS 0.0627664f $X=0.135 $Y=0.054
r160 133 134 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.03 $Y2=0.189
r161 130 133 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.027 $Y2=0.189
r162 122 123 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.729 $Y=0.18
+ $X2=0.729 $Y2=0.18
r163 104 123 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.729 $Y=0.189 $X2=0.729
+ $Y2=0.189
r164 101 102 13.3086 $w=1.8e-08 $l=1.96e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.175 $Y=0.189 $X2=0.371 $Y2=0.189
r165 99 104 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.729 $Y2=0.189
r166 99 102 13.3086 $w=1.8e-08 $l=1.96e-07 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.371 $Y2=0.189
r167 99 100 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.567 $Y=0.189 $X2=0.567
+ $Y2=0.189
r168 96 101 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.175 $Y2=0.189
r169 96 97 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.135 $Y=0.189 $X2=0.135
+ $Y2=0.189
r170 93 134 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.03 $Y2=0.189
r171 92 96 6.92593 $w=1.8e-08 $l=1.02e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.135 $Y2=0.189
r172 92 93 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.189 $X2=0.033
+ $Y2=0.189
r173 90 100 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.18 $X2=0.567 $Y2=0.189
r174 89 90 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.171 $X2=0.567 $Y2=0.18
r175 86 89 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.171
r176 83 97 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.18 $X2=0.135 $Y2=0.189
r177 82 83 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.164 $X2=0.135 $Y2=0.18
r178 79 82 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.164
r179 74 75 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r180 72 75 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r181 70 74 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r182 67 68 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r183 65 68 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r184 63 67 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r185 61 62 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.207 $X2=0.018 $Y2=0.216
r186 60 70 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r187 60 62 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.216
r188 59 130 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.189
r189 59 61 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.207
r190 57 58 5.6358 $w=1.8e-08 $l=8.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.164
r191 56 130 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.189
r192 56 58 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.164
r193 55 63 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r194 55 57 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r195 53 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r196 50 53 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r197 48 65 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r198 45 48 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r199 28 31 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.178 $X2=0.945 $Y2=0.2295
r200 25 28 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08 $X=0.837
+ $Y=0.178 $X2=0.945 $Y2=0.178
r201 25 122 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.837 $Y=0.178 $X2=0.729 $Y2=0.178
r202 22 25 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0405 $X2=0.837 $Y2=0.178
r203 19 122 43.022 $w=2.6e-08 $l=5.4e-08 $layer=LISD $thickness=2.8e-08 $X=0.675
+ $Y=0.178 $X2=0.729 $Y2=0.178
r204 16 19 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.178
r205 10 86 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r206 10 13 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1355 $X2=0.567 $Y2=0.2025
r207 5 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r208 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r209 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%SE 2 5 7 10 13 15 19 22 23 24 31 33 41 44 45 46 47
+ 54 58 59 62 63 VSS
c80 63 VSS 5.91978e-19 $X=1.215 $Y=0.113
c81 62 VSS 0.00161589f $X=1.215 $Y=0.09
c82 59 VSS 2.63823e-19 $X=0.225 $Y=0.099
c83 58 VSS 5.90201e-19 $X=0.225 $Y=0.081
c84 54 VSS 0.00204823f $X=1.215 $Y=0.136
c85 47 VSS 0.0381131f $X=1.175 $Y=0.045
c86 46 VSS 0.00642311f $X=0.337 $Y=0.045
c87 45 VSS 0.00708497f $X=1.215 $Y=0.045
c88 44 VSS 0.00325301f $X=1.215 $Y=0.045
c89 41 VSS 0.00531f $X=0.225 $Y=0.045
c90 31 VSS 0.00110873f $X=0.225 $Y=0.126
c91 24 VSS 2.51525e-19 $X=0.279 $Y=0.135
c92 23 VSS 1.48251e-19 $X=0.261 $Y=0.135
c93 22 VSS 6.38823e-20 $X=0.258 $Y=0.135
c94 21 VSS 0.00134071f $X=0.255 $Y=0.135
c95 19 VSS 6.89032e-19 $X=0.297 $Y=0.135
c96 13 VSS 0.00265978f $X=1.215 $Y=0.136
c97 10 VSS 0.0624472f $X=1.215 $Y=0.0675
c98 5 VSS 0.0031928f $X=0.297 $Y=0.135
c99 2 VSS 0.063344f $X=0.297 $Y=0.0675
r100 62 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.09 $X2=1.215 $Y2=0.113
r101 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.081 $X2=0.225 $Y2=0.099
r102 54 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.136 $X2=1.215 $Y2=0.113
r103 46 47 56.9012 $w=1.8e-08 $l=8.38e-07 $layer=M2 $thickness=3.6e-08 $X=0.337
+ $Y=0.045 $X2=1.175 $Y2=0.045
r104 45 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.215 $Y2=0.09
r105 44 47 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.175 $Y2=0.045
r106 44 45 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.215 $Y=0.045 $X2=1.215
+ $Y2=0.045
r107 41 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.081
r108 40 46 7.60494 $w=1.8e-08 $l=1.12e-07 $layer=M2 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.337 $Y2=0.045
r109 40 41 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.225 $Y=0.045 $X2=0.225
+ $Y2=0.045
r110 31 59 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.099
r111 31 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r112 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.135 $X2=0.279 $Y2=0.135
r113 22 23 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.258
+ $Y=0.135 $X2=0.261 $Y2=0.135
r114 21 22 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.255
+ $Y=0.135 $X2=0.258 $Y2=0.135
r115 19 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.279 $Y2=0.135
r116 17 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.225 $Y2=0.135
r117 17 21 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.255 $Y2=0.135
r118 13 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.215 $Y=0.136 $X2=1.215
+ $Y2=0.136
r119 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.136 $X2=1.215 $Y2=0.2025
r120 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.0675 $X2=1.215 $Y2=0.136
r121 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r122 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r123 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%6 2 5 7 9 12 14 17 23 26 28 29 33 36 38 39 43 51
+ 57 58 65 VSS
c72 65 VSS 1.50983e-19 $X=1.161 $Y=0.2125
c73 58 VSS 5.45782e-19 $X=0.351 $Y=0.126
c74 57 VSS 8.0335e-19 $X=0.351 $Y=0.099
c75 51 VSS 0.00278599f $X=1.161 $Y=0.049
c76 43 VSS 3.76741e-19 $X=0.351 $Y=0.135
c77 39 VSS 9.89222e-19 $X=0.936 $Y=0.081
c78 38 VSS 0.00675922f $X=0.9 $Y=0.081
c79 36 VSS 0.00203618f $X=1.161 $Y=0.081
c80 33 VSS 8.1122e-19 $X=0.351 $Y=0.081
c81 29 VSS 6.98259e-19 $X=1.179 $Y=0.234
c82 28 VSS 0.00240687f $X=1.17 $Y=0.234
c83 26 VSS 0.00313492f $X=1.188 $Y=0.234
c84 23 VSS 4.80083e-20 $X=1.161 $Y=0.225
c85 17 VSS 0.00673327f $X=1.19 $Y=0.2025
c86 14 VSS 3.79317e-19 $X=1.205 $Y=0.2025
c87 12 VSS 0.0657106f $X=1.19 $Y=0.0675
c88 9 VSS 3.99927e-19 $X=1.205 $Y=0.0675
c89 5 VSS 0.00125227f $X=0.351 $Y=0.135
c90 2 VSS 0.0585837f $X=0.351 $Y=0.0675
r91 64 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.2 $X2=1.161 $Y2=0.2125
r92 57 58 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.099 $X2=0.351 $Y2=0.126
r93 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.161 $Y=0.049 $X2=1.161
+ $Y2=0.049
r94 43 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.126
r95 38 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.9
+ $Y=0.081 $X2=0.936 $Y2=0.081
r96 37 64 8.08025 $w=1.8e-08 $l=1.19e-07 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.2
r97 37 51 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.049
r98 36 39 15.2778 $w=1.8e-08 $l=2.25e-07 $layer=M2 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=0.936 $Y2=0.081
r99 36 37 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.161 $Y=0.081 $X2=1.161
+ $Y2=0.081
r100 33 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.099
r101 32 38 37.2778 $w=1.8e-08 $l=5.49e-07 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.9 $Y2=0.081
r102 32 33 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.081 $X2=0.351
+ $Y2=0.081
r103 28 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.17
+ $Y=0.234 $X2=1.179 $Y2=0.234
r104 26 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.188
+ $Y=0.234 $X2=1.179 $Y2=0.234
r105 23 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.225 $X2=1.161 $Y2=0.2125
r106 22 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.17 $Y2=0.234
r107 22 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.161 $Y2=0.225
r108 17 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.188 $Y=0.234
+ $X2=1.188 $Y2=0.234
r109 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.2025 $X2=1.19 $Y2=0.2025
r110 12 50 7.35229 $w=8.1e-08 $l=2.9e-08 $layer=LISD $thickness=2.8e-08 $X=1.19
+ $Y=0.0675 $X2=1.161 $Y2=0.0675
r111 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.0675 $X2=1.19 $Y2=0.0675
r112 5 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r113 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r114 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%D 2 5 7 11 VSS
c18 11 VSS 0.00145113f $X=0.405 $Y=0.134
c19 5 VSS 0.00106786f $X=0.405 $Y=0.135
c20 2 VSS 0.0589243f $X=0.405 $Y=0.0675
r21 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%SI 2 7 11 14 VSS
c21 14 VSS 0.00329293f $X=0.475 $Y=0.135
c22 11 VSS 0.00333153f $X=0.473 $Y=0.135
c23 2 VSS 0.0640988f $X=0.459 $Y=0.0675
r24 11 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.475 $Y=0.135 $X2=0.475
+ $Y2=0.135
r25 5 14 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.475 $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%9 2 5 7 10 13 15 17 20 22 25 27 29 36 43 45 51 55
+ 56 57 59 61 62 69 79 80 81 82 84 85 VSS
c76 86 VSS 5.63033e-20 $X=0.189 $Y=0.216
c77 85 VSS 4.28571e-19 $X=0.189 $Y=0.207
c78 84 VSS 4.04265e-19 $X=0.189 $Y=0.189
c79 82 VSS 2.19344e-19 $X=0.189 $Y=0.1485
c80 81 VSS 3.0092e-19 $X=0.189 $Y=0.144
c81 80 VSS 4.92067e-19 $X=0.189 $Y=0.121
c82 79 VSS 8.32677e-19 $X=0.189 $Y=0.099
c83 69 VSS 0.001222f $X=0.891 $Y=0.135
c84 62 VSS 0.0020506f $X=0.817 $Y=0.153
c85 61 VSS 0.00277455f $X=0.743 $Y=0.153
c86 59 VSS 0.00276294f $X=0.891 $Y=0.153
c87 57 VSS 0.00120333f $X=0.337 $Y=0.153
c88 56 VSS 0.00116325f $X=0.211 $Y=0.153
c89 55 VSS 9.40943e-19 $X=0.621 $Y=0.153
c90 51 VSS 5.62309e-19 $X=0.189 $Y=0.153
c91 48 VSS 5.43917e-20 $X=0.189 $Y=0.225
c92 45 VSS 0.00373046f $X=0.18 $Y=0.036
c93 43 VSS 0.00194932f $X=0.189 $Y=0.036
c94 36 VSS 5.26559e-19 $X=0.621 $Y=0.135
c95 29 VSS 0.00311772f $X=0.162 $Y=0.234
c96 27 VSS 0.00522825f $X=0.18 $Y=0.234
c97 25 VSS 0.00583113f $X=0.16 $Y=0.216
c98 20 VSS 0.00576958f $X=0.16 $Y=0.054
c99 13 VSS 0.00216055f $X=0.891 $Y=0.135
c100 10 VSS 0.0585656f $X=0.891 $Y=0.0405
c101 5 VSS 0.00201792f $X=0.621 $Y=0.135
c102 2 VSS 0.0601628f $X=0.621 $Y=0.0675
r103 85 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.207 $X2=0.189 $Y2=0.216
r104 84 85 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.207
r105 83 84 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.189
r106 81 82 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.1485
r107 80 81 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.121 $X2=0.189 $Y2=0.144
r108 79 80 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.099 $X2=0.189 $Y2=0.121
r109 61 62 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.743
+ $Y=0.153 $X2=0.817 $Y2=0.153
r110 59 62 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.817 $Y2=0.153
r111 59 69 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r112 56 57 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.211
+ $Y=0.153 $X2=0.337 $Y2=0.153
r113 54 61 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.743 $Y2=0.153
r114 54 57 19.284 $w=1.8e-08 $l=2.84e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.337 $Y2=0.153
r115 54 55 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.621 $Y=0.153 $X2=0.621
+ $Y2=0.153
r116 51 83 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.164
r117 51 82 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.1485
r118 50 56 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.211 $Y2=0.153
r119 50 51 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.153 $X2=0.189
+ $Y2=0.153
r120 48 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.216
r121 45 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r122 44 79 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.099
r123 43 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r124 43 44 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r125 40 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r126 36 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.153
r127 27 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.234 $X2=0.189 $Y2=0.225
r128 27 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.162 $Y2=0.234
r129 25 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r130 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r131 20 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r132 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r133 13 69 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.135 $X2=0.891
+ $Y2=0.135
r134 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.135 $X2=0.891 $Y2=0.2295
r135 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.0405 $X2=0.891 $Y2=0.135
r136 5 36 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r137 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2295
r138 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%10 2 7 9 10 13 14 17 19 22 27 28 29 31 33 38 40 46
+ 47 48 49 50 51 52 56 VSS
c49 58 VSS 5.19568e-19 $X=0.828 $Y=0.09
c50 57 VSS 3.9329e-19 $X=0.819 $Y=0.09
c51 56 VSS 4.29e-19 $X=0.837 $Y=0.09
c52 52 VSS 5.92996e-19 $X=0.837 $Y=0.207
c53 51 VSS 1.19762e-19 $X=0.837 $Y=0.167
c54 50 VSS 1.86299e-19 $X=0.837 $Y=0.165
c55 49 VSS 3.05662e-19 $X=0.837 $Y=0.14
c56 48 VSS 4.69487e-19 $X=0.837 $Y=0.122
c57 47 VSS 1.91116e-19 $X=0.837 $Y=0.101
c58 46 VSS 4.02479e-19 $X=0.837 $Y=0.225
c59 44 VSS 3.58124e-20 $X=0.81 $Y=0.0715
c60 40 VSS 0.00112276f $X=0.81 $Y=0.054
c61 33 VSS 0.00268883f $X=0.81 $Y=0.234
c62 31 VSS 0.00427376f $X=0.828 $Y=0.234
c63 30 VSS 2.64081e-19 $X=0.799 $Y=0.09
c64 29 VSS 0.00133552f $X=0.797 $Y=0.09
c65 28 VSS 0.00410211f $X=0.747 $Y=0.09
c66 27 VSS 4.49532e-19 $X=0.747 $Y=0.09
c67 24 VSS 4.45336e-20 $X=0.801 $Y=0.09
c68 22 VSS 0.0178238f $X=0.866 $Y=0.2295
c69 19 VSS 3.14771e-19 $X=0.881 $Y=0.2295
c70 17 VSS 2.5391e-19 $X=0.808 $Y=0.2295
c71 13 VSS 0.0201369f $X=0.81 $Y=0.0405
c72 9 VSS 6.29543e-19 $X=0.827 $Y=0.0405
c73 2 VSS 0.0580179f $X=0.729 $Y=0.0405
r74 57 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.819
+ $Y=0.09 $X2=0.828 $Y2=0.09
r75 56 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.09 $X2=0.828 $Y2=0.09
r76 55 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.09 $X2=0.819 $Y2=0.09
r77 51 52 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.167 $X2=0.837 $Y2=0.207
r78 50 51 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.165 $X2=0.837 $Y2=0.167
r79 49 50 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.14 $X2=0.837 $Y2=0.165
r80 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.122 $X2=0.837 $Y2=0.14
r81 47 48 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.101 $X2=0.837 $Y2=0.122
r82 46 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.207
r83 45 56 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.09
r84 45 47 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.101
r85 43 44 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.062 $X2=0.81 $Y2=0.0715
r86 40 43 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.054 $X2=0.81 $Y2=0.062
r87 38 55 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.09
r88 38 44 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.0715
r89 31 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r90 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.81 $Y2=0.234
r91 29 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.797
+ $Y=0.09 $X2=0.799 $Y2=0.09
r92 27 29 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.09 $X2=0.797 $Y2=0.09
r93 27 28 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.747 $Y=0.09 $X2=0.747
+ $Y2=0.09
r94 24 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.81 $Y2=0.09
r95 24 30 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.799 $Y2=0.09
r96 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2295 $X2=0.866 $Y2=0.2295
r97 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.808
+ $Y=0.2295 $X2=0.866 $Y2=0.2295
r98 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.234 $X2=0.81
+ $Y2=0.234
r99 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2295 $X2=0.808 $Y2=0.2295
r100 13 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.054 $X2=0.81
+ $Y2=0.054
r101 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.0405 $X2=0.81 $Y2=0.0405
r102 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.0405 $X2=0.81 $Y2=0.0405
r103 5 28 16.3636 $w=2.2e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.09 $X2=0.747 $Y2=0.09
r104 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.09 $X2=0.729 $Y2=0.2295
r105 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0405 $X2=0.729 $Y2=0.09
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%11 2 5 7 9 14 17 21 22 25 30 31 33 34 37 39 40 43
+ 44 45 46 48 50 51 52 53 54 55 56 59 61 62 65 VSS
c72 65 VSS 1.00162e-19 $X=0.693 $Y=0.131
c73 61 VSS 9.09188e-19 $X=0.72 $Y=0.131
c74 59 VSS 8.5526e-19 $X=0.783 $Y=0.131
c75 56 VSS 1.82087e-19 $X=0.693 $Y=0.216
c76 55 VSS 1.40959e-19 $X=0.693 $Y=0.207
c77 54 VSS 1.07888e-19 $X=0.693 $Y=0.189
c78 53 VSS 1.66071e-19 $X=0.693 $Y=0.171
c79 52 VSS 2.71272e-19 $X=0.693 $Y=0.165
c80 51 VSS 3.53682e-19 $X=0.693 $Y=0.153
c81 50 VSS 2.11704e-19 $X=0.693 $Y=0.225
c82 48 VSS 4.15228e-19 $X=0.693 $Y=0.114
c83 47 VSS 2.7378e-19 $X=0.693 $Y=0.106
c84 46 VSS 5.46003e-20 $X=0.693 $Y=0.099
c85 45 VSS 5.96385e-20 $X=0.693 $Y=0.081
c86 43 VSS 1.65771e-19 $X=0.693 $Y=0.062
c87 42 VSS 2.30403e-19 $X=0.693 $Y=0.122
c88 40 VSS 0.00145015f $X=0.6665 $Y=0.036
c89 39 VSS 0.00201121f $X=0.649 $Y=0.036
c90 37 VSS 0.00303728f $X=0.648 $Y=0.036
c91 34 VSS 0.00412969f $X=0.684 $Y=0.036
c92 33 VSS 0.00297725f $X=0.649 $Y=0.234
c93 32 VSS 2.2805e-19 $X=0.612 $Y=0.234
c94 31 VSS 0.00126734f $X=0.609 $Y=0.234
c95 30 VSS 0.0016591f $X=0.595 $Y=0.234
c96 25 VSS 0.00558865f $X=0.684 $Y=0.234
c97 24 VSS 5.62656e-19 $X=0.594 $Y=0.2295
c98 21 VSS 0.00254121f $X=0.594 $Y=0.2025
c99 18 VSS 1.02475e-19 $X=0.5895 $Y=0.216
c100 16 VSS 5.70081e-19 $X=0.648 $Y=0.0405
c101 10 VSS 7.61325e-20 $X=0.6435 $Y=0.054
c102 5 VSS 0.00231049f $X=0.783 $Y=0.131
c103 2 VSS 0.0591968f $X=0.783 $Y=0.0405
r104 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.131 $X2=0.738 $Y2=0.131
r105 59 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.131 $X2=0.738 $Y2=0.131
r106 57 65 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.693 $Y2=0.131
r107 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.72 $Y2=0.131
r108 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.207 $X2=0.693 $Y2=0.216
r109 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.189 $X2=0.693 $Y2=0.207
r110 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.171 $X2=0.693 $Y2=0.189
r111 52 53 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.165 $X2=0.693 $Y2=0.171
r112 51 52 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.153 $X2=0.693 $Y2=0.165
r113 50 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.225 $X2=0.693 $Y2=0.216
r114 49 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.131
r115 49 51 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.153
r116 47 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.106 $X2=0.693 $Y2=0.114
r117 46 47 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.099 $X2=0.693 $Y2=0.106
r118 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.081 $X2=0.693 $Y2=0.099
r119 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.063 $X2=0.693 $Y2=0.081
r120 43 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.062 $X2=0.693 $Y2=0.063
r121 42 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.131
r122 42 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.114
r123 41 43 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.045 $X2=0.693 $Y2=0.062
r124 39 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.649
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r125 36 39 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.649 $Y2=0.036
r126 36 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r127 34 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.036 $X2=0.693 $Y2=0.045
r128 34 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r129 32 33 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.649 $Y2=0.234
r130 31 32 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.609
+ $Y=0.234 $X2=0.612 $Y2=0.234
r131 30 31 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.595
+ $Y=0.234 $X2=0.609 $Y2=0.234
r132 27 30 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.595 $Y2=0.234
r133 25 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.234 $X2=0.693 $Y2=0.225
r134 25 33 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.234 $X2=0.649 $Y2=0.234
r135 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2295 $X2=0.594 $Y2=0.2295
r136 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r137 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.594 $Y2=0.2295
r138 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.5895 $Y2=0.189
r139 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.189 $X2=0.5895 $Y2=0.189
r140 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r141 13 37 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r142 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.648 $Y2=0.0405
r143 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.6435 $Y2=0.081
r144 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.081 $X2=0.6435 $Y2=0.081
r145 5 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.131 $X2=0.783
+ $Y2=0.131
r146 5 7 369.03 $w=2e-08 $l=9.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.131 $X2=0.783 $Y2=0.2295
r147 2 5 339.058 $w=2e-08 $l=9.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.131
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%12 2 5 7 9 12 14 17 21 25 26 30 31 35 36 37 43 VSS
c33 43 VSS 0.00419842f $X=1.098 $Y=0.234
c34 42 VSS 0.00204425f $X=1.107 $Y=0.234
c35 37 VSS 0.00106107f $X=1.107 $Y=0.171
c36 36 VSS 0.00114275f $X=1.107 $Y=0.117
c37 35 VSS 0.00149546f $X=1.107 $Y=0.225
c38 33 VSS 7.70286e-19 $X=1.073 $Y=0.036
c39 32 VSS 4.41014e-19 $X=1.066 $Y=0.036
c40 31 VSS 0.00146362f $X=1.062 $Y=0.036
c41 30 VSS 0.00481311f $X=1.044 $Y=0.036
c42 26 VSS 0.00226308f $X=1.008 $Y=0.036
c43 25 VSS 0.00460331f $X=1.098 $Y=0.036
c44 21 VSS 7.16657e-19 $X=0.999 $Y=0.105
c45 17 VSS 0.00426839f $X=1.078 $Y=0.2295
c46 12 VSS 0.00485453f $X=1.078 $Y=0.0405
c47 5 VSS 0.00227106f $X=0.999 $Y=0.1055
c48 2 VSS 0.0590816f $X=0.999 $Y=0.0405
r49 43 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r50 42 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r51 39 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.098 $Y2=0.234
r52 36 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.117 $X2=1.107 $Y2=0.171
r53 35 42 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.234
r54 35 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.171
r55 34 36 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.045 $X2=1.107 $Y2=0.117
r56 32 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.066
+ $Y=0.036 $X2=1.073 $Y2=0.036
r57 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=1.062
+ $Y=0.036 $X2=1.066 $Y2=0.036
r58 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=1.062 $Y2=0.036
r59 28 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.036 $X2=1.073 $Y2=0.036
r60 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.008
+ $Y=0.036 $X2=1.044 $Y2=0.036
r61 25 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.098 $Y=0.036 $X2=1.107 $Y2=0.045
r62 25 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.036 $X2=1.08 $Y2=0.036
r63 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.999 $Y=0.045 $X2=1.008 $Y2=0.036
r64 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.045 $X2=0.999 $Y2=0.105
r65 17 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234 $X2=1.08
+ $Y2=0.234
r66 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2295 $X2=1.078 $Y2=0.2295
r67 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.036 $X2=1.08
+ $Y2=0.036
r68 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.0405 $X2=1.078 $Y2=0.0405
r69 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.105 $X2=0.999
+ $Y2=0.105
r70 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.1055 $X2=0.999 $Y2=0.2295
r71 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.0405 $X2=0.999 $Y2=0.1055
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%13 2 7 10 13 15 17 18 21 22 23 26 27 32 33 35 38
+ 39 40 41 43 46 47 50 60 65 68 70 71 78 VSS
c70 78 VSS 0.00312516f $X=1.269 $Y=0.136
c71 71 VSS 0.00157729f $X=1.229 $Y=0.153
c72 70 VSS 0.00790597f $X=1.175 $Y=0.153
c73 68 VSS 0.00415759f $X=1.269 $Y=0.153
c74 65 VSS 1.90327e-19 $X=0.945 $Y=0.153
c75 60 VSS 0.0033916f $X=0.936 $Y=0.234
c76 59 VSS 0.00253671f $X=0.945 $Y=0.234
c77 50 VSS 4.04001e-19 $X=1.053 $Y=0.14
c78 47 VSS 3.26354e-19 $X=1.008 $Y=0.162
c79 46 VSS 0.00199114f $X=0.99 $Y=0.162
c80 44 VSS 0.00235839f $X=1.044 $Y=0.162
c81 43 VSS 0.00104404f $X=0.945 $Y=0.225
c82 41 VSS 2.07499e-19 $X=0.945 $Y=0.136
c83 40 VSS 2.77769e-19 $X=0.945 $Y=0.119
c84 39 VSS 2.61356e-19 $X=0.945 $Y=0.101
c85 38 VSS 6.393e-19 $X=0.945 $Y=0.081
c86 37 VSS 3.04251e-19 $X=0.945 $Y=0.153
c87 35 VSS 0.00136569f $X=0.92 $Y=0.036
c88 34 VSS 4.8751e-19 $X=0.904 $Y=0.036
c89 33 VSS 0.00146362f $X=0.9 $Y=0.036
c90 32 VSS 0.00358427f $X=0.882 $Y=0.036
c91 27 VSS 0.00347893f $X=0.936 $Y=0.036
c92 26 VSS 0.00276615f $X=0.918 $Y=0.2295
c93 22 VSS 5.63046e-19 $X=0.935 $Y=0.2295
c94 21 VSS 0.0201056f $X=0.864 $Y=0.0405
c95 17 VSS 5.63046e-19 $X=0.881 $Y=0.0405
c96 13 VSS 0.00278011f $X=1.269 $Y=0.136
c97 10 VSS 0.0625639f $X=1.269 $Y=0.0675
c98 5 VSS 0.00302777f $X=1.053 $Y=0.14
c99 2 VSS 0.0627731f $X=1.053 $Y=0.0405
r100 70 71 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=1.175
+ $Y=0.153 $X2=1.229 $Y2=0.153
r101 68 71 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.269
+ $Y=0.153 $X2=1.229 $Y2=0.153
r102 68 78 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.269 $Y=0.153 $X2=1.269
+ $Y2=0.153
r103 64 70 15.6173 $w=1.8e-08 $l=2.3e-07 $layer=M2 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=1.175 $Y2=0.153
r104 64 65 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.945 $Y=0.153 $X2=0.945
+ $Y2=0.153
r105 60 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r106 59 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r107 56 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.234 $X2=0.936 $Y2=0.234
r108 48 50 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.153 $X2=1.053 $Y2=0.14
r109 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.99
+ $Y=0.162 $X2=1.008 $Y2=0.162
r110 45 65 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.945 $Y2=0.162
r111 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.99 $Y2=0.162
r112 44 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.162 $X2=1.053 $Y2=0.153
r113 44 47 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.162 $X2=1.008 $Y2=0.162
r114 43 59 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.234
r115 42 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.162
r116 42 43 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.225
r117 40 41 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.119 $X2=0.945 $Y2=0.136
r118 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.101 $X2=0.945 $Y2=0.119
r119 38 39 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.081 $X2=0.945 $Y2=0.101
r120 37 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.162
r121 37 41 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.136
r122 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.081
r123 34 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.904
+ $Y=0.036 $X2=0.92 $Y2=0.036
r124 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.036 $X2=0.904 $Y2=0.036
r125 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r126 29 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r127 27 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r128 27 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.92 $Y2=0.036
r129 26 56 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.234
+ $X2=0.918 $Y2=0.234
r130 23 26 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.2295 $X2=0.918 $Y2=0.2295
r131 22 26 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.935 $Y=0.2295 $X2=0.918 $Y2=0.2295
r132 21 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036
+ $X2=0.864 $Y2=0.036
r133 18 21 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.864 $Y2=0.0405
r134 17 21 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0405 $X2=0.864 $Y2=0.0405
r135 13 78 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.269 $Y=0.136 $X2=1.269
+ $Y2=0.136
r136 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.136 $X2=1.269 $Y2=0.2025
r137 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.0675 $X2=1.269 $Y2=0.136
r138 5 50 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.053 $Y=0.14 $X2=1.053
+ $Y2=0.14
r139 5 7 335.312 $w=2e-08 $l=8.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.14 $X2=1.053 $Y2=0.2295
r140 2 5 372.777 $w=2e-08 $l=9.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.0405 $X2=1.053 $Y2=0.14
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%14 1 4 6 11 14 21 23 24 25 VSS
c29 26 VSS 0.00225833f $X=0.485 $Y=0.234
c30 25 VSS 0.00141737f $X=0.461 $Y=0.234
c31 24 VSS 0.0134342f $X=0.447 $Y=0.234
c32 23 VSS 0.00523898f $X=0.309 $Y=0.234
c33 21 VSS 0.00168783f $X=0.486 $Y=0.234
c34 14 VSS 0.0195485f $X=0.542 $Y=0.2025
c35 11 VSS 3.25039e-19 $X=0.557 $Y=0.2025
c36 9 VSS 4.57278e-19 $X=0.484 $Y=0.2025
c37 4 VSS 0.00250858f $X=0.272 $Y=0.2025
c38 1 VSS 3.31752e-19 $X=0.287 $Y=0.2025
r39 25 26 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.461
+ $Y=0.234 $X2=0.485 $Y2=0.234
r40 24 25 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.234 $X2=0.461 $Y2=0.234
r41 23 24 9.37037 $w=1.8e-08 $l=1.38e-07 $layer=M1 $thickness=3.6e-08 $X=0.309
+ $Y=0.234 $X2=0.447 $Y2=0.234
r42 21 26 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.485 $Y2=0.234
r43 17 23 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.309 $Y2=0.234
r44 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.542 $Y2=0.2025
r45 9 14 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.484
+ $Y=0.2025 $X2=0.542 $Y2=0.2025
r46 9 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r47 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.2025 $X2=0.484 $Y2=0.2025
r48 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r49 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.272 $Y2=0.2025
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%16 1 2 5 6 7 10 12 18 20 21 22 23 24 25 VSS
c21 25 VSS 3.8923e-20 $X=0.423 $Y=0.198
c22 24 VSS 8.46035e-21 $X=0.414 $Y=0.198
c23 23 VSS 0.00116854f $X=0.396 $Y=0.198
c24 22 VSS 0.00154511f $X=0.379 $Y=0.198
c25 21 VSS 8.46035e-21 $X=0.36 $Y=0.198
c26 20 VSS 2.61077e-19 $X=0.342 $Y=0.198
c27 18 VSS 3.31089e-19 $X=0.432 $Y=0.198
c28 12 VSS 5.32749e-19 $X=0.324 $Y=0.198
c29 10 VSS 0.00631853f $X=0.432 $Y=0.2025
c30 6 VSS 5.67296e-19 $X=0.449 $Y=0.2025
c31 5 VSS 0.00790786f $X=0.324 $Y=0.2025
c32 1 VSS 6.05629e-19 $X=0.341 $Y=0.2025
r33 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.423 $Y2=0.198
r34 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.414 $Y2=0.198
r35 22 23 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.198 $X2=0.396 $Y2=0.198
r36 21 22 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.198 $X2=0.379 $Y2=0.198
r37 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r38 18 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.423 $Y2=0.198
r39 12 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.342 $Y2=0.198
r40 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r41 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r42 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r43 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198 $X2=0.324
+ $Y2=0.198
r44 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
r45 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%QN 1 6 9 14 15 16 19 22 30 VSS
c9 30 VSS 0.0042609f $X=1.314 $Y=0.234
c10 29 VSS 0.00278493f $X=1.323 $Y=0.234
c11 22 VSS 0.00408512f $X=1.314 $Y=0.036
c12 21 VSS 0.00278493f $X=1.323 $Y=0.036
c13 19 VSS 0.00657307f $X=1.296 $Y=0.036
c14 16 VSS 0.00487569f $X=1.323 $Y=0.2
c15 15 VSS 0.00226847f $X=1.323 $Y=0.09
c16 12 VSS 0.00136544f $X=1.323 $Y=0.225
c17 9 VSS 0.00693684f $X=1.294 $Y=0.2025
c18 4 VSS 3.77696e-19 $X=1.294 $Y=0.0675
r19 30 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.314
+ $Y=0.234 $X2=1.3185 $Y2=0.234
r20 29 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.234 $X2=1.3185 $Y2=0.234
r21 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.234 $X2=1.314 $Y2=0.234
r22 22 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.314
+ $Y=0.036 $X2=1.3185 $Y2=0.036
r23 21 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.036 $X2=1.3185 $Y2=0.036
r24 18 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.036 $X2=1.314 $Y2=0.036
r25 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.036 $X2=1.296
+ $Y2=0.036
r26 15 16 7.46914 $w=1.8e-08 $l=1.1e-07 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.09 $X2=1.323 $Y2=0.2
r27 14 16 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.223 $X2=1.323 $Y2=0.2
r28 12 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.225 $X2=1.323 $Y2=0.234
r29 12 14 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.225 $X2=1.323 $Y2=0.223
r30 11 21 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.045 $X2=1.323 $Y2=0.036
r31 11 15 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.045 $X2=1.323 $Y2=0.09
r32 9 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.234 $X2=1.296
+ $Y2=0.234
r33 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=1.279
+ $Y=0.2025 $X2=1.294 $Y2=0.2025
r34 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.296
+ $Y=0.0675 $X2=1.296 $Y2=0.036
r35 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.279
+ $Y=0.0675 $X2=1.294 $Y2=0.0675
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%19 1 6 9 VSS
c10 9 VSS 0.0140217f $X=0.704 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.719 $Y=0.2295
c12 4 VSS 2.70811e-19 $X=0.646 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.646
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.631
+ $Y=0.2295 $X2=0.646 $Y2=0.2295
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%20 1 6 9 VSS
c9 9 VSS 0.0145746f $X=0.974 $Y=0.0405
c10 6 VSS 3.14771e-19 $X=0.989 $Y=0.0405
c11 4 VSS 2.65708e-19 $X=0.916 $Y=0.0405
r12 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r13 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.916
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r14 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.901
+ $Y=0.0405 $X2=0.916 $Y2=0.0405
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%22 1 2 VSS
c2 1 VSS 0.00203573f $X=0.719 $Y=0.0405
r3 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0405 $X2=0.685 $Y2=0.0405
.ends

.subckt PM_SDFLX1_ASAP7_75T_SRAM%23 1 2 VSS
c0 1 VSS 0.00214045f $X=0.989 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.2295 $X2=0.955 $Y2=0.2295
.ends


* END of "./SDFLx1_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt SDFLx1_ASAP7_75t_SRAM  VSS VDD CLK SE D SI QN
* 
* QN	QN
* SI	SI
* D	D
* SE	SE
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_9_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_SE_M2_g noxref_15 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 noxref_21 N_6_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 noxref_17 N_D_M4_g noxref_21 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 noxref_15 N_SI_M5_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 N_11_M6_d N_9_M6_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M7 N_22_M7_d N_4_M7_g N_11_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M8 VSS N_10_M8_g N_22_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.027
M9 N_10_M9_d N_11_M9_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_13_M10_d N_4_M10_g N_10_M10_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.827 $Y=0.027
M11 N_20_M11_d N_9_M11_g N_13_M11_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.027
M12 VSS N_12_M12_g N_20_M12_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.027
M13 N_12_M13_d N_13_M13_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.027
M14 VSS N_SE_M14_g N_6_M14_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.027
M15 N_QN_M15_d N_13_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M16 VDD N_CLK_M16_g N_4_M16_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M17 N_9_M17_d N_4_M17_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M18 N_16_M18_d N_SE_M18_g N_14_M18_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M19 VDD N_6_M19_g N_16_M19_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M20 N_16_M20_d N_D_M20_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M21 N_14_M21_d N_SI_M21_g N_16_M21_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M22 N_11_M22_d N_4_M22_g N_14_M22_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M23 N_19_M23_d N_9_M23_g N_11_M23_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.611 $Y=0.216
M24 VDD N_10_M24_g N_19_M24_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.216
M25 N_10_M25_d N_11_M25_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M26 N_13_M26_d N_9_M26_g N_10_M26_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.216
M27 N_23_M27_d N_4_M27_g N_13_M27_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.935 $Y=0.216
M28 VDD N_12_M28_g N_23_M28_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.216
M29 N_12_M29_d N_13_M29_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.216
M30 VDD N_SE_M30_g N_6_M30_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.162
M31 N_QN_M31_d N_13_M31_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
*
* 
* .include "SDFLx1_ASAP7_75t_SRAM.pex.sp.SDFLX1_ASAP7_75T_SRAM.pxi"
* BEGIN of "./SDFLx1_ASAP7_75t_SRAM.pex.sp.SDFLX1_ASAP7_75T_SRAM.pxi"
* File: SDFLx1_ASAP7_75t_SRAM.pex.sp.SDFLX1_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 13:04:33 2017
* 
x_PM_SDFLX1_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M16_g N_CLK_c_3_p CLK
+ VSS PM_SDFLX1_ASAP7_75T_SRAM%CLK
x_PM_SDFLX1_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_14_n N_4_M17_g N_4_c_25_p N_4_M22_g
+ N_4_M7_g N_4_c_91_p N_4_M10_g N_4_c_75_p N_4_c_24_p N_4_M27_g N_4_M0_s
+ N_4_c_15_n N_4_M16_s N_4_c_16_n N_4_c_17_n N_4_c_18_n N_4_c_41_p N_4_c_19_n
+ N_4_c_59_p N_4_c_26_p N_4_c_27_p N_4_c_37_p N_4_c_28_p N_4_c_20_n N_4_c_21_p
+ N_4_c_29_p N_4_c_56_p VSS PM_SDFLX1_ASAP7_75T_SRAM%4
x_PM_SDFLX1_ASAP7_75T_SRAM%SE N_SE_M2_g N_SE_c_138_p N_SE_M18_g N_SE_M14_g
+ N_SE_c_175_p N_SE_M30_g N_SE_c_144_p N_SE_c_189_p N_SE_c_187_p N_SE_c_205_p
+ N_SE_c_135_n SE N_SE_c_134_n N_SE_c_139_p N_SE_c_140_p N_SE_c_136_n
+ N_SE_c_141_p N_SE_c_142_p N_SE_c_153_p N_SE_c_158_p N_SE_c_147_p N_SE_c_186_p
+ VSS PM_SDFLX1_ASAP7_75T_SRAM%SE
x_PM_SDFLX1_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_217_n N_6_M19_g N_6_M14_s N_6_c_218_n
+ N_6_M30_s N_6_c_221_n N_6_c_256_p N_6_c_266_p N_6_c_253_p N_6_c_262_p
+ N_6_c_270_p N_6_c_248_p N_6_c_214_n N_6_c_215_n N_6_c_223_n N_6_c_224_n
+ N_6_c_227_n N_6_c_228_n N_6_c_255_p VSS PM_SDFLX1_ASAP7_75T_SRAM%6
x_PM_SDFLX1_ASAP7_75T_SRAM%D N_D_M4_g N_D_c_288_n N_D_M20_g D VSS
+ PM_SDFLX1_ASAP7_75T_SRAM%D
x_PM_SDFLX1_ASAP7_75T_SRAM%SI N_SI_M5_g N_SI_M21_g SI N_SI_c_309_n VSS
+ PM_SDFLX1_ASAP7_75T_SRAM%SI
x_PM_SDFLX1_ASAP7_75T_SRAM%9 N_9_M6_g N_9_c_330_n N_9_M23_g N_9_M11_g N_9_c_333_n
+ N_9_M26_g N_9_M1_d N_9_c_400_p N_9_M17_d N_9_c_334_n N_9_c_336_n N_9_c_337_n
+ N_9_c_341_n N_9_c_360_n N_9_c_325_n N_9_c_343_n N_9_c_345_n N_9_c_346_n
+ N_9_c_348_n N_9_c_349_n N_9_c_350_n N_9_c_365_n N_9_c_354_n N_9_c_326_n
+ N_9_c_327_n N_9_c_355_n N_9_c_356_n N_9_c_357_n N_9_c_359_n VSS
+ PM_SDFLX1_ASAP7_75T_SRAM%9
x_PM_SDFLX1_ASAP7_75T_SRAM%10 N_10_M8_g N_10_M24_g N_10_M10_s N_10_M9_d
+ N_10_c_405_n N_10_M25_d N_10_c_406_n N_10_M26_s N_10_c_408_n N_10_c_419_n
+ N_10_c_420_n N_10_c_417_n N_10_c_448_p N_10_c_425_n N_10_c_422_n N_10_c_418_n
+ N_10_c_435_p N_10_c_449_p N_10_c_410_n N_10_c_437_p N_10_c_411_n N_10_c_412_n
+ N_10_c_413_n N_10_c_415_n VSS PM_SDFLX1_ASAP7_75T_SRAM%10
x_PM_SDFLX1_ASAP7_75T_SRAM%11 N_11_M9_g N_11_c_485_n N_11_M25_g N_11_M6_d N_11_M7_s
+ N_11_M22_d N_11_c_453_n N_11_M23_s N_11_c_515_p N_11_c_455_n N_11_c_456_n
+ N_11_c_487_n N_11_c_457_n N_11_c_477_n N_11_c_478_n N_11_c_479_n N_11_c_480_n
+ N_11_c_498_n N_11_c_458_n N_11_c_459_n N_11_c_489_n N_11_c_518_p N_11_c_490_n
+ N_11_c_460_n N_11_c_461_n N_11_c_463_n N_11_c_466_n N_11_c_519_p N_11_c_471_n
+ N_11_c_472_n N_11_c_473_n N_11_c_475_n VSS PM_SDFLX1_ASAP7_75T_SRAM%11
x_PM_SDFLX1_ASAP7_75T_SRAM%12 N_12_M12_g N_12_c_544_p N_12_M28_g N_12_M13_d
+ N_12_c_529_n N_12_M29_d N_12_c_531_n N_12_c_523_n N_12_c_524_n N_12_c_525_n
+ N_12_c_526_n N_12_c_527_n N_12_c_535_n N_12_c_528_n N_12_c_538_n N_12_c_553_p
+ VSS PM_SDFLX1_ASAP7_75T_SRAM%12
x_PM_SDFLX1_ASAP7_75T_SRAM%13 N_13_M13_g N_13_M29_g N_13_M15_g N_13_c_565_n
+ N_13_M31_g N_13_M11_s N_13_M10_d N_13_c_556_n N_13_M27_s N_13_M26_d
+ N_13_c_558_n N_13_c_567_n N_13_c_568_n N_13_c_569_n N_13_c_570_n N_13_c_571_n
+ N_13_c_559_n N_13_c_589_n N_13_c_560_n N_13_c_561_n N_13_c_624_p N_13_c_609_n
+ N_13_c_611_n N_13_c_562_n N_13_c_563_n N_13_c_572_n N_13_c_573_n N_13_c_574_n
+ N_13_c_576_n VSS PM_SDFLX1_ASAP7_75T_SRAM%13
x_PM_SDFLX1_ASAP7_75T_SRAM%14 N_14_M18_s N_14_c_625_n N_14_M21_d N_14_M22_s
+ N_14_c_626_n N_14_c_636_n N_14_c_628_n N_14_c_633_n N_14_c_629_n VSS
+ PM_SDFLX1_ASAP7_75T_SRAM%14
x_PM_SDFLX1_ASAP7_75T_SRAM%16 N_16_M19_s N_16_M18_d N_16_c_668_n N_16_M21_s
+ N_16_M20_d N_16_c_670_n N_16_c_654_n N_16_c_655_n N_16_c_656_n N_16_c_657_n
+ N_16_c_658_n N_16_c_659_n N_16_c_660_n N_16_c_661_n VSS
+ PM_SDFLX1_ASAP7_75T_SRAM%16
x_PM_SDFLX1_ASAP7_75T_SRAM%QN N_QN_M15_d N_QN_M31_d N_QN_c_677_n QN N_QN_c_675_n
+ N_QN_c_681_n N_QN_c_678_n N_QN_c_676_n N_QN_c_679_n VSS
+ PM_SDFLX1_ASAP7_75T_SRAM%QN
x_PM_SDFLX1_ASAP7_75T_SRAM%19 N_19_M23_d N_19_M24_s N_19_c_685_n VSS
+ PM_SDFLX1_ASAP7_75T_SRAM%19
x_PM_SDFLX1_ASAP7_75T_SRAM%20 N_20_M11_d N_20_M12_s N_20_c_694_n VSS
+ PM_SDFLX1_ASAP7_75T_SRAM%20
x_PM_SDFLX1_ASAP7_75T_SRAM%22 N_22_M8_s N_22_M7_d VSS PM_SDFLX1_ASAP7_75T_SRAM%22
x_PM_SDFLX1_ASAP7_75T_SRAM%23 N_23_M28_s N_23_M27_d VSS PM_SDFLX1_ASAP7_75T_SRAM%23
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_CLK_c_2_p N_4_c_14_n 9.79748e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_CLK_c_3_p N_4_c_15_n 2.66516e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.054
cc_4 N_CLK_c_3_p N_4_c_16_n 3.97017e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.081
cc_5 N_CLK_c_3_p N_4_c_17_n 0.00342695f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.164
cc_6 N_CLK_c_3_p N_4_c_18_n 4.97741e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.036
cc_7 N_CLK_c_3_p N_4_c_19_n 0.00171874f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_8 N_CLK_c_3_p N_4_c_20_n 8.1621e-19 $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.189
cc_9 N_CLK_c_3_p N_SE_c_134_n 2.45198e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_10 N_CLK_c_3_p N_9_c_325_n 6.32319e-19 $X=0.081 $Y=0.135 $X2=0.071 $Y2=0.054
cc_11 N_CLK_c_3_p N_9_c_326_n 0.00114506f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_12 N_CLK_c_3_p N_9_c_327_n 4.4946e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_13 N_4_c_21_p N_SE_c_135_n 4.53301e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_14 N_4_c_21_p N_SE_c_136_n 3.907e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_15 N_4_c_21_p N_6_c_214_n 0.0011956f $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_16 N_4_c_24_p N_6_c_215_n 3.37164e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_17 N_4_c_25_p N_SI_M5_g 2.94371e-19 $X=0.567 $Y=0.1355 $X2=0.081 $Y2=0.054
cc_18 N_4_c_26_p SI 0.00114959f $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.135
cc_19 N_4_c_27_p SI 0.00114959f $X=0.567 $Y=0.18 $X2=0.081 $Y2=0.135
cc_20 N_4_c_28_p SI 0.00239259f $X=0.567 $Y=0.189 $X2=0.081 $Y2=0.135
cc_21 N_4_c_29_p SI 0.00167124f $X=0.729 $Y=0.189 $X2=0.081 $Y2=0.135
cc_22 N_4_c_25_p N_SI_c_309_n 5.18435e-19 $X=0.567 $Y=0.1355 $X2=0 $Y2=0
cc_23 N_4_c_25_p N_9_M6_g 0.00365763f $X=0.567 $Y=0.1355 $X2=0.081 $Y2=0.054
cc_24 N_4_M7_g N_9_M6_g 0.00355599f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_25 N_4_c_25_p N_9_c_330_n 9.97803e-19 $X=0.567 $Y=0.1355 $X2=0.081 $Y2=0.135
cc_26 N_4_M10_g N_9_M11_g 0.00355599f $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_27 N_4_c_24_p N_9_M11_g 0.00605856f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.135
cc_28 N_4_c_24_p N_9_c_333_n 0.00180656f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_29 N_4_c_37_p N_9_c_334_n 3.29411e-19 $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_30 N_4_c_20_n N_9_c_334_n 3.38615e-19 $X=0.175 $Y=0.189 $X2=0 $Y2=0
cc_31 N_4_c_21_p N_9_c_336_n 2.67996e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_32 N_4_M1_g N_9_c_337_n 2.57258e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_33 N_4_c_41_p N_9_c_337_n 3.72764e-19 $X=0.054 $Y=0.234 $X2=0 $Y2=0
cc_34 N_4_c_37_p N_9_c_337_n 0.00209054f $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_35 N_4_c_20_n N_9_c_337_n 2.67996e-19 $X=0.175 $Y=0.189 $X2=0 $Y2=0
cc_36 N_4_c_26_p N_9_c_341_n 0.00279251f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_20_n N_9_c_325_n 2.60625e-19 $X=0.175 $Y=0.189 $X2=0 $Y2=0
cc_38 N_4_c_37_p N_9_c_343_n 9.44301e-19 $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_39 N_4_c_21_p N_9_c_343_n 2.46239e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_40 N_4_c_29_p N_9_c_345_n 3.80004e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_41 N_4_c_19_n N_9_c_346_n 3.53344e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_42 N_4_c_21_p N_9_c_346_n 0.0235609f $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_43 N_4_c_29_p N_9_c_348_n 0.0235609f $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_44 N_4_c_24_p N_9_c_349_n 5.51712e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_45 N_4_c_24_p N_9_c_350_n 0.00168667f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_46 N_4_c_26_p N_9_c_350_n 9.87747e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_47 N_4_c_28_p N_9_c_350_n 2.46239e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_48 N_4_c_56_p N_9_c_350_n 2.81643e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_49 N_4_c_24_p N_9_c_354_n 0.00123876f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_50 N_4_c_19_n N_9_c_355_n 9.44301e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_51 N_4_c_59_p N_9_c_356_n 9.44301e-19 $X=0.135 $Y=0.18 $X2=0 $Y2=0
cc_52 N_4_c_37_p N_9_c_357_n 0.00103771f $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_53 N_4_c_21_p N_9_c_357_n 5.9968e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_54 N_4_c_21_p N_9_c_359_n 4.92128e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_55 N_4_M7_g N_10_M8_g 0.00341068f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_56 N_4_M10_g N_10_M8_g 2.13359e-19 $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_57 N_4_c_24_p N_10_M8_g 0.00205997f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_58 N_4_c_56_p N_10_M8_g 3.19768e-19 $X=0.729 $Y=0.18 $X2=0.081 $Y2=0.054
cc_59 N_4_c_24_p N_10_c_405_n 5.49754e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_60 N_4_c_24_p N_10_c_406_n 2.12581e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_61 N_4_c_24_p N_10_M26_s 2.50995e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_62 N_4_M10_g N_10_c_408_n 0.00200065f $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_63 N_4_c_24_p N_10_c_408_n 0.00303373f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_64 N_4_M10_g N_10_c_410_n 2.74825e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_65 N_4_M10_g N_10_c_411_n 2.10136e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_66 N_4_c_56_p N_10_c_412_n 6.73839e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_67 N_4_c_75_p N_10_c_413_n 0.00195059f $X=0.837 $Y=0.178 $X2=0 $Y2=0
cc_68 N_4_c_24_p N_10_c_413_n 0.00191847f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_69 N_4_M10_g N_10_c_415_n 3.61755e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_70 N_4_M7_g N_11_M9_g 2.13359e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_71 N_4_M10_g N_11_M9_g 0.00341068f $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_72 N_4_c_24_p N_11_M9_g 0.00302156f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_73 N_4_c_26_p N_11_c_453_n 7.70794e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_74 N_4_c_28_p N_11_c_453_n 0.001307f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_75 N_4_c_28_p N_11_c_455_n 0.00138499f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_76 N_4_c_29_p N_11_c_456_n 0.00160025f $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_77 N_4_M7_g N_11_c_457_n 4.38308e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_78 N_4_M7_g N_11_c_458_n 2.0845e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_79 N_4_M7_g N_11_c_459_n 2.27141e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_80 N_4_c_24_p N_11_c_460_n 0.0361494f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_81 N_4_c_24_p N_11_c_461_n 2.38252e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_82 N_4_c_56_p N_11_c_461_n 0.00386452f $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_83 N_4_c_91_p N_11_c_463_n 7.00743e-19 $X=0.675 $Y=0.178 $X2=0 $Y2=0
cc_84 N_4_c_24_p N_11_c_463_n 7.89771e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_85 N_4_c_29_p N_11_c_463_n 4.88732e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_86 N_4_M7_g N_11_c_466_n 2.5554e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_87 N_4_c_24_p N_11_c_466_n 3.47488e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_88 N_4_c_28_p N_11_c_466_n 2.13133e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_89 N_4_c_29_p N_11_c_466_n 4.32971e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_90 N_4_c_56_p N_11_c_466_n 2.60223e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_91 N_4_c_24_p N_11_c_471_n 4.76652e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_92 N_4_c_24_p N_11_c_472_n 4.41163e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_93 N_4_c_24_p N_11_c_473_n 3.33141e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_94 N_4_c_56_p N_11_c_473_n 9.1388e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_95 N_4_M7_g N_11_c_475_n 2.12062e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_96 N_4_c_24_p N_12_M12_g 0.00341068f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_97 N_4_c_24_p N_13_M13_g 2.13359e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_98 N_4_c_24_p N_13_c_556_n 8.27183e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_99 N_4_c_24_p N_13_M27_s 3.37661e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_100 N_4_c_24_p N_13_c_558_n 0.00145657f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_101 N_4_c_24_p N_13_c_559_n 3.13444e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_102 N_4_c_24_p N_13_c_560_n 2.6418e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_103 N_4_c_24_p N_13_c_561_n 0.00294656f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_104 N_4_c_24_p N_13_c_562_n 3.75802e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_105 N_4_c_24_p N_13_c_563_n 5.46321e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_106 N_4_c_21_p N_14_c_625_n 4.92298e-19 $X=0.371 $Y=0.189 $X2=0.081 $Y2=0.135
cc_107 N_4_c_26_p N_14_c_626_n 9.68946e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_108 N_4_c_29_p N_14_c_626_n 6.49405e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_109 N_4_c_21_p N_14_c_628_n 7.84624e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_110 N_4_c_29_p N_14_c_629_n 6.22262e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_111 N_4_c_21_p N_16_c_654_n 2.13751e-19 $X=0.371 $Y=0.189 $X2=0.081 $Y2=0.135
cc_112 N_4_c_29_p N_16_c_655_n 7.1298e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_113 N_4_c_21_p N_16_c_656_n 6.46208e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_114 N_4_c_21_p N_16_c_657_n 4.50553e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_115 N_4_c_21_p N_16_c_658_n 2.85141e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_116 N_4_c_29_p N_16_c_659_n 4.60071e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_117 N_4_c_29_p N_16_c_660_n 4.38038e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_118 N_4_c_29_p N_16_c_661_n 2.31538e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_119 VSS N_4_c_25_p 3.33061e-19 $X=0.567 $Y=0.1355 $X2=0 $Y2=0
cc_120 VSS N_4_c_26_p 0.00110314f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_121 N_4_c_24_p N_19_M24_s 2.33161e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.216
cc_122 N_4_M7_g N_19_c_685_n 0.00248549f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_123 N_4_c_24_p N_19_c_685_n 0.00208457f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_124 N_4_c_29_p N_19_c_685_n 7.88525e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_125 N_4_c_24_p N_20_c_694_n 0.00250239f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_126 N_SE_M2_g N_6_M3_g 0.00304756f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_127 N_SE_c_138_p N_6_c_217_n 0.00126421f $X=0.297 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_128 N_SE_c_139_p N_6_c_218_n 2.80156e-19 $X=1.215 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_129 N_SE_c_140_p N_6_c_218_n 0.00154788f $X=1.215 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_130 N_SE_c_141_p N_6_c_218_n 2.41437e-19 $X=1.175 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_131 N_SE_c_142_p N_6_c_221_n 0.00114532f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_132 N_SE_c_141_p N_6_c_214_n 0.0681088f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_133 N_SE_c_144_p N_6_c_223_n 8.79603e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_134 N_SE_c_140_p N_6_c_224_n 0.00603469f $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_135 N_SE_c_141_p N_6_c_224_n 0.00103045f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_136 N_SE_c_147_p N_6_c_224_n 3.73635e-19 $X=1.215 $Y=0.09 $X2=0 $Y2=0
cc_137 N_SE_c_141_p N_6_c_227_n 2.46239e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_138 N_SE_c_135_n N_6_c_228_n 3.24594e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_139 N_SE_M2_g N_D_M4_g 2.13359e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_140 N_SE_c_134_n N_9_c_360_n 0.00266639f $X=0.225 $Y=0.045 $X2=0 $Y2=0
cc_141 N_SE_c_136_n N_9_c_360_n 4.45368e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_142 N_SE_c_153_p N_9_c_360_n 2.64176e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_143 N_SE_c_135_n N_9_c_348_n 8.13669e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_144 N_SE_c_136_n N_9_c_348_n 0.00228611f $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_145 N_SE_c_141_p N_9_c_365_n 0.00228611f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_146 N_SE_c_153_p N_9_c_326_n 0.00292661f $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_147 N_SE_c_158_p N_9_c_327_n 0.00266639f $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_148 N_SE_c_135_n N_9_c_355_n 0.00266639f $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_149 N_SE_c_141_p N_10_c_405_n 4.38905e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_150 N_SE_c_141_p N_10_c_417_n 3.0053e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_151 N_SE_c_141_p N_10_c_418_n 7.16568e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_152 N_SE_c_141_p N_11_c_457_n 0.00113636f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_153 N_SE_c_141_p N_11_c_477_n 2.78297e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_154 N_SE_c_141_p N_11_c_478_n 5.99401e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_155 N_SE_c_141_p N_11_c_479_n 4.8504e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_156 N_SE_c_141_p N_11_c_480_n 4.65038e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_157 N_SE_c_141_p N_12_c_523_n 5.48108e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_158 N_SE_c_141_p N_12_c_524_n 0.00109158f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_159 N_SE_c_141_p N_12_c_525_n 5.50727e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_160 N_SE_c_141_p N_12_c_526_n 9.11285e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_161 N_SE_c_141_p N_12_c_527_n 4.62125e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_162 N_SE_c_141_p N_12_c_528_n 5.48546e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_163 N_SE_M14_g N_13_M15_g 0.00268443f $X=1.215 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_164 N_SE_c_175_p N_13_c_565_n 0.00112344f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_165 N_SE_c_141_p N_13_c_556_n 2.30689e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_166 N_SE_c_141_p N_13_c_567_n 9.08574e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_167 N_SE_c_141_p N_13_c_568_n 0.00124317f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_168 N_SE_c_141_p N_13_c_569_n 4.54245e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_169 N_SE_c_141_p N_13_c_570_n 4.39544e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_170 N_SE_c_141_p N_13_c_571_n 5.37888e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_171 N_SE_c_140_p N_13_c_572_n 3.26078e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_172 N_SE_c_141_p N_13_c_573_n 9.30198e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_173 N_SE_c_139_p N_13_c_574_n 9.30198e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_174 N_SE_c_142_p N_13_c_574_n 0.00114818f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_175 N_SE_c_186_p N_13_c_576_n 0.00409247f $X=1.215 $Y=0.113 $X2=0 $Y2=0
cc_176 N_SE_c_187_p N_14_c_625_n 2.31793e-19 $X=0.261 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_177 N_SE_M2_g N_14_c_628_n 3.83731e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_178 N_SE_c_189_p N_14_c_628_n 6.51345e-19 $X=0.258 $Y=0.135 $X2=0 $Y2=0
cc_179 VSS N_SE_c_134_n 2.40719e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.135
cc_180 VSS N_SE_c_136_n 5.30841e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.135
cc_181 VSS N_SE_c_153_p 9.86432e-19 $X=0.225 $Y=0.081 $X2=0.081 $Y2=0.135
cc_182 VSS N_SE_c_144_p 0.00129447f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_183 VSS N_SE_c_136_n 7.061e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_184 VSS N_SE_c_153_p 7.68051e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_185 VSS N_SE_c_134_n 8.44602e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.15
cc_186 VSS N_SE_c_136_n 5.36527e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.15
cc_187 VSS N_SE_c_141_p 0.00141783f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_188 VSS N_SE_c_141_p 2.35788e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_189 VSS N_SE_c_136_n 6.93145e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_190 VSS N_SE_c_141_p 9.13621e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_191 VSS N_SE_c_141_p 4.6862e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_192 VSS N_SE_c_141_p 5.41611e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_193 VSS N_SE_c_141_p 8.51044e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_194 VSS N_SE_c_205_p 0.00129447f $X=0.279 $Y=0.135 $X2=0 $Y2=0
cc_195 VSS N_SE_c_136_n 3.48715e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_196 VSS N_SE_c_158_p 9.77595e-19 $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_197 VSS N_SE_c_141_p 2.40178e-19 $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.135
cc_198 VSS N_SE_c_141_p 6.42719e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_199 VSS N_SE_c_141_p 0.00110738f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_200 N_SE_c_147_p N_QN_c_675_n 3.2291e-19 $X=1.215 $Y=0.09 $X2=0.081 $Y2=0.15
cc_201 N_SE_c_140_p N_QN_c_676_n 8.07872e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_202 N_SE_c_141_p N_20_c_694_n 4.98441e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_203 N_6_M3_g N_D_M4_g 0.00304756f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_204 N_6_c_217_n N_D_c_288_n 9.71463e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_205 N_6_c_214_n D 3.33994e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_206 N_6_c_223_n D 0.00195518f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_207 N_6_c_228_n D 9.77589e-19 $X=0.351 $Y=0.126 $X2=0 $Y2=0
cc_208 N_6_M3_g N_SI_M5_g 2.48122e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_209 N_6_c_214_n SI 3.40688e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_210 N_6_c_214_n N_9_c_341_n 3.98881e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_211 N_6_c_214_n N_9_c_350_n 0.0176005f $X=0.9 $Y=0.081 $X2=0.018 $Y2=0.207
cc_212 N_6_c_223_n N_9_c_350_n 0.00113948f $X=0.351 $Y=0.135 $X2=0.018 $Y2=0.207
cc_213 N_6_c_214_n N_10_c_419_n 5.04077e-19 $X=0.9 $Y=0.081 $X2=0.945 $Y2=0.178
cc_214 N_6_c_214_n N_10_c_420_n 2.53924e-19 $X=0.9 $Y=0.081 $X2=0.945 $Y2=0.178
cc_215 N_6_c_214_n N_10_c_417_n 9.03945e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_216 N_6_c_214_n N_10_c_422_n 5.75824e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_217 N_6_c_214_n N_10_c_415_n 7.91051e-19 $X=0.9 $Y=0.081 $X2=0.018 $Y2=0.18
cc_218 N_6_c_214_n N_11_c_477_n 4.20387e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_219 N_6_c_214_n N_11_c_458_n 4.92006e-19 $X=0.9 $Y=0.081 $X2=0.071 $Y2=0.054
cc_220 N_6_c_214_n N_11_c_459_n 7.19039e-19 $X=0.9 $Y=0.081 $X2=0.056 $Y2=0.054
cc_221 N_6_c_218_n N_12_c_529_n 0.00122694f $X=1.19 $Y=0.0675 $X2=0.567
+ $Y2=0.2025
cc_222 N_6_c_248_p N_12_c_529_n 2.40393e-19 $X=1.161 $Y=0.081 $X2=0.567
+ $Y2=0.2025
cc_223 N_6_c_221_n N_12_c_531_n 4.63408e-19 $X=1.19 $Y=0.2025 $X2=0 $Y2=0
cc_224 N_6_c_248_p N_12_c_523_n 9.95523e-19 $X=1.161 $Y=0.081 $X2=0.837
+ $Y2=0.0405
cc_225 N_6_c_218_n N_12_c_524_n 9.66531e-19 $X=1.19 $Y=0.0675 $X2=0.837
+ $Y2=0.178
cc_226 N_6_c_224_n N_12_c_524_n 0.00241878f $X=1.161 $Y=0.049 $X2=0.837
+ $Y2=0.178
cc_227 N_6_c_253_p N_12_c_535_n 0.00241878f $X=1.17 $Y=0.234 $X2=0 $Y2=0
cc_228 N_6_c_248_p N_12_c_528_n 0.0012739f $X=1.161 $Y=0.081 $X2=0 $Y2=0
cc_229 N_6_c_255_p N_12_c_528_n 0.00241878f $X=1.161 $Y=0.2125 $X2=0 $Y2=0
cc_230 N_6_c_256_p N_12_c_538_n 0.00241878f $X=1.161 $Y=0.225 $X2=0 $Y2=0
cc_231 N_6_c_215_n N_13_c_568_n 6.23859e-19 $X=0.936 $Y=0.081 $X2=0 $Y2=0
cc_232 N_6_c_248_p N_13_c_571_n 3.66836e-19 $X=1.161 $Y=0.081 $X2=0 $Y2=0
cc_233 N_6_c_248_p N_13_c_559_n 5.24665e-19 $X=1.161 $Y=0.081 $X2=0 $Y2=0
cc_234 N_6_c_215_n N_13_c_562_n 3.12147e-19 $X=0.936 $Y=0.081 $X2=0.018
+ $Y2=0.225
cc_235 N_6_c_218_n N_13_c_573_n 2.31667e-19 $X=1.19 $Y=0.0675 $X2=0.027
+ $Y2=0.234
cc_236 N_6_c_262_p N_13_c_573_n 2.53206e-19 $X=1.179 $Y=0.234 $X2=0.027
+ $Y2=0.234
cc_237 N_6_c_248_p N_13_c_573_n 0.00813033f $X=1.161 $Y=0.081 $X2=0.027
+ $Y2=0.234
cc_238 N_6_c_224_n N_13_c_573_n 0.00109426f $X=1.161 $Y=0.049 $X2=0.027
+ $Y2=0.234
cc_239 N_6_c_221_n N_13_c_574_n 3.0124e-19 $X=1.19 $Y=0.2025 $X2=0.054 $Y2=0.234
cc_240 N_6_c_266_p N_13_c_574_n 2.53206e-19 $X=1.188 $Y=0.234 $X2=0.054
+ $Y2=0.234
cc_241 N_6_M3_g N_14_c_633_n 2.37298e-19 $X=0.351 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_242 VSS N_6_c_214_n 3.90811e-19 $X=0.9 $Y=0.081 $X2=0.567 $Y2=0.2025
cc_243 VSS N_6_c_227_n 7.35661e-19 $X=0.351 $Y=0.099 $X2=0.567 $Y2=0.2025
cc_244 VSS N_6_c_270_p 6.42252e-19 $X=0.351 $Y=0.081 $X2=0 $Y2=0
cc_245 VSS N_6_c_270_p 0.00369658f $X=0.351 $Y=0.081 $X2=0.837 $Y2=0.0405
cc_246 N_6_M3_g N_16_c_657_n 2.50526e-19 $X=0.351 $Y=0.0675 $X2=0.837 $Y2=0.0405
cc_247 N_6_c_223_n N_16_c_657_n 0.00110314f $X=0.351 $Y=0.135 $X2=0.837
+ $Y2=0.0405
cc_248 VSS N_6_c_227_n 2.30452e-19 $X=0.351 $Y=0.099 $X2=0.135 $Y2=0.135
cc_249 VSS N_6_c_214_n 7.92007e-19 $X=0.9 $Y=0.081 $X2=0.675 $Y2=0.0405
cc_250 VSS N_6_c_270_p 8.14481e-19 $X=0.351 $Y=0.081 $X2=0.675 $Y2=0.178
cc_251 VSS N_6_c_214_n 2.67459e-19 $X=0.9 $Y=0.081 $X2=0.675 $Y2=0.178
cc_252 VSS N_6_c_214_n 3.16736e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_253 VSS N_6_c_214_n 2.43408e-19 $X=0.9 $Y=0.081 $X2=0.837 $Y2=0.0405
cc_254 VSS N_6_c_214_n 5.19239e-19 $X=0.9 $Y=0.081 $X2=0.837 $Y2=0.178
cc_255 N_6_c_221_n N_QN_c_677_n 3.12696e-19 $X=1.19 $Y=0.2025 $X2=0.567
+ $Y2=0.1355
cc_256 N_6_c_218_n N_QN_c_678_n 3.35016e-19 $X=1.19 $Y=0.0675 $X2=0.675
+ $Y2=0.178
cc_257 N_6_c_266_p N_QN_c_679_n 2.64332e-19 $X=1.188 $Y=0.234 $X2=0.945
+ $Y2=0.2295
cc_258 N_6_c_215_n N_20_c_694_n 5.02041e-19 $X=0.936 $Y=0.081 $X2=0.567
+ $Y2=0.1355
cc_259 VSS N_6_c_270_p 2.73492e-19 $X=0.351 $Y=0.081 $X2=0.135 $Y2=0.054
cc_260 N_D_M4_g N_SI_M5_g 0.00348334f $X=0.405 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_261 D SI 7.00288e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_262 N_D_c_288_n N_SI_c_309_n 0.00109838f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_263 D N_9_c_350_n 0.00102191f $X=0.405 $Y=0.134 $X2=0.018 $Y2=0.207
cc_264 N_D_M4_g N_14_c_633_n 2.37298e-19 $X=0.405 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_265 VSS N_D_M4_g 3.08888e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_266 VSS D 5.77345e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_267 N_D_M4_g N_16_c_660_n 2.43567e-19 $X=0.405 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_268 D N_16_c_660_n 0.00108212f $X=0.405 $Y=0.134 $X2=0.837 $Y2=0.178
cc_269 D N_16_c_661_n 3.4434e-19 $X=0.405 $Y=0.134 $X2=0.837 $Y2=0.178
cc_270 VSS D 8.86227e-19 $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.135
cc_271 VSS D 0.00161923f $X=0.405 $Y=0.134 $X2=0.675 $Y2=0.178
cc_272 SI N_9_c_350_n 0.00138386f $X=0.473 $Y=0.135 $X2=0.018 $Y2=0.207
cc_273 SI N_14_c_626_n 0.00560919f $X=0.473 $Y=0.135 $X2=0 $Y2=0
cc_274 SI N_14_c_636_n 0.00167456f $X=0.473 $Y=0.135 $X2=0.837 $Y2=0.0405
cc_275 N_SI_M5_g N_14_c_629_n 2.70361e-19 $X=0.459 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_276 SI N_16_c_655_n 6.69571e-19 $X=0.473 $Y=0.135 $X2=0.675 $Y2=0.178
cc_277 VSS N_SI_M5_g 3.10987e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_278 VSS N_SI_c_309_n 2.08525e-19 $X=0.475 $Y=0.135 $X2=0 $Y2=0
cc_279 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.837 $Y2=0.0405
cc_280 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.837 $Y2=0.0405
cc_281 VSS SI 0.00110314f $X=0.473 $Y=0.135 $X2=0 $Y2=0
cc_282 N_9_M6_g N_10_M8_g 2.82885e-19 $X=0.621 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_283 N_9_c_349_n N_10_c_425_n 2.61213e-19 $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_284 N_9_c_365_n N_10_c_425_n 2.61213e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_285 N_9_c_354_n N_10_c_410_n 0.00318254f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_286 N_9_c_349_n N_10_c_411_n 0.00128311f $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_287 N_9_M11_g N_11_M9_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_288 N_9_c_333_n N_11_c_485_n 3.1781e-19 $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.135
cc_289 N_9_c_345_n N_11_c_453_n 3.24488e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_290 N_9_M6_g N_11_c_487_n 3.41974e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_291 N_9_c_345_n N_11_c_487_n 0.00102727f $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_292 N_9_c_341_n N_11_c_489_n 0.00133858f $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_293 N_9_c_350_n N_11_c_490_n 7.726e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_294 N_9_c_345_n N_11_c_460_n 8.63476e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_295 N_9_c_350_n N_11_c_460_n 5.92766e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_296 N_9_c_365_n N_11_c_471_n 3.86765e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_297 N_9_c_350_n N_11_c_472_n 3.86765e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_298 N_9_M11_g N_12_M12_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_299 N_9_M11_g N_13_c_569_n 3.18506e-19 $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_300 N_9_c_354_n N_13_c_569_n 4.09234e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_301 N_9_c_354_n N_13_c_589_n 0.00320381f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_302 N_9_c_354_n N_13_c_563_n 3.56772e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_303 N_9_c_349_n N_13_c_573_n 9.40125e-19 $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_304 N_9_c_334_n N_14_c_625_n 0.0010034f $X=0.16 $Y=0.216 $X2=0.081 $Y2=0.135
cc_305 N_9_c_343_n N_14_c_625_n 0.00105265f $X=0.189 $Y=0.153 $X2=0.081
+ $Y2=0.135
cc_306 N_9_c_350_n N_14_c_626_n 4.24134e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_307 N_9_c_336_n N_14_c_628_n 7.83928e-19 $X=0.18 $Y=0.234 $X2=0 $Y2=0
cc_308 VSS N_9_c_400_p 9.30745e-19 $X=0.16 $Y=0.054 $X2=0.081 $Y2=0.135
cc_309 N_10_M8_g N_11_M9_g 0.00268443f $X=0.729 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_310 N_10_c_417_n N_11_M9_g 3.80603e-19 $X=0.797 $Y=0.09 $X2=0.135 $Y2=0.054
cc_311 N_10_c_418_n N_11_c_480_n 2.46574e-19 $X=0.81 $Y=0.054 $X2=0 $Y2=0
cc_312 N_10_c_419_n N_11_c_498_n 0.00360624f $X=0.747 $Y=0.09 $X2=0 $Y2=0
cc_313 N_10_c_420_n N_11_c_458_n 3.99428e-19 $X=0.747 $Y=0.09 $X2=0.071
+ $Y2=0.054
cc_314 N_10_c_411_n N_11_c_490_n 2.22221e-19 $X=0.837 $Y=0.165 $X2=0.056
+ $Y2=0.216
cc_315 N_10_c_435_p N_11_c_466_n 2.22221e-19 $X=0.837 $Y=0.225 $X2=0.018
+ $Y2=0.045
cc_316 N_10_c_417_n N_11_c_471_n 0.00219679f $X=0.797 $Y=0.09 $X2=0.018
+ $Y2=0.198
cc_317 N_10_c_437_p N_11_c_471_n 9.66928e-19 $X=0.837 $Y=0.14 $X2=0.018
+ $Y2=0.198
cc_318 N_10_M8_g N_11_c_473_n 3.21351e-19 $X=0.729 $Y=0.0405 $X2=0.018 $Y2=0.216
cc_319 N_10_c_419_n N_11_c_473_n 0.00219679f $X=0.747 $Y=0.09 $X2=0.018
+ $Y2=0.216
cc_320 N_10_c_405_n N_13_c_556_n 0.00379158f $X=0.81 $Y=0.0405 $X2=0.837
+ $Y2=0.0405
cc_321 N_10_c_418_n N_13_c_556_n 2.84891e-19 $X=0.81 $Y=0.054 $X2=0.837
+ $Y2=0.0405
cc_322 N_10_c_415_n N_13_c_556_n 2.08929e-19 $X=0.837 $Y=0.09 $X2=0.837
+ $Y2=0.0405
cc_323 N_10_c_408_n N_13_c_558_n 0.00222825f $X=0.866 $Y=0.2295 $X2=0 $Y2=0
cc_324 N_10_c_405_n N_13_c_568_n 3.41768e-19 $X=0.81 $Y=0.0405 $X2=0 $Y2=0
cc_325 N_10_c_415_n N_13_c_559_n 4.2911e-19 $X=0.837 $Y=0.09 $X2=0 $Y2=0
cc_326 N_10_c_413_n N_13_c_561_n 4.2911e-19 $X=0.837 $Y=0.207 $X2=0 $Y2=0
cc_327 N_10_c_408_n N_13_c_562_n 3.64454e-19 $X=0.866 $Y=0.2295 $X2=0.018
+ $Y2=0.225
cc_328 N_10_c_448_p N_13_c_562_n 4.86017e-19 $X=0.828 $Y=0.234 $X2=0.018
+ $Y2=0.225
cc_329 N_10_c_449_p N_13_c_563_n 4.2911e-19 $X=0.837 $Y=0.101 $X2=0.054
+ $Y2=0.036
cc_330 N_11_c_453_n N_14_c_626_n 0.00424458f $X=0.594 $Y=0.2025 $X2=0 $Y2=0
cc_331 N_11_c_455_n N_14_c_626_n 4.3429e-19 $X=0.595 $Y=0.234 $X2=0 $Y2=0
cc_332 N_11_c_455_n N_14_c_636_n 2.8677e-19 $X=0.595 $Y=0.234 $X2=0.837
+ $Y2=0.0405
cc_333 VSS N_11_c_453_n 0.0016174f $X=0.594 $Y=0.2025 $X2=0.567 $Y2=0.1355
cc_334 VSS N_11_c_477_n 0.00414127f $X=0.648 $Y=0.036 $X2=0.567 $Y2=0.1355
cc_335 VSS N_11_c_478_n 3.30384e-19 $X=0.649 $Y=0.036 $X2=0.567 $Y2=0.1355
cc_336 VSS N_11_c_477_n 2.79363e-19 $X=0.648 $Y=0.036 $X2=0.675 $Y2=0.0405
cc_337 VSS N_11_c_458_n 2.70508e-19 $X=0.693 $Y=0.081 $X2=0.675 $Y2=0.0405
cc_338 N_11_c_453_n N_19_c_685_n 0.00167238f $X=0.594 $Y=0.2025 $X2=0.567
+ $Y2=0.1355
cc_339 N_11_c_515_p N_19_c_685_n 0.00315491f $X=0.684 $Y=0.234 $X2=0.567
+ $Y2=0.1355
cc_340 N_11_c_487_n N_19_c_685_n 0.00111131f $X=0.649 $Y=0.234 $X2=0.567
+ $Y2=0.1355
cc_341 N_11_c_477_n N_19_c_685_n 5.67227e-19 $X=0.648 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_342 N_11_c_518_p N_19_c_685_n 4.0515e-19 $X=0.693 $Y=0.225 $X2=0.567
+ $Y2=0.1355
cc_343 N_11_c_519_p N_19_c_685_n 0.0409693f $X=0.693 $Y=0.216 $X2=0.567
+ $Y2=0.1355
cc_344 N_11_c_457_n N_22_M8_s 2.44135e-19 $X=0.684 $Y=0.036 $X2=0.135 $Y2=0.054
cc_345 N_11_c_480_n N_22_M8_s 3.62465e-19 $X=0.693 $Y=0.062 $X2=0.135 $Y2=0.054
cc_346 N_12_M12_g N_13_M13_g 0.00268443f $X=0.999 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_347 N_12_c_527_n N_13_M13_g 3.55314e-19 $X=1.062 $Y=0.036 $X2=0.135 $Y2=0.054
cc_348 N_12_c_525_n N_13_c_567_n 0.00136796f $X=1.008 $Y=0.036 $X2=0.945
+ $Y2=0.178
cc_349 N_12_c_523_n N_13_c_571_n 0.00136796f $X=0.999 $Y=0.105 $X2=0 $Y2=0
cc_350 N_12_c_544_p N_13_c_559_n 3.34766e-19 $X=0.999 $Y=0.1055 $X2=0 $Y2=0
cc_351 N_12_c_523_n N_13_c_559_n 0.00136796f $X=0.999 $Y=0.105 $X2=0 $Y2=0
cc_352 N_12_c_535_n N_13_c_561_n 5.28703e-19 $X=1.107 $Y=0.225 $X2=0 $Y2=0
cc_353 N_12_M12_g N_13_c_609_n 6.35734e-19 $X=0.999 $Y=0.0405 $X2=0 $Y2=0
cc_354 N_12_c_523_n N_13_c_609_n 7.99759e-19 $X=0.999 $Y=0.105 $X2=0 $Y2=0
cc_355 N_12_c_527_n N_13_c_611_n 2.75024e-19 $X=1.062 $Y=0.036 $X2=0.071
+ $Y2=0.216
cc_356 N_12_c_538_n N_13_c_611_n 0.00266503f $X=1.107 $Y=0.171 $X2=0.071
+ $Y2=0.216
cc_357 N_12_c_531_n N_13_c_573_n 2.19627e-19 $X=1.078 $Y=0.2295 $X2=0.027
+ $Y2=0.234
cc_358 N_12_c_538_n N_13_c_573_n 0.00106087f $X=1.107 $Y=0.171 $X2=0.027
+ $Y2=0.234
cc_359 N_12_c_553_p N_13_c_573_n 5.80975e-19 $X=1.098 $Y=0.234 $X2=0.027
+ $Y2=0.234
cc_360 N_12_c_525_n N_20_c_694_n 5.06067e-19 $X=1.008 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_361 N_13_c_576_n N_QN_c_677_n 0.00114532f $X=1.269 $Y=0.136 $X2=0.567
+ $Y2=0.1355
cc_362 N_13_c_572_n N_QN_c_681_n 2.31819e-19 $X=1.269 $Y=0.153 $X2=0.675
+ $Y2=0.0405
cc_363 N_13_c_576_n N_QN_c_681_n 0.00431194f $X=1.269 $Y=0.136 $X2=0.675
+ $Y2=0.0405
cc_364 N_13_c_576_n N_QN_c_678_n 5.42522e-19 $X=1.269 $Y=0.136 $X2=0.675
+ $Y2=0.178
cc_365 N_13_c_556_n N_20_c_694_n 0.00210698f $X=0.864 $Y=0.0405 $X2=0.567
+ $Y2=0.1355
cc_366 N_13_c_567_n N_20_c_694_n 0.00203632f $X=0.936 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_367 N_13_c_570_n N_20_c_694_n 0.00129774f $X=0.92 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_368 N_13_c_571_n N_20_c_694_n 0.00104094f $X=0.945 $Y=0.081 $X2=0.567
+ $Y2=0.1355
cc_369 N_13_c_624_p N_20_c_694_n 2.5109e-19 $X=0.99 $Y=0.162 $X2=0.567
+ $Y2=0.1355
cc_370 VSS N_14_c_625_n 0.00156967f $X=0.272 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_371 VSS N_14_c_626_n 0.00145872f $X=0.542 $Y=0.2025 $X2=0.675 $Y2=0.178
cc_372 N_14_c_625_n N_16_c_668_n 0.003872f $X=0.272 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_373 N_14_c_633_n N_16_c_668_n 0.00248801f $X=0.447 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_374 N_14_c_626_n N_16_c_670_n 0.00434154f $X=0.542 $Y=0.2025 $X2=0.567
+ $Y2=0.1355
cc_375 N_14_c_633_n N_16_c_670_n 0.0025506f $X=0.447 $Y=0.234 $X2=0.567
+ $Y2=0.1355
cc_376 N_14_c_625_n N_16_c_654_n 3.19827e-19 $X=0.272 $Y=0.2025 $X2=0.567
+ $Y2=0.2025
cc_377 N_14_c_633_n N_16_c_654_n 0.0113176f $X=0.447 $Y=0.234 $X2=0.567
+ $Y2=0.2025
cc_378 VSS N_14_c_626_n 4.53012e-19 $X=0.542 $Y=0.2025 $X2=0.837 $Y2=0.178
cc_379 VSS N_16_c_670_n 0.00141703f $X=0.432 $Y=0.2025 $X2=0.135 $Y2=0.135

* END of "./SDFLx1_ASAP7_75t_SRAM.pex.sp.SDFLX1_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: SDFLx2_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 13:04:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "SDFLx2_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./SDFLx2_ASAP7_75t_SRAM.pex.sp.pex"
* File: SDFLx2_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 13:04:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_SDFLX2_ASAP7_75T_SRAM%CLK 2 5 7 11 16 VSS
c12 11 VSS 0.00713456f $X=0.081 $Y=0.135
c13 5 VSS 0.00188964f $X=0.081 $Y=0.135
c14 2 VSS 0.0628473f $X=0.081 $Y=0.054
r15 11 16 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.15
r16 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%4 2 5 7 10 13 16 19 22 25 28 31 45 48 50 57 58 65
+ 72 79 83 86 90 97 100 101 102 104 123 VSS
c122 134 VSS 7.0154e-20 $X=0.03 $Y=0.189
c123 133 VSS 5.9624e-19 $X=0.027 $Y=0.189
c124 123 VSS 6.49238e-19 $X=0.729 $Y=0.18
c125 104 VSS 0.00976003f $X=0.729 $Y=0.189
c126 102 VSS 0.00542037f $X=0.371 $Y=0.189
c127 101 VSS 0.00609885f $X=0.175 $Y=0.189
c128 100 VSS 0.0013748f $X=0.567 $Y=0.189
c129 97 VSS 0.00291011f $X=0.135 $Y=0.189
c130 93 VSS 5.52785e-19 $X=0.033 $Y=0.189
c131 90 VSS 9.61695e-20 $X=0.567 $Y=0.18
c132 86 VSS 5.76385e-19 $X=0.567 $Y=0.135
c133 83 VSS 1.05495e-19 $X=0.135 $Y=0.18
c134 79 VSS 6.50523e-19 $X=0.135 $Y=0.135
c135 75 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c136 74 VSS 0.00169428f $X=0.047 $Y=0.234
c137 72 VSS 0.0024557f $X=0.054 $Y=0.234
c138 70 VSS 0.00306385f $X=0.027 $Y=0.234
c139 68 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c140 67 VSS 0.00205521f $X=0.047 $Y=0.036
c141 65 VSS 0.00239525f $X=0.054 $Y=0.036
c142 63 VSS 0.00305101f $X=0.027 $Y=0.036
c143 62 VSS 3.84318e-19 $X=0.018 $Y=0.216
c144 61 VSS 3.30259e-19 $X=0.018 $Y=0.207
c145 60 VSS 3.64183e-19 $X=0.018 $Y=0.225
c146 58 VSS 0.0039492f $X=0.018 $Y=0.164
c147 57 VSS 0.00142827f $X=0.018 $Y=0.081
c148 56 VSS 8.21418e-19 $X=0.018 $Y=0.18
c149 53 VSS 0.00514186f $X=0.056 $Y=0.216
c150 50 VSS 2.98509e-19 $X=0.071 $Y=0.216
c151 48 VSS 0.00458629f $X=0.056 $Y=0.054
c152 45 VSS 2.98509e-19 $X=0.071 $Y=0.054
c153 28 VSS 0.108836f $X=0.945 $Y=0.178
c154 25 VSS 1.08457e-19 $X=0.837 $Y=0.178
c155 22 VSS 0.0600244f $X=0.837 $Y=0.0405
c156 19 VSS 2.24613e-19 $X=0.675 $Y=0.178
c157 16 VSS 0.0602569f $X=0.675 $Y=0.0405
c158 10 VSS 0.0660345f $X=0.567 $Y=0.1355
c159 5 VSS 0.00179729f $X=0.135 $Y=0.135
c160 2 VSS 0.0627664f $X=0.135 $Y=0.054
r161 133 134 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.03 $Y2=0.189
r162 130 133 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.027 $Y2=0.189
r163 122 123 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.729 $Y=0.18
+ $X2=0.729 $Y2=0.18
r164 104 123 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.729 $Y=0.189 $X2=0.729
+ $Y2=0.189
r165 101 102 13.3086 $w=1.8e-08 $l=1.96e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.175 $Y=0.189 $X2=0.371 $Y2=0.189
r166 99 104 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.729 $Y2=0.189
r167 99 102 13.3086 $w=1.8e-08 $l=1.96e-07 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.371 $Y2=0.189
r168 99 100 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.567 $Y=0.189 $X2=0.567
+ $Y2=0.189
r169 96 101 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.175 $Y2=0.189
r170 96 97 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.135 $Y=0.189 $X2=0.135
+ $Y2=0.189
r171 93 134 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.03 $Y2=0.189
r172 92 96 6.92593 $w=1.8e-08 $l=1.02e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.135 $Y2=0.189
r173 92 93 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.189 $X2=0.033
+ $Y2=0.189
r174 90 100 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.18 $X2=0.567 $Y2=0.189
r175 89 90 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.171 $X2=0.567 $Y2=0.18
r176 86 89 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.171
r177 83 97 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.18 $X2=0.135 $Y2=0.189
r178 82 83 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.164 $X2=0.135 $Y2=0.18
r179 79 82 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.164
r180 74 75 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r181 72 75 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r182 70 74 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r183 67 68 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r184 65 68 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r185 63 67 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r186 61 62 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.207 $X2=0.018 $Y2=0.216
r187 60 70 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r188 60 62 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.216
r189 59 130 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.189
r190 59 61 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.207
r191 57 58 5.6358 $w=1.8e-08 $l=8.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.164
r192 56 130 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.189
r193 56 58 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.164
r194 55 63 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r195 55 57 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r196 53 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r197 50 53 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r198 48 65 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r199 45 48 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r200 28 31 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.178 $X2=0.945 $Y2=0.2295
r201 25 28 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08 $X=0.837
+ $Y=0.178 $X2=0.945 $Y2=0.178
r202 25 122 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.837 $Y=0.178 $X2=0.729 $Y2=0.178
r203 22 25 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0405 $X2=0.837 $Y2=0.178
r204 19 122 43.022 $w=2.6e-08 $l=5.4e-08 $layer=LISD $thickness=2.8e-08 $X=0.675
+ $Y=0.178 $X2=0.729 $Y2=0.178
r205 16 19 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.178
r206 10 86 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r207 10 13 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1355 $X2=0.567 $Y2=0.2025
r208 5 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r209 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r210 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%SE 2 5 7 10 13 15 19 22 23 24 31 33 41 44 45 46 47
+ 54 58 59 62 63 VSS
c80 63 VSS 5.91978e-19 $X=1.215 $Y=0.113
c81 62 VSS 0.00217892f $X=1.215 $Y=0.09
c82 59 VSS 2.63823e-19 $X=0.225 $Y=0.099
c83 58 VSS 5.90201e-19 $X=0.225 $Y=0.081
c84 54 VSS 0.00209141f $X=1.215 $Y=0.136
c85 47 VSS 0.0381258f $X=1.175 $Y=0.045
c86 46 VSS 0.00642311f $X=0.337 $Y=0.045
c87 45 VSS 0.00700109f $X=1.215 $Y=0.045
c88 44 VSS 0.0031469f $X=1.215 $Y=0.045
c89 41 VSS 0.00531f $X=0.225 $Y=0.045
c90 31 VSS 0.00110873f $X=0.225 $Y=0.126
c91 24 VSS 2.51525e-19 $X=0.279 $Y=0.135
c92 23 VSS 1.48251e-19 $X=0.261 $Y=0.135
c93 22 VSS 6.38823e-20 $X=0.258 $Y=0.135
c94 21 VSS 0.00134071f $X=0.255 $Y=0.135
c95 19 VSS 6.89032e-19 $X=0.297 $Y=0.135
c96 13 VSS 0.0019468f $X=1.215 $Y=0.136
c97 10 VSS 0.0611074f $X=1.215 $Y=0.0675
c98 5 VSS 0.0031928f $X=0.297 $Y=0.135
c99 2 VSS 0.063344f $X=0.297 $Y=0.0675
r100 62 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.09 $X2=1.215 $Y2=0.113
r101 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.081 $X2=0.225 $Y2=0.099
r102 54 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.136 $X2=1.215 $Y2=0.113
r103 46 47 56.9012 $w=1.8e-08 $l=8.38e-07 $layer=M2 $thickness=3.6e-08 $X=0.337
+ $Y=0.045 $X2=1.175 $Y2=0.045
r104 45 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.215 $Y2=0.09
r105 44 47 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.175 $Y2=0.045
r106 44 45 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.215 $Y=0.045 $X2=1.215
+ $Y2=0.045
r107 41 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.081
r108 40 46 7.60494 $w=1.8e-08 $l=1.12e-07 $layer=M2 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.337 $Y2=0.045
r109 40 41 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.225 $Y=0.045 $X2=0.225
+ $Y2=0.045
r110 31 59 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.099
r111 31 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r112 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.135 $X2=0.279 $Y2=0.135
r113 22 23 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.258
+ $Y=0.135 $X2=0.261 $Y2=0.135
r114 21 22 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.255
+ $Y=0.135 $X2=0.258 $Y2=0.135
r115 19 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.279 $Y2=0.135
r116 17 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.225 $Y2=0.135
r117 17 21 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.255 $Y2=0.135
r118 13 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.215 $Y=0.136 $X2=1.215
+ $Y2=0.136
r119 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.136 $X2=1.215 $Y2=0.2025
r120 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.0675 $X2=1.215 $Y2=0.136
r121 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r122 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r123 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%6 2 5 7 9 12 14 17 23 26 28 29 33 36 38 39 43 51
+ 57 58 65 VSS
c72 65 VSS 8.50758e-20 $X=1.161 $Y=0.2125
c73 58 VSS 5.45782e-19 $X=0.351 $Y=0.126
c74 57 VSS 8.0335e-19 $X=0.351 $Y=0.099
c75 51 VSS 0.00278401f $X=1.161 $Y=0.049
c76 43 VSS 3.76741e-19 $X=0.351 $Y=0.135
c77 39 VSS 9.89222e-19 $X=0.936 $Y=0.081
c78 38 VSS 0.00685031f $X=0.9 $Y=0.081
c79 36 VSS 0.00203618f $X=1.161 $Y=0.081
c80 33 VSS 8.1122e-19 $X=0.351 $Y=0.081
c81 29 VSS 6.98259e-19 $X=1.179 $Y=0.234
c82 28 VSS 0.00240687f $X=1.17 $Y=0.234
c83 26 VSS 0.00313492f $X=1.188 $Y=0.234
c84 23 VSS 2.83663e-20 $X=1.161 $Y=0.225
c85 17 VSS 0.00673327f $X=1.19 $Y=0.2025
c86 14 VSS 3.02808e-19 $X=1.205 $Y=0.2025
c87 12 VSS 0.0657106f $X=1.19 $Y=0.0675
c88 9 VSS 3.25039e-19 $X=1.205 $Y=0.0675
c89 5 VSS 0.00125227f $X=0.351 $Y=0.135
c90 2 VSS 0.0585837f $X=0.351 $Y=0.0675
r91 64 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.2 $X2=1.161 $Y2=0.2125
r92 57 58 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.099 $X2=0.351 $Y2=0.126
r93 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.161 $Y=0.049 $X2=1.161
+ $Y2=0.049
r94 43 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.126
r95 38 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.9
+ $Y=0.081 $X2=0.936 $Y2=0.081
r96 37 64 8.08025 $w=1.8e-08 $l=1.19e-07 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.2
r97 37 51 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.049
r98 36 39 15.2778 $w=1.8e-08 $l=2.25e-07 $layer=M2 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=0.936 $Y2=0.081
r99 36 37 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.161 $Y=0.081 $X2=1.161
+ $Y2=0.081
r100 33 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.099
r101 32 38 37.2778 $w=1.8e-08 $l=5.49e-07 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.9 $Y2=0.081
r102 32 33 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.081 $X2=0.351
+ $Y2=0.081
r103 28 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.17
+ $Y=0.234 $X2=1.179 $Y2=0.234
r104 26 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.188
+ $Y=0.234 $X2=1.179 $Y2=0.234
r105 23 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.225 $X2=1.161 $Y2=0.2125
r106 22 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.17 $Y2=0.234
r107 22 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.161 $Y2=0.225
r108 17 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.188 $Y=0.234
+ $X2=1.188 $Y2=0.234
r109 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.2025 $X2=1.19 $Y2=0.2025
r110 12 50 7.35229 $w=8.1e-08 $l=2.9e-08 $layer=LISD $thickness=2.8e-08 $X=1.19
+ $Y=0.0675 $X2=1.161 $Y2=0.0675
r111 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.0675 $X2=1.19 $Y2=0.0675
r112 5 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r113 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r114 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%D 2 5 7 11 VSS
c18 11 VSS 0.00145113f $X=0.405 $Y=0.134
c19 5 VSS 0.00106786f $X=0.405 $Y=0.135
c20 2 VSS 0.0589243f $X=0.405 $Y=0.0675
r21 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%SI 2 7 11 14 VSS
c21 14 VSS 0.00329293f $X=0.475 $Y=0.135
c22 11 VSS 0.00333153f $X=0.473 $Y=0.135
c23 2 VSS 0.0640988f $X=0.459 $Y=0.0675
r24 11 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.475 $Y=0.135 $X2=0.475
+ $Y2=0.135
r25 5 14 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.475 $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%9 2 5 7 10 13 15 17 20 22 25 27 29 36 43 45 51 55
+ 56 57 59 61 62 69 79 80 81 82 84 85 VSS
c75 86 VSS 5.63033e-20 $X=0.189 $Y=0.216
c76 85 VSS 4.28571e-19 $X=0.189 $Y=0.207
c77 84 VSS 4.04265e-19 $X=0.189 $Y=0.189
c78 82 VSS 2.19344e-19 $X=0.189 $Y=0.1485
c79 81 VSS 3.0092e-19 $X=0.189 $Y=0.144
c80 80 VSS 4.92067e-19 $X=0.189 $Y=0.121
c81 79 VSS 8.32677e-19 $X=0.189 $Y=0.099
c82 69 VSS 0.001222f $X=0.891 $Y=0.135
c83 62 VSS 0.00209834f $X=0.817 $Y=0.153
c84 61 VSS 0.00277455f $X=0.743 $Y=0.153
c85 59 VSS 0.00277965f $X=0.891 $Y=0.153
c86 57 VSS 0.00120333f $X=0.337 $Y=0.153
c87 56 VSS 0.00116325f $X=0.211 $Y=0.153
c88 55 VSS 9.40943e-19 $X=0.621 $Y=0.153
c89 51 VSS 5.62309e-19 $X=0.189 $Y=0.153
c90 48 VSS 5.43917e-20 $X=0.189 $Y=0.225
c91 45 VSS 0.00373046f $X=0.18 $Y=0.036
c92 43 VSS 0.00194932f $X=0.189 $Y=0.036
c93 36 VSS 5.26559e-19 $X=0.621 $Y=0.135
c94 29 VSS 0.00311772f $X=0.162 $Y=0.234
c95 27 VSS 0.00522825f $X=0.18 $Y=0.234
c96 25 VSS 0.00583113f $X=0.16 $Y=0.216
c97 20 VSS 0.00576958f $X=0.16 $Y=0.054
c98 13 VSS 0.00216055f $X=0.891 $Y=0.135
c99 10 VSS 0.0585656f $X=0.891 $Y=0.0405
c100 5 VSS 0.00201785f $X=0.621 $Y=0.135
c101 2 VSS 0.0601628f $X=0.621 $Y=0.0675
r102 85 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.207 $X2=0.189 $Y2=0.216
r103 84 85 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.207
r104 83 84 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.189
r105 81 82 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.1485
r106 80 81 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.121 $X2=0.189 $Y2=0.144
r107 79 80 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.099 $X2=0.189 $Y2=0.121
r108 61 62 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.743
+ $Y=0.153 $X2=0.817 $Y2=0.153
r109 59 62 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.817 $Y2=0.153
r110 59 69 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r111 56 57 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.211
+ $Y=0.153 $X2=0.337 $Y2=0.153
r112 54 61 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.743 $Y2=0.153
r113 54 57 19.284 $w=1.8e-08 $l=2.84e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.337 $Y2=0.153
r114 54 55 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.621 $Y=0.153 $X2=0.621
+ $Y2=0.153
r115 51 83 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.164
r116 51 82 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.1485
r117 50 56 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.211 $Y2=0.153
r118 50 51 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.153 $X2=0.189
+ $Y2=0.153
r119 48 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.216
r120 45 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r121 44 79 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.099
r122 43 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r123 43 44 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r124 40 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r125 36 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.153
r126 27 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.234 $X2=0.189 $Y2=0.225
r127 27 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.162 $Y2=0.234
r128 25 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r129 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r130 20 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r131 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r132 13 69 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.135 $X2=0.891
+ $Y2=0.135
r133 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.135 $X2=0.891 $Y2=0.2295
r134 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.0405 $X2=0.891 $Y2=0.135
r135 5 36 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r136 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2295
r137 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%10 2 7 9 10 13 14 17 19 22 27 28 29 31 36 38 44 45
+ 46 47 48 49 50 54 VSS
c49 56 VSS 5.19568e-19 $X=0.828 $Y=0.09
c50 55 VSS 4.09996e-19 $X=0.819 $Y=0.09
c51 54 VSS 4.29e-19 $X=0.837 $Y=0.09
c52 50 VSS 5.92996e-19 $X=0.837 $Y=0.207
c53 49 VSS 1.19762e-19 $X=0.837 $Y=0.167
c54 48 VSS 1.59501e-19 $X=0.837 $Y=0.165
c55 47 VSS 3.13056e-19 $X=0.837 $Y=0.14
c56 46 VSS 5.61414e-19 $X=0.837 $Y=0.122
c57 45 VSS 1.91116e-19 $X=0.837 $Y=0.101
c58 44 VSS 4.02479e-19 $X=0.837 $Y=0.225
c59 42 VSS 3.58124e-20 $X=0.81 $Y=0.0715
c60 38 VSS 0.00112276f $X=0.81 $Y=0.054
c61 31 VSS 0.00670205f $X=0.828 $Y=0.234
c62 30 VSS 4.74851e-19 $X=0.7965 $Y=0.09
c63 29 VSS 0.00125276f $X=0.792 $Y=0.09
c64 28 VSS 0.00410211f $X=0.747 $Y=0.09
c65 27 VSS 4.49532e-19 $X=0.747 $Y=0.09
c66 24 VSS 1.65079e-19 $X=0.801 $Y=0.09
c67 22 VSS 0.0178177f $X=0.866 $Y=0.2295
c68 19 VSS 3.14771e-19 $X=0.881 $Y=0.2295
c69 17 VSS 2.67274e-19 $X=0.808 $Y=0.2295
c70 13 VSS 0.020153f $X=0.81 $Y=0.0405
c71 9 VSS 6.29543e-19 $X=0.827 $Y=0.0405
c72 2 VSS 0.0580179f $X=0.729 $Y=0.0405
r73 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.819
+ $Y=0.09 $X2=0.828 $Y2=0.09
r74 54 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.09 $X2=0.828 $Y2=0.09
r75 53 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.09 $X2=0.819 $Y2=0.09
r76 49 50 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.167 $X2=0.837 $Y2=0.207
r77 48 49 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.165 $X2=0.837 $Y2=0.167
r78 47 48 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.14 $X2=0.837 $Y2=0.165
r79 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.122 $X2=0.837 $Y2=0.14
r80 45 46 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.101 $X2=0.837 $Y2=0.122
r81 44 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.207
r82 43 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.09
r83 43 45 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.101
r84 41 42 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.062 $X2=0.81 $Y2=0.0715
r85 38 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.054 $X2=0.81 $Y2=0.062
r86 36 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.09
r87 36 42 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.0715
r88 31 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r89 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.81 $Y2=0.234
r90 29 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.09 $X2=0.7965 $Y2=0.09
r91 27 29 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.09 $X2=0.792 $Y2=0.09
r92 27 28 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.747 $Y=0.09 $X2=0.747
+ $Y2=0.09
r93 24 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.81 $Y2=0.09
r94 24 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.7965 $Y2=0.09
r95 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2295 $X2=0.866 $Y2=0.2295
r96 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.808
+ $Y=0.2295 $X2=0.866 $Y2=0.2295
r97 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.234 $X2=0.81
+ $Y2=0.234
r98 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2295 $X2=0.808 $Y2=0.2295
r99 13 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.054 $X2=0.81
+ $Y2=0.054
r100 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.0405 $X2=0.81 $Y2=0.0405
r101 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.0405 $X2=0.81 $Y2=0.0405
r102 5 28 16.3636 $w=2.2e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.09 $X2=0.747 $Y2=0.09
r103 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.09 $X2=0.729 $Y2=0.2295
r104 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0405 $X2=0.729 $Y2=0.09
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%11 2 5 7 9 14 17 21 22 25 30 31 33 34 37 39 40 43
+ 44 45 46 48 50 51 52 53 54 55 56 59 61 62 64 VSS
c72 64 VSS 1.00092e-19 $X=0.693 $Y=0.131
c73 61 VSS 9.09188e-19 $X=0.72 $Y=0.131
c74 59 VSS 6.42979e-19 $X=0.783 $Y=0.131
c75 56 VSS 1.82087e-19 $X=0.693 $Y=0.216
c76 55 VSS 1.40959e-19 $X=0.693 $Y=0.207
c77 54 VSS 1.07888e-19 $X=0.693 $Y=0.189
c78 53 VSS 1.66071e-19 $X=0.693 $Y=0.171
c79 52 VSS 2.71272e-19 $X=0.693 $Y=0.165
c80 51 VSS 3.53682e-19 $X=0.693 $Y=0.153
c81 50 VSS 2.11704e-19 $X=0.693 $Y=0.225
c82 48 VSS 4.15228e-19 $X=0.693 $Y=0.114
c83 47 VSS 2.7378e-19 $X=0.693 $Y=0.106
c84 46 VSS 5.46003e-20 $X=0.693 $Y=0.099
c85 45 VSS 5.96385e-20 $X=0.693 $Y=0.081
c86 43 VSS 1.65771e-19 $X=0.693 $Y=0.062
c87 42 VSS 2.30403e-19 $X=0.693 $Y=0.122
c88 40 VSS 0.00145015f $X=0.6665 $Y=0.036
c89 39 VSS 0.00201121f $X=0.649 $Y=0.036
c90 37 VSS 0.00303728f $X=0.648 $Y=0.036
c91 34 VSS 0.00412969f $X=0.684 $Y=0.036
c92 33 VSS 0.00297725f $X=0.649 $Y=0.234
c93 32 VSS 2.2805e-19 $X=0.612 $Y=0.234
c94 31 VSS 0.00126734f $X=0.609 $Y=0.234
c95 30 VSS 0.0016591f $X=0.595 $Y=0.234
c96 25 VSS 0.00558865f $X=0.684 $Y=0.234
c97 24 VSS 5.62656e-19 $X=0.594 $Y=0.2295
c98 21 VSS 0.00254121f $X=0.594 $Y=0.2025
c99 18 VSS 1.02475e-19 $X=0.5895 $Y=0.216
c100 16 VSS 5.70081e-19 $X=0.648 $Y=0.0405
c101 10 VSS 7.61325e-20 $X=0.6435 $Y=0.054
c102 5 VSS 0.00241128f $X=0.783 $Y=0.131
c103 2 VSS 0.0591782f $X=0.783 $Y=0.0405
r104 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.131 $X2=0.738 $Y2=0.131
r105 59 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.131 $X2=0.738 $Y2=0.131
r106 57 64 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.693 $Y2=0.131
r107 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.72 $Y2=0.131
r108 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.207 $X2=0.693 $Y2=0.216
r109 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.189 $X2=0.693 $Y2=0.207
r110 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.171 $X2=0.693 $Y2=0.189
r111 52 53 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.165 $X2=0.693 $Y2=0.171
r112 51 52 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.153 $X2=0.693 $Y2=0.165
r113 50 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.225 $X2=0.693 $Y2=0.216
r114 49 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.131
r115 49 51 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.153
r116 47 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.106 $X2=0.693 $Y2=0.114
r117 46 47 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.099 $X2=0.693 $Y2=0.106
r118 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.081 $X2=0.693 $Y2=0.099
r119 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.063 $X2=0.693 $Y2=0.081
r120 43 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.062 $X2=0.693 $Y2=0.063
r121 42 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.131
r122 42 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.114
r123 41 43 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.045 $X2=0.693 $Y2=0.062
r124 39 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.649
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r125 36 39 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.649 $Y2=0.036
r126 36 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r127 34 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.036 $X2=0.693 $Y2=0.045
r128 34 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r129 32 33 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.649 $Y2=0.234
r130 31 32 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.609
+ $Y=0.234 $X2=0.612 $Y2=0.234
r131 30 31 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.595
+ $Y=0.234 $X2=0.609 $Y2=0.234
r132 27 30 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.595 $Y2=0.234
r133 25 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.234 $X2=0.693 $Y2=0.225
r134 25 33 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.234 $X2=0.649 $Y2=0.234
r135 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2295 $X2=0.594 $Y2=0.2295
r136 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r137 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.594 $Y2=0.2295
r138 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.5895 $Y2=0.189
r139 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.189 $X2=0.5895 $Y2=0.189
r140 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r141 13 37 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r142 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.648 $Y2=0.0405
r143 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.6435 $Y2=0.081
r144 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.081 $X2=0.6435 $Y2=0.081
r145 5 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.131 $X2=0.783
+ $Y2=0.131
r146 5 7 369.03 $w=2e-08 $l=9.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.131 $X2=0.783 $Y2=0.2295
r147 2 5 339.058 $w=2e-08 $l=9.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.131
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%12 2 5 7 9 12 14 17 21 25 26 30 31 35 36 37 43 VSS
c33 43 VSS 0.00419842f $X=1.098 $Y=0.234
c34 42 VSS 0.00204425f $X=1.107 $Y=0.234
c35 37 VSS 0.00106107f $X=1.107 $Y=0.171
c36 36 VSS 0.00114275f $X=1.107 $Y=0.117
c37 35 VSS 0.00149546f $X=1.107 $Y=0.225
c38 33 VSS 7.70286e-19 $X=1.073 $Y=0.036
c39 32 VSS 4.41014e-19 $X=1.066 $Y=0.036
c40 31 VSS 0.00146362f $X=1.062 $Y=0.036
c41 30 VSS 0.00481311f $X=1.044 $Y=0.036
c42 26 VSS 0.00226308f $X=1.008 $Y=0.036
c43 25 VSS 0.00460331f $X=1.098 $Y=0.036
c44 21 VSS 7.16657e-19 $X=0.999 $Y=0.105
c45 17 VSS 0.00426839f $X=1.078 $Y=0.2295
c46 12 VSS 0.00485453f $X=1.078 $Y=0.0405
c47 5 VSS 0.00227106f $X=0.999 $Y=0.1055
c48 2 VSS 0.0590816f $X=0.999 $Y=0.0405
r49 43 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r50 42 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r51 39 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.098 $Y2=0.234
r52 36 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.117 $X2=1.107 $Y2=0.171
r53 35 42 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.234
r54 35 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.171
r55 34 36 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.045 $X2=1.107 $Y2=0.117
r56 32 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.066
+ $Y=0.036 $X2=1.073 $Y2=0.036
r57 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=1.062
+ $Y=0.036 $X2=1.066 $Y2=0.036
r58 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=1.062 $Y2=0.036
r59 28 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.036 $X2=1.073 $Y2=0.036
r60 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.008
+ $Y=0.036 $X2=1.044 $Y2=0.036
r61 25 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.098 $Y=0.036 $X2=1.107 $Y2=0.045
r62 25 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.036 $X2=1.08 $Y2=0.036
r63 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.999 $Y=0.045 $X2=1.008 $Y2=0.036
r64 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.045 $X2=0.999 $Y2=0.105
r65 17 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234 $X2=1.08
+ $Y2=0.234
r66 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2295 $X2=1.078 $Y2=0.2295
r67 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.036 $X2=1.08
+ $Y2=0.036
r68 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.0405 $X2=1.078 $Y2=0.0405
r69 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.105 $X2=0.999
+ $Y2=0.105
r70 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.1055 $X2=0.999 $Y2=0.2295
r71 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.0405 $X2=0.999 $Y2=0.1055
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%13 2 7 10 15 18 21 23 25 26 29 30 31 34 35 40 41
+ 43 46 47 48 49 51 54 55 58 68 73 76 78 79 86 VSS
c79 86 VSS 0.0031785f $X=1.269 $Y=0.136
c80 79 VSS 0.00159305f $X=1.229 $Y=0.153
c81 78 VSS 0.00790597f $X=1.175 $Y=0.153
c82 76 VSS 0.00438702f $X=1.269 $Y=0.153
c83 73 VSS 1.90327e-19 $X=0.945 $Y=0.153
c84 68 VSS 0.0033916f $X=0.936 $Y=0.234
c85 67 VSS 0.00253671f $X=0.945 $Y=0.234
c86 58 VSS 4.04001e-19 $X=1.053 $Y=0.14
c87 55 VSS 3.26354e-19 $X=1.008 $Y=0.162
c88 54 VSS 0.00199114f $X=0.99 $Y=0.162
c89 52 VSS 0.00235839f $X=1.044 $Y=0.162
c90 51 VSS 0.00104404f $X=0.945 $Y=0.225
c91 49 VSS 2.07499e-19 $X=0.945 $Y=0.136
c92 48 VSS 2.77769e-19 $X=0.945 $Y=0.119
c93 47 VSS 2.61356e-19 $X=0.945 $Y=0.101
c94 46 VSS 6.393e-19 $X=0.945 $Y=0.081
c95 45 VSS 3.04251e-19 $X=0.945 $Y=0.153
c96 43 VSS 0.00136569f $X=0.92 $Y=0.036
c97 42 VSS 4.8751e-19 $X=0.904 $Y=0.036
c98 41 VSS 0.00146362f $X=0.9 $Y=0.036
c99 40 VSS 0.00358427f $X=0.882 $Y=0.036
c100 35 VSS 0.00347893f $X=0.936 $Y=0.036
c101 34 VSS 0.00276615f $X=0.918 $Y=0.2295
c102 30 VSS 5.63046e-19 $X=0.935 $Y=0.2295
c103 29 VSS 0.0201056f $X=0.864 $Y=0.0405
c104 25 VSS 5.63046e-19 $X=0.881 $Y=0.0405
c105 21 VSS 0.0041584f $X=1.323 $Y=0.136
c106 18 VSS 0.0615048f $X=1.323 $Y=0.0675
c107 10 VSS 0.0581342f $X=1.269 $Y=0.0675
c108 5 VSS 0.00302777f $X=1.053 $Y=0.14
c109 2 VSS 0.0627731f $X=1.053 $Y=0.0405
r110 78 79 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=1.175
+ $Y=0.153 $X2=1.229 $Y2=0.153
r111 76 79 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.269
+ $Y=0.153 $X2=1.229 $Y2=0.153
r112 76 86 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.269 $Y=0.153 $X2=1.269
+ $Y2=0.153
r113 72 78 15.6173 $w=1.8e-08 $l=2.3e-07 $layer=M2 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=1.175 $Y2=0.153
r114 72 73 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.945 $Y=0.153 $X2=0.945
+ $Y2=0.153
r115 68 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r116 67 69 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r117 64 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.234 $X2=0.936 $Y2=0.234
r118 56 58 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.153 $X2=1.053 $Y2=0.14
r119 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.99
+ $Y=0.162 $X2=1.008 $Y2=0.162
r120 53 73 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.945 $Y2=0.162
r121 53 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.99 $Y2=0.162
r122 52 56 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.162 $X2=1.053 $Y2=0.153
r123 52 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.162 $X2=1.008 $Y2=0.162
r124 51 67 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.234
r125 50 73 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.162
r126 50 51 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.225
r127 48 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.119 $X2=0.945 $Y2=0.136
r128 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.101 $X2=0.945 $Y2=0.119
r129 46 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.081 $X2=0.945 $Y2=0.101
r130 45 73 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.162
r131 45 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.136
r132 44 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.081
r133 42 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.904
+ $Y=0.036 $X2=0.92 $Y2=0.036
r134 41 42 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.036 $X2=0.904 $Y2=0.036
r135 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r136 37 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r137 35 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r138 35 43 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.92 $Y2=0.036
r139 34 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.234
+ $X2=0.918 $Y2=0.234
r140 31 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.2295 $X2=0.918 $Y2=0.2295
r141 30 34 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.935 $Y=0.2295 $X2=0.918 $Y2=0.2295
r142 29 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036
+ $X2=0.864 $Y2=0.036
r143 26 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.864 $Y2=0.0405
r144 25 29 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0405 $X2=0.864 $Y2=0.0405
r145 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.136 $X2=1.323 $Y2=0.2025
r146 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.0675 $X2=1.323 $Y2=0.136
r147 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.269
+ $Y=0.136 $X2=1.323 $Y2=0.136
r148 13 86 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.269 $Y=0.136 $X2=1.269
+ $Y2=0.136
r149 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.136 $X2=1.269 $Y2=0.2025
r150 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.0675 $X2=1.269 $Y2=0.136
r151 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.053 $Y=0.14 $X2=1.053
+ $Y2=0.14
r152 5 7 335.312 $w=2e-08 $l=8.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.14 $X2=1.053 $Y2=0.2295
r153 2 5 372.777 $w=2e-08 $l=9.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.0405 $X2=1.053 $Y2=0.14
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%14 1 4 6 11 14 21 23 24 25 VSS
c29 26 VSS 0.00225833f $X=0.485 $Y=0.234
c30 25 VSS 0.00141737f $X=0.461 $Y=0.234
c31 24 VSS 0.0134342f $X=0.447 $Y=0.234
c32 23 VSS 0.00523898f $X=0.309 $Y=0.234
c33 21 VSS 0.00168783f $X=0.486 $Y=0.234
c34 14 VSS 0.0195485f $X=0.542 $Y=0.2025
c35 11 VSS 3.25039e-19 $X=0.557 $Y=0.2025
c36 9 VSS 4.57278e-19 $X=0.484 $Y=0.2025
c37 4 VSS 0.00250858f $X=0.272 $Y=0.2025
c38 1 VSS 3.31752e-19 $X=0.287 $Y=0.2025
r39 25 26 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.461
+ $Y=0.234 $X2=0.485 $Y2=0.234
r40 24 25 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.234 $X2=0.461 $Y2=0.234
r41 23 24 9.37037 $w=1.8e-08 $l=1.38e-07 $layer=M1 $thickness=3.6e-08 $X=0.309
+ $Y=0.234 $X2=0.447 $Y2=0.234
r42 21 26 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.485 $Y2=0.234
r43 17 23 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.309 $Y2=0.234
r44 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.542 $Y2=0.2025
r45 9 14 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.484
+ $Y=0.2025 $X2=0.542 $Y2=0.2025
r46 9 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r47 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.2025 $X2=0.484 $Y2=0.2025
r48 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r49 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.272 $Y2=0.2025
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%16 1 2 5 6 7 10 12 18 20 21 22 23 24 25 VSS
c21 25 VSS 3.8923e-20 $X=0.423 $Y=0.198
c22 24 VSS 8.46035e-21 $X=0.414 $Y=0.198
c23 23 VSS 0.00116854f $X=0.396 $Y=0.198
c24 22 VSS 0.00154511f $X=0.379 $Y=0.198
c25 21 VSS 8.46035e-21 $X=0.36 $Y=0.198
c26 20 VSS 2.61077e-19 $X=0.342 $Y=0.198
c27 18 VSS 3.31089e-19 $X=0.432 $Y=0.198
c28 12 VSS 5.32749e-19 $X=0.324 $Y=0.198
c29 10 VSS 0.00631853f $X=0.432 $Y=0.2025
c30 6 VSS 5.67296e-19 $X=0.449 $Y=0.2025
c31 5 VSS 0.00790786f $X=0.324 $Y=0.2025
c32 1 VSS 6.05629e-19 $X=0.341 $Y=0.2025
r33 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.423 $Y2=0.198
r34 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.414 $Y2=0.198
r35 22 23 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.198 $X2=0.396 $Y2=0.198
r36 21 22 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.198 $X2=0.379 $Y2=0.198
r37 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r38 18 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.423 $Y2=0.198
r39 12 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.342 $Y2=0.198
r40 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r41 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r42 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r43 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198 $X2=0.324
+ $Y2=0.198
r44 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
r45 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%QN 1 2 6 7 10 11 14 16 24 26 VSS
c16 26 VSS 0.00603734f $X=1.377 $Y=0.2
c17 25 VSS 0.0025598f $X=1.377 $Y=0.09
c18 24 VSS 0.00130307f $X=1.377 $Y=0.223
c19 16 VSS 0.0146181f $X=1.368 $Y=0.234
c20 14 VSS 0.00967599f $X=1.296 $Y=0.036
c21 11 VSS 0.0144374f $X=1.368 $Y=0.036
c22 10 VSS 0.010161f $X=1.296 $Y=0.2025
c23 6 VSS 5.72268e-19 $X=1.313 $Y=0.2025
c24 1 VSS 5.72268e-19 $X=1.313 $Y=0.0675
r25 25 26 7.46914 $w=1.8e-08 $l=1.1e-07 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.09 $X2=1.377 $Y2=0.2
r26 24 26 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.223 $X2=1.377 $Y2=0.2
r27 22 24 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.225 $X2=1.377 $Y2=0.223
r28 21 25 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.045 $X2=1.377 $Y2=0.09
r29 16 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.368 $Y=0.234 $X2=1.377 $Y2=0.225
r30 16 18 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.368
+ $Y=0.234 $X2=1.296 $Y2=0.234
r31 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.036 $X2=1.296
+ $Y2=0.036
r32 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.368 $Y=0.036 $X2=1.377 $Y2=0.045
r33 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.368
+ $Y=0.036 $X2=1.296 $Y2=0.036
r34 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.234 $X2=1.296
+ $Y2=0.234
r35 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.279 $Y=0.2025 $X2=1.296 $Y2=0.2025
r36 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.313 $Y=0.2025 $X2=1.296 $Y2=0.2025
r37 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.296
+ $Y=0.0675 $X2=1.296 $Y2=0.036
r38 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.279
+ $Y=0.0675 $X2=1.296 $Y2=0.0675
r39 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.313
+ $Y=0.0675 $X2=1.296 $Y2=0.0675
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%19 1 6 9 VSS
c10 9 VSS 0.0140217f $X=0.704 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.719 $Y=0.2295
c12 4 VSS 2.70811e-19 $X=0.646 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.646
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.631
+ $Y=0.2295 $X2=0.646 $Y2=0.2295
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%20 1 6 9 VSS
c9 9 VSS 0.0145746f $X=0.974 $Y=0.0405
c10 6 VSS 3.14771e-19 $X=0.989 $Y=0.0405
c11 4 VSS 2.65708e-19 $X=0.916 $Y=0.0405
r12 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r13 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.916
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r14 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.901
+ $Y=0.0405 $X2=0.916 $Y2=0.0405
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%22 1 2 VSS
c2 1 VSS 0.00203573f $X=0.719 $Y=0.0405
r3 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0405 $X2=0.685 $Y2=0.0405
.ends

.subckt PM_SDFLX2_ASAP7_75T_SRAM%23 1 2 VSS
c0 1 VSS 0.00214045f $X=0.989 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.2295 $X2=0.955 $Y2=0.2295
.ends


* END of "./SDFLx2_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt SDFLx2_ASAP7_75t_SRAM  VSS VDD CLK SE D SI QN
* 
* QN	QN
* SI	SI
* D	D
* SE	SE
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_9_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_SE_M2_g noxref_15 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 noxref_21 N_6_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 noxref_17 N_D_M4_g noxref_21 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 noxref_15 N_SI_M5_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 N_11_M6_d N_9_M6_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M7 N_22_M7_d N_4_M7_g N_11_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M8 VSS N_10_M8_g N_22_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.027
M9 N_10_M9_d N_11_M9_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_13_M10_d N_4_M10_g N_10_M10_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.827 $Y=0.027
M11 N_20_M11_d N_9_M11_g N_13_M11_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.027
M12 VSS N_12_M12_g N_20_M12_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.027
M13 N_12_M13_d N_13_M13_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.027
M14 VSS N_SE_M14_g N_6_M14_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.027
M15 N_QN_M15_d N_13_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M16 N_QN_M16_d N_13_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.027
M17 VDD N_CLK_M17_g N_4_M17_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M18 N_9_M18_d N_4_M18_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M19 N_16_M19_d N_SE_M19_g N_14_M19_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M20 VDD N_6_M20_g N_16_M20_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M21 N_16_M21_d N_D_M21_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M22 N_14_M22_d N_SI_M22_g N_16_M22_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M23 N_11_M23_d N_4_M23_g N_14_M23_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M24 N_19_M24_d N_9_M24_g N_11_M24_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.611 $Y=0.216
M25 VDD N_10_M25_g N_19_M25_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.216
M26 N_10_M26_d N_11_M26_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M27 N_13_M27_d N_9_M27_g N_10_M27_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.216
M28 N_23_M28_d N_4_M28_g N_13_M28_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.935 $Y=0.216
M29 VDD N_12_M29_g N_23_M29_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.216
M30 N_12_M30_d N_13_M30_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.216
M31 VDD N_SE_M31_g N_6_M31_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.162
M32 N_QN_M32_d N_13_M32_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
M33 N_QN_M33_d N_13_M33_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.162
*
* 
* .include "SDFLx2_ASAP7_75t_SRAM.pex.sp.SDFLX2_ASAP7_75T_SRAM.pxi"
* BEGIN of "./SDFLx2_ASAP7_75t_SRAM.pex.sp.SDFLX2_ASAP7_75T_SRAM.pxi"
* File: SDFLx2_ASAP7_75t_SRAM.pex.sp.SDFLX2_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 13:04:55 2017
* 
x_PM_SDFLX2_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M17_g N_CLK_c_3_p CLK
+ VSS PM_SDFLX2_ASAP7_75T_SRAM%CLK
x_PM_SDFLX2_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_14_n N_4_M18_g N_4_c_25_p N_4_M23_g
+ N_4_M7_g N_4_c_92_p N_4_M10_g N_4_c_76_p N_4_c_24_p N_4_M28_g N_4_M0_s
+ N_4_c_15_n N_4_M17_s N_4_c_16_n N_4_c_17_n N_4_c_18_n N_4_c_41_p N_4_c_19_n
+ N_4_c_59_p N_4_c_26_p N_4_c_27_p N_4_c_37_p N_4_c_28_p N_4_c_20_n N_4_c_21_p
+ N_4_c_29_p N_4_c_56_p VSS PM_SDFLX2_ASAP7_75T_SRAM%4
x_PM_SDFLX2_ASAP7_75T_SRAM%SE N_SE_M2_g N_SE_c_139_p N_SE_M19_g N_SE_M14_g
+ N_SE_c_177_p N_SE_M31_g N_SE_c_145_p N_SE_c_191_p N_SE_c_189_p N_SE_c_207_p
+ N_SE_c_136_n SE N_SE_c_135_n N_SE_c_140_p N_SE_c_141_p N_SE_c_137_n
+ N_SE_c_142_p N_SE_c_143_p N_SE_c_154_p N_SE_c_159_p N_SE_c_148_p N_SE_c_188_p
+ VSS PM_SDFLX2_ASAP7_75T_SRAM%SE
x_PM_SDFLX2_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_218_n N_6_M20_g N_6_M14_s N_6_c_219_n
+ N_6_M31_s N_6_c_222_n N_6_c_257_p N_6_c_267_p N_6_c_254_p N_6_c_263_p
+ N_6_c_271_p N_6_c_249_p N_6_c_215_n N_6_c_216_n N_6_c_224_n N_6_c_225_n
+ N_6_c_228_n N_6_c_229_n N_6_c_256_p VSS PM_SDFLX2_ASAP7_75T_SRAM%6
x_PM_SDFLX2_ASAP7_75T_SRAM%D N_D_M4_g N_D_c_289_n N_D_M21_g D VSS
+ PM_SDFLX2_ASAP7_75T_SRAM%D
x_PM_SDFLX2_ASAP7_75T_SRAM%SI N_SI_M5_g N_SI_M22_g SI N_SI_c_310_n VSS
+ PM_SDFLX2_ASAP7_75T_SRAM%SI
x_PM_SDFLX2_ASAP7_75T_SRAM%9 N_9_M6_g N_9_c_331_n N_9_M24_g N_9_M11_g N_9_c_334_n
+ N_9_M27_g N_9_M1_d N_9_c_400_p N_9_M18_d N_9_c_335_n N_9_c_337_n N_9_c_338_n
+ N_9_c_342_n N_9_c_361_n N_9_c_326_n N_9_c_344_n N_9_c_346_n N_9_c_347_n
+ N_9_c_349_n N_9_c_350_n N_9_c_351_n N_9_c_366_n N_9_c_355_n N_9_c_327_n
+ N_9_c_328_n N_9_c_356_n N_9_c_357_n N_9_c_358_n N_9_c_360_n VSS
+ PM_SDFLX2_ASAP7_75T_SRAM%9
x_PM_SDFLX2_ASAP7_75T_SRAM%10 N_10_M8_g N_10_M25_g N_10_M10_s N_10_M9_d
+ N_10_c_405_n N_10_M26_d N_10_c_406_n N_10_M27_s N_10_c_408_n N_10_c_420_n
+ N_10_c_421_n N_10_c_418_n N_10_c_410_n N_10_c_423_n N_10_c_419_n N_10_c_435_p
+ N_10_c_449_p N_10_c_411_n N_10_c_437_p N_10_c_412_n N_10_c_413_n N_10_c_414_n
+ N_10_c_416_n VSS PM_SDFLX2_ASAP7_75T_SRAM%10
x_PM_SDFLX2_ASAP7_75T_SRAM%11 N_11_M9_g N_11_c_485_n N_11_M26_g N_11_M6_d N_11_M7_s
+ N_11_M23_d N_11_c_453_n N_11_M24_s N_11_c_515_p N_11_c_455_n N_11_c_456_n
+ N_11_c_487_n N_11_c_457_n N_11_c_477_n N_11_c_478_n N_11_c_479_n N_11_c_480_n
+ N_11_c_498_n N_11_c_458_n N_11_c_459_n N_11_c_489_n N_11_c_518_p N_11_c_490_n
+ N_11_c_460_n N_11_c_461_n N_11_c_463_n N_11_c_466_n N_11_c_519_p N_11_c_471_n
+ N_11_c_472_n N_11_c_473_n N_11_c_475_n VSS PM_SDFLX2_ASAP7_75T_SRAM%11
x_PM_SDFLX2_ASAP7_75T_SRAM%12 N_12_M12_g N_12_c_544_p N_12_M29_g N_12_M13_d
+ N_12_c_529_n N_12_M30_d N_12_c_531_n N_12_c_523_n N_12_c_524_n N_12_c_525_n
+ N_12_c_526_n N_12_c_527_n N_12_c_535_n N_12_c_528_n N_12_c_538_n N_12_c_553_p
+ VSS PM_SDFLX2_ASAP7_75T_SRAM%12
x_PM_SDFLX2_ASAP7_75T_SRAM%13 N_13_M13_g N_13_M30_g N_13_M15_g N_13_M32_g
+ N_13_M16_g N_13_c_566_n N_13_M33_g N_13_M11_s N_13_M10_d N_13_c_556_n
+ N_13_M28_s N_13_M27_d N_13_c_558_n N_13_c_568_n N_13_c_569_n N_13_c_570_n
+ N_13_c_571_n N_13_c_572_n N_13_c_559_n N_13_c_590_n N_13_c_560_n N_13_c_561_n
+ N_13_c_633_p N_13_c_610_n N_13_c_612_n N_13_c_562_n N_13_c_563_n N_13_c_573_n
+ N_13_c_574_n N_13_c_575_n N_13_c_577_n VSS PM_SDFLX2_ASAP7_75T_SRAM%13
x_PM_SDFLX2_ASAP7_75T_SRAM%14 N_14_M19_s N_14_c_634_n N_14_M22_d N_14_M23_s
+ N_14_c_635_n N_14_c_645_n N_14_c_637_n N_14_c_642_n N_14_c_638_n VSS
+ PM_SDFLX2_ASAP7_75T_SRAM%14
x_PM_SDFLX2_ASAP7_75T_SRAM%16 N_16_M20_s N_16_M19_d N_16_c_677_n N_16_M22_s
+ N_16_M21_d N_16_c_679_n N_16_c_663_n N_16_c_664_n N_16_c_665_n N_16_c_666_n
+ N_16_c_667_n N_16_c_668_n N_16_c_669_n N_16_c_670_n VSS
+ PM_SDFLX2_ASAP7_75T_SRAM%16
x_PM_SDFLX2_ASAP7_75T_SRAM%QN N_QN_M16_d N_QN_M15_d N_QN_M33_d N_QN_M32_d
+ N_QN_c_685_n N_QN_c_684_n N_QN_c_686_n N_QN_c_687_n QN N_QN_c_698_n VSS
+ PM_SDFLX2_ASAP7_75T_SRAM%QN
x_PM_SDFLX2_ASAP7_75T_SRAM%19 N_19_M24_d N_19_M25_s N_19_c_701_n VSS
+ PM_SDFLX2_ASAP7_75T_SRAM%19
x_PM_SDFLX2_ASAP7_75T_SRAM%20 N_20_M11_d N_20_M12_s N_20_c_710_n VSS
+ PM_SDFLX2_ASAP7_75T_SRAM%20
x_PM_SDFLX2_ASAP7_75T_SRAM%22 N_22_M8_s N_22_M7_d VSS PM_SDFLX2_ASAP7_75T_SRAM%22
x_PM_SDFLX2_ASAP7_75T_SRAM%23 N_23_M29_s N_23_M28_d VSS PM_SDFLX2_ASAP7_75T_SRAM%23
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_CLK_c_2_p N_4_c_14_n 9.79748e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_CLK_c_3_p N_4_c_15_n 2.66516e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.054
cc_4 N_CLK_c_3_p N_4_c_16_n 3.97017e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.081
cc_5 N_CLK_c_3_p N_4_c_17_n 0.00342695f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.164
cc_6 N_CLK_c_3_p N_4_c_18_n 4.97741e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.036
cc_7 N_CLK_c_3_p N_4_c_19_n 0.00171874f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_8 N_CLK_c_3_p N_4_c_20_n 8.1621e-19 $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.189
cc_9 N_CLK_c_3_p N_SE_c_135_n 2.45198e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_10 N_CLK_c_3_p N_9_c_326_n 6.32319e-19 $X=0.081 $Y=0.135 $X2=0.071 $Y2=0.054
cc_11 N_CLK_c_3_p N_9_c_327_n 0.00114506f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_12 N_CLK_c_3_p N_9_c_328_n 4.4946e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_13 N_4_c_21_p N_SE_c_136_n 4.53301e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_14 N_4_c_21_p N_SE_c_137_n 3.907e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_15 N_4_c_21_p N_6_c_215_n 0.0011956f $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_16 N_4_c_24_p N_6_c_216_n 3.37164e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_17 N_4_c_25_p N_SI_M5_g 2.94371e-19 $X=0.567 $Y=0.1355 $X2=0.081 $Y2=0.054
cc_18 N_4_c_26_p SI 0.00114959f $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.135
cc_19 N_4_c_27_p SI 0.00114959f $X=0.567 $Y=0.18 $X2=0.081 $Y2=0.135
cc_20 N_4_c_28_p SI 0.00239259f $X=0.567 $Y=0.189 $X2=0.081 $Y2=0.135
cc_21 N_4_c_29_p SI 0.00167124f $X=0.729 $Y=0.189 $X2=0.081 $Y2=0.135
cc_22 N_4_c_25_p N_SI_c_310_n 5.18435e-19 $X=0.567 $Y=0.1355 $X2=0 $Y2=0
cc_23 N_4_c_25_p N_9_M6_g 0.00365763f $X=0.567 $Y=0.1355 $X2=0.081 $Y2=0.054
cc_24 N_4_M7_g N_9_M6_g 0.00355599f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_25 N_4_c_25_p N_9_c_331_n 9.97803e-19 $X=0.567 $Y=0.1355 $X2=0.081 $Y2=0.135
cc_26 N_4_M10_g N_9_M11_g 0.00355599f $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_27 N_4_c_24_p N_9_M11_g 0.00605856f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.135
cc_28 N_4_c_24_p N_9_c_334_n 0.00180656f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_29 N_4_c_37_p N_9_c_335_n 3.29411e-19 $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_30 N_4_c_20_n N_9_c_335_n 3.38615e-19 $X=0.175 $Y=0.189 $X2=0 $Y2=0
cc_31 N_4_c_21_p N_9_c_337_n 2.67996e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_32 N_4_M1_g N_9_c_338_n 2.57258e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_33 N_4_c_41_p N_9_c_338_n 3.72764e-19 $X=0.054 $Y=0.234 $X2=0 $Y2=0
cc_34 N_4_c_37_p N_9_c_338_n 0.00209054f $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_35 N_4_c_20_n N_9_c_338_n 2.67996e-19 $X=0.175 $Y=0.189 $X2=0 $Y2=0
cc_36 N_4_c_26_p N_9_c_342_n 0.00279251f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_20_n N_9_c_326_n 2.60625e-19 $X=0.175 $Y=0.189 $X2=0 $Y2=0
cc_38 N_4_c_37_p N_9_c_344_n 9.44301e-19 $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_39 N_4_c_21_p N_9_c_344_n 2.46239e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_40 N_4_c_29_p N_9_c_346_n 3.80004e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_41 N_4_c_19_n N_9_c_347_n 3.53344e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_42 N_4_c_21_p N_9_c_347_n 0.0235609f $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_43 N_4_c_29_p N_9_c_349_n 0.0235609f $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_44 N_4_c_24_p N_9_c_350_n 5.51712e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_45 N_4_c_24_p N_9_c_351_n 0.00168667f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_46 N_4_c_26_p N_9_c_351_n 9.87747e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_47 N_4_c_28_p N_9_c_351_n 2.46239e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_48 N_4_c_56_p N_9_c_351_n 2.81643e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_49 N_4_c_24_p N_9_c_355_n 0.00123876f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_50 N_4_c_19_n N_9_c_356_n 9.44301e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_51 N_4_c_59_p N_9_c_357_n 9.44301e-19 $X=0.135 $Y=0.18 $X2=0 $Y2=0
cc_52 N_4_c_37_p N_9_c_358_n 0.00103771f $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_53 N_4_c_21_p N_9_c_358_n 5.9968e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_54 N_4_c_21_p N_9_c_360_n 4.92128e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_55 N_4_M7_g N_10_M8_g 0.00341068f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_56 N_4_M10_g N_10_M8_g 2.13359e-19 $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_57 N_4_c_24_p N_10_M8_g 0.00205997f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_58 N_4_c_56_p N_10_M8_g 3.19768e-19 $X=0.729 $Y=0.18 $X2=0.081 $Y2=0.054
cc_59 N_4_c_24_p N_10_c_405_n 5.52012e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_60 N_4_c_24_p N_10_c_406_n 2.12581e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_61 N_4_c_24_p N_10_M27_s 2.50995e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_62 N_4_M10_g N_10_c_408_n 0.00200065f $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_63 N_4_c_24_p N_10_c_408_n 0.00322783f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_64 N_4_c_24_p N_10_c_410_n 3.41745e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_65 N_4_M10_g N_10_c_411_n 2.74825e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_66 N_4_M10_g N_10_c_412_n 2.10136e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_67 N_4_c_56_p N_10_c_413_n 6.73839e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_68 N_4_c_76_p N_10_c_414_n 0.00195059f $X=0.837 $Y=0.178 $X2=0 $Y2=0
cc_69 N_4_c_24_p N_10_c_414_n 0.00191847f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_70 N_4_M10_g N_10_c_416_n 3.61755e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_71 N_4_M7_g N_11_M9_g 2.13359e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_72 N_4_M10_g N_11_M9_g 0.00341068f $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_73 N_4_c_24_p N_11_M9_g 0.00302156f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_74 N_4_c_26_p N_11_c_453_n 7.70794e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_75 N_4_c_28_p N_11_c_453_n 0.001307f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_76 N_4_c_28_p N_11_c_455_n 0.00138499f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_77 N_4_c_29_p N_11_c_456_n 0.00160025f $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_78 N_4_M7_g N_11_c_457_n 4.38308e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_79 N_4_M7_g N_11_c_458_n 2.0845e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_80 N_4_M7_g N_11_c_459_n 2.27141e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_81 N_4_c_24_p N_11_c_460_n 0.0361494f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_82 N_4_c_24_p N_11_c_461_n 2.38252e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_83 N_4_c_56_p N_11_c_461_n 0.00386452f $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_84 N_4_c_92_p N_11_c_463_n 7.00743e-19 $X=0.675 $Y=0.178 $X2=0 $Y2=0
cc_85 N_4_c_24_p N_11_c_463_n 7.89771e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_86 N_4_c_29_p N_11_c_463_n 4.88732e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_87 N_4_M7_g N_11_c_466_n 2.5554e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_88 N_4_c_24_p N_11_c_466_n 3.47488e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_89 N_4_c_28_p N_11_c_466_n 2.13133e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_90 N_4_c_29_p N_11_c_466_n 4.32971e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_91 N_4_c_56_p N_11_c_466_n 2.60223e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_92 N_4_c_24_p N_11_c_471_n 4.26771e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_93 N_4_c_24_p N_11_c_472_n 4.41163e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_94 N_4_c_24_p N_11_c_473_n 3.33141e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_95 N_4_c_56_p N_11_c_473_n 9.1388e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_96 N_4_M7_g N_11_c_475_n 2.11651e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_97 N_4_c_24_p N_12_M12_g 0.00341068f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_98 N_4_c_24_p N_13_M13_g 2.13359e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_99 N_4_c_24_p N_13_c_556_n 8.27183e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_100 N_4_c_24_p N_13_M28_s 3.37661e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_101 N_4_c_24_p N_13_c_558_n 0.00145657f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_102 N_4_c_24_p N_13_c_559_n 3.13444e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_103 N_4_c_24_p N_13_c_560_n 2.6418e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_104 N_4_c_24_p N_13_c_561_n 0.00294656f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_105 N_4_c_24_p N_13_c_562_n 3.75802e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_106 N_4_c_24_p N_13_c_563_n 5.46321e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_107 N_4_c_21_p N_14_c_634_n 4.92298e-19 $X=0.371 $Y=0.189 $X2=0.081 $Y2=0.135
cc_108 N_4_c_26_p N_14_c_635_n 9.68946e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_109 N_4_c_29_p N_14_c_635_n 6.49405e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_110 N_4_c_21_p N_14_c_637_n 7.84624e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_111 N_4_c_29_p N_14_c_638_n 6.22262e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_112 N_4_c_21_p N_16_c_663_n 2.13751e-19 $X=0.371 $Y=0.189 $X2=0.081 $Y2=0.135
cc_113 N_4_c_29_p N_16_c_664_n 7.1298e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_114 N_4_c_21_p N_16_c_665_n 6.46208e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_115 N_4_c_21_p N_16_c_666_n 4.50553e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_116 N_4_c_21_p N_16_c_667_n 2.85141e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_117 N_4_c_29_p N_16_c_668_n 4.60071e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_118 N_4_c_29_p N_16_c_669_n 4.38038e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_119 N_4_c_29_p N_16_c_670_n 2.31538e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_120 VSS N_4_c_25_p 3.33061e-19 $X=0.567 $Y=0.1355 $X2=0 $Y2=0
cc_121 VSS N_4_c_26_p 0.00110314f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_122 N_4_c_24_p N_19_M25_s 2.33161e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.216
cc_123 N_4_M7_g N_19_c_701_n 0.00248549f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_124 N_4_c_24_p N_19_c_701_n 0.00208457f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_125 N_4_c_29_p N_19_c_701_n 7.88525e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_126 N_4_c_24_p N_20_c_710_n 0.00250239f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_127 N_SE_M2_g N_6_M3_g 0.00304756f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_128 N_SE_c_139_p N_6_c_218_n 0.00126421f $X=0.297 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_129 N_SE_c_140_p N_6_c_219_n 2.80156e-19 $X=1.215 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_130 N_SE_c_141_p N_6_c_219_n 0.00154788f $X=1.215 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_131 N_SE_c_142_p N_6_c_219_n 2.41437e-19 $X=1.175 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_132 N_SE_c_143_p N_6_c_222_n 0.00114532f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_133 N_SE_c_142_p N_6_c_215_n 0.0681088f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_134 N_SE_c_145_p N_6_c_224_n 8.79603e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_135 N_SE_c_141_p N_6_c_225_n 0.00603765f $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_136 N_SE_c_142_p N_6_c_225_n 0.00103045f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_137 N_SE_c_148_p N_6_c_225_n 3.73635e-19 $X=1.215 $Y=0.09 $X2=0 $Y2=0
cc_138 N_SE_c_142_p N_6_c_228_n 2.46239e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_139 N_SE_c_136_n N_6_c_229_n 3.24594e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_140 N_SE_M2_g N_D_M4_g 2.13359e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_141 N_SE_c_135_n N_9_c_361_n 0.00266639f $X=0.225 $Y=0.045 $X2=0 $Y2=0
cc_142 N_SE_c_137_n N_9_c_361_n 4.45368e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_143 N_SE_c_154_p N_9_c_361_n 2.64176e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_144 N_SE_c_136_n N_9_c_349_n 8.13669e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_145 N_SE_c_137_n N_9_c_349_n 0.00228623f $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_146 N_SE_c_142_p N_9_c_366_n 0.00228623f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_147 N_SE_c_154_p N_9_c_327_n 0.00292661f $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_148 N_SE_c_159_p N_9_c_328_n 0.00266639f $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_149 N_SE_c_136_n N_9_c_356_n 0.00266639f $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_150 N_SE_c_142_p N_10_c_405_n 4.38905e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_151 N_SE_c_142_p N_10_c_418_n 3.00479e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_152 N_SE_c_142_p N_10_c_419_n 7.16568e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_153 N_SE_c_142_p N_11_c_457_n 0.00113636f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_154 N_SE_c_142_p N_11_c_477_n 2.78297e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_155 N_SE_c_142_p N_11_c_478_n 5.99401e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_156 N_SE_c_142_p N_11_c_479_n 4.8504e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_157 N_SE_c_142_p N_11_c_480_n 4.65038e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_158 N_SE_c_142_p N_12_c_523_n 5.48108e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_159 N_SE_c_142_p N_12_c_524_n 0.00109158f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_160 N_SE_c_142_p N_12_c_525_n 5.50727e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_161 N_SE_c_142_p N_12_c_526_n 9.11285e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_162 N_SE_c_142_p N_12_c_527_n 4.62125e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_163 N_SE_c_142_p N_12_c_528_n 5.48546e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_164 N_SE_M14_g N_13_M15_g 0.00268443f $X=1.215 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_165 N_SE_M14_g N_13_M16_g 2.13359e-19 $X=1.215 $Y=0.0675 $X2=0 $Y2=0
cc_166 N_SE_c_177_p N_13_c_566_n 0.00112169f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_167 N_SE_c_142_p N_13_c_556_n 2.30689e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_168 N_SE_c_142_p N_13_c_568_n 9.08574e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_169 N_SE_c_142_p N_13_c_569_n 0.00124317f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_170 N_SE_c_142_p N_13_c_570_n 4.54245e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_171 N_SE_c_142_p N_13_c_571_n 4.39544e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_172 N_SE_c_142_p N_13_c_572_n 5.37888e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_173 N_SE_c_141_p N_13_c_573_n 3.26078e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_174 N_SE_c_142_p N_13_c_574_n 9.31342e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_175 N_SE_c_140_p N_13_c_575_n 9.31342e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_176 N_SE_c_143_p N_13_c_575_n 0.00114818f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_177 N_SE_c_188_p N_13_c_577_n 0.00409622f $X=1.215 $Y=0.113 $X2=0 $Y2=0
cc_178 N_SE_c_189_p N_14_c_634_n 2.31793e-19 $X=0.261 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_179 N_SE_M2_g N_14_c_637_n 3.83731e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_180 N_SE_c_191_p N_14_c_637_n 6.51345e-19 $X=0.258 $Y=0.135 $X2=0 $Y2=0
cc_181 VSS N_SE_c_135_n 2.40719e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.135
cc_182 VSS N_SE_c_137_n 5.30841e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.135
cc_183 VSS N_SE_c_154_p 9.86432e-19 $X=0.225 $Y=0.081 $X2=0.081 $Y2=0.135
cc_184 VSS N_SE_c_145_p 0.00129447f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_185 VSS N_SE_c_137_n 7.061e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_186 VSS N_SE_c_154_p 7.68051e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_187 VSS N_SE_c_135_n 8.44602e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.15
cc_188 VSS N_SE_c_137_n 5.36527e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.15
cc_189 VSS N_SE_c_142_p 0.00141783f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_190 VSS N_SE_c_142_p 2.35788e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_191 VSS N_SE_c_137_n 6.93145e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_192 VSS N_SE_c_142_p 9.13621e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_193 VSS N_SE_c_142_p 4.6862e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_194 VSS N_SE_c_142_p 5.41611e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_195 VSS N_SE_c_142_p 8.51044e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_196 VSS N_SE_c_207_p 0.00129447f $X=0.279 $Y=0.135 $X2=0 $Y2=0
cc_197 VSS N_SE_c_137_n 3.48715e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_198 VSS N_SE_c_159_p 9.77595e-19 $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_199 VSS N_SE_c_142_p 2.40178e-19 $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.135
cc_200 VSS N_SE_c_142_p 6.42719e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_201 VSS N_SE_c_142_p 0.00110738f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_202 N_SE_c_141_p N_QN_c_684_n 8.29488e-19 $X=1.215 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_203 N_SE_c_142_p N_20_c_710_n 4.98441e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_204 N_6_M3_g N_D_M4_g 0.00304756f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_205 N_6_c_218_n N_D_c_289_n 9.71463e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_206 N_6_c_215_n D 3.33994e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_207 N_6_c_224_n D 0.00195518f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_208 N_6_c_229_n D 9.77589e-19 $X=0.351 $Y=0.126 $X2=0 $Y2=0
cc_209 N_6_M3_g N_SI_M5_g 2.48122e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_210 N_6_c_215_n SI 3.40688e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_211 N_6_c_215_n N_9_c_342_n 3.98881e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_212 N_6_c_215_n N_9_c_351_n 0.0176151f $X=0.9 $Y=0.081 $X2=0.018 $Y2=0.207
cc_213 N_6_c_224_n N_9_c_351_n 0.00113948f $X=0.351 $Y=0.135 $X2=0.018 $Y2=0.207
cc_214 N_6_c_215_n N_10_c_420_n 5.04077e-19 $X=0.9 $Y=0.081 $X2=0.945 $Y2=0.178
cc_215 N_6_c_215_n N_10_c_421_n 2.53924e-19 $X=0.9 $Y=0.081 $X2=0.945 $Y2=0.178
cc_216 N_6_c_215_n N_10_c_418_n 8.29294e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_217 N_6_c_215_n N_10_c_423_n 5.75824e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_218 N_6_c_215_n N_10_c_416_n 7.91051e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_219 N_6_c_215_n N_11_c_477_n 4.20387e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_220 N_6_c_215_n N_11_c_458_n 4.92006e-19 $X=0.9 $Y=0.081 $X2=0.071 $Y2=0.054
cc_221 N_6_c_215_n N_11_c_459_n 7.19039e-19 $X=0.9 $Y=0.081 $X2=0.056 $Y2=0.054
cc_222 N_6_c_219_n N_12_c_529_n 0.00122694f $X=1.19 $Y=0.0675 $X2=0.567
+ $Y2=0.2025
cc_223 N_6_c_249_p N_12_c_529_n 2.40393e-19 $X=1.161 $Y=0.081 $X2=0.567
+ $Y2=0.2025
cc_224 N_6_c_222_n N_12_c_531_n 4.63408e-19 $X=1.19 $Y=0.2025 $X2=0 $Y2=0
cc_225 N_6_c_249_p N_12_c_523_n 9.95523e-19 $X=1.161 $Y=0.081 $X2=0.837
+ $Y2=0.0405
cc_226 N_6_c_219_n N_12_c_524_n 9.66531e-19 $X=1.19 $Y=0.0675 $X2=0.837
+ $Y2=0.178
cc_227 N_6_c_225_n N_12_c_524_n 0.00241878f $X=1.161 $Y=0.049 $X2=0.837
+ $Y2=0.178
cc_228 N_6_c_254_p N_12_c_535_n 0.00241878f $X=1.17 $Y=0.234 $X2=0 $Y2=0
cc_229 N_6_c_249_p N_12_c_528_n 0.0012739f $X=1.161 $Y=0.081 $X2=0 $Y2=0
cc_230 N_6_c_256_p N_12_c_528_n 0.00241878f $X=1.161 $Y=0.2125 $X2=0 $Y2=0
cc_231 N_6_c_257_p N_12_c_538_n 0.00241878f $X=1.161 $Y=0.225 $X2=0 $Y2=0
cc_232 N_6_c_216_n N_13_c_569_n 6.23859e-19 $X=0.936 $Y=0.081 $X2=0 $Y2=0
cc_233 N_6_c_249_p N_13_c_572_n 3.66836e-19 $X=1.161 $Y=0.081 $X2=0.056
+ $Y2=0.054
cc_234 N_6_c_249_p N_13_c_559_n 5.24665e-19 $X=1.161 $Y=0.081 $X2=0 $Y2=0
cc_235 N_6_c_216_n N_13_c_562_n 3.12147e-19 $X=0.936 $Y=0.081 $X2=0.0505
+ $Y2=0.036
cc_236 N_6_c_219_n N_13_c_574_n 2.31667e-19 $X=1.19 $Y=0.0675 $X2=0.135
+ $Y2=0.135
cc_237 N_6_c_263_p N_13_c_574_n 2.53206e-19 $X=1.179 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_238 N_6_c_249_p N_13_c_574_n 0.00813033f $X=1.161 $Y=0.081 $X2=0.135
+ $Y2=0.135
cc_239 N_6_c_225_n N_13_c_574_n 0.00109426f $X=1.161 $Y=0.049 $X2=0.135
+ $Y2=0.135
cc_240 N_6_c_222_n N_13_c_575_n 3.0124e-19 $X=1.19 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_241 N_6_c_267_p N_13_c_575_n 2.53206e-19 $X=1.188 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_242 N_6_M3_g N_14_c_642_n 2.37298e-19 $X=0.351 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_243 VSS N_6_c_215_n 3.90811e-19 $X=0.9 $Y=0.081 $X2=0.567 $Y2=0.2025
cc_244 VSS N_6_c_228_n 7.35661e-19 $X=0.351 $Y=0.099 $X2=0.567 $Y2=0.2025
cc_245 VSS N_6_c_271_p 6.42252e-19 $X=0.351 $Y=0.081 $X2=0 $Y2=0
cc_246 VSS N_6_c_271_p 0.00369658f $X=0.351 $Y=0.081 $X2=0.837 $Y2=0.0405
cc_247 N_6_M3_g N_16_c_666_n 2.50526e-19 $X=0.351 $Y=0.0675 $X2=0.837 $Y2=0.0405
cc_248 N_6_c_224_n N_16_c_666_n 0.00110314f $X=0.351 $Y=0.135 $X2=0.837
+ $Y2=0.0405
cc_249 VSS N_6_c_228_n 2.30452e-19 $X=0.351 $Y=0.099 $X2=0.135 $Y2=0.135
cc_250 VSS N_6_c_215_n 7.92007e-19 $X=0.9 $Y=0.081 $X2=0.675 $Y2=0.0405
cc_251 VSS N_6_c_271_p 8.14481e-19 $X=0.351 $Y=0.081 $X2=0.675 $Y2=0.178
cc_252 VSS N_6_c_215_n 2.67459e-19 $X=0.9 $Y=0.081 $X2=0.675 $Y2=0.178
cc_253 VSS N_6_c_215_n 3.16736e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_254 VSS N_6_c_215_n 2.43408e-19 $X=0.9 $Y=0.081 $X2=0.837 $Y2=0.0405
cc_255 VSS N_6_c_215_n 5.19239e-19 $X=0.9 $Y=0.081 $X2=0.837 $Y2=0.178
cc_256 N_6_c_222_n N_QN_c_685_n 2.39643e-19 $X=1.19 $Y=0.2025 $X2=0.567
+ $Y2=0.1355
cc_257 N_6_c_219_n N_QN_c_686_n 2.66287e-19 $X=1.19 $Y=0.0675 $X2=0 $Y2=0
cc_258 N_6_c_267_p N_QN_c_687_n 2.72644e-19 $X=1.188 $Y=0.234 $X2=0.675
+ $Y2=0.0405
cc_259 N_6_c_216_n N_20_c_710_n 5.02041e-19 $X=0.936 $Y=0.081 $X2=0.567
+ $Y2=0.1355
cc_260 VSS N_6_c_271_p 2.73492e-19 $X=0.351 $Y=0.081 $X2=0.135 $Y2=0.054
cc_261 N_D_M4_g N_SI_M5_g 0.00348334f $X=0.405 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_262 D SI 7.00288e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_263 N_D_c_289_n N_SI_c_310_n 0.00109838f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_264 D N_9_c_351_n 0.00102191f $X=0.405 $Y=0.134 $X2=0.018 $Y2=0.207
cc_265 N_D_M4_g N_14_c_642_n 2.37298e-19 $X=0.405 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_266 VSS N_D_M4_g 3.08888e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_267 VSS D 5.77345e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_268 N_D_M4_g N_16_c_669_n 2.43567e-19 $X=0.405 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_269 D N_16_c_669_n 0.00108212f $X=0.405 $Y=0.134 $X2=0.837 $Y2=0.178
cc_270 D N_16_c_670_n 3.4434e-19 $X=0.405 $Y=0.134 $X2=0.837 $Y2=0.178
cc_271 VSS D 8.86227e-19 $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.135
cc_272 VSS D 0.00161923f $X=0.405 $Y=0.134 $X2=0.675 $Y2=0.178
cc_273 SI N_9_c_351_n 0.00138386f $X=0.473 $Y=0.135 $X2=0.018 $Y2=0.207
cc_274 SI N_14_c_635_n 0.00560919f $X=0.473 $Y=0.135 $X2=0 $Y2=0
cc_275 SI N_14_c_645_n 0.00167456f $X=0.473 $Y=0.135 $X2=0.837 $Y2=0.0405
cc_276 N_SI_M5_g N_14_c_638_n 2.70361e-19 $X=0.459 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_277 SI N_16_c_664_n 6.69571e-19 $X=0.473 $Y=0.135 $X2=0.675 $Y2=0.178
cc_278 VSS N_SI_M5_g 3.10987e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_279 VSS N_SI_c_310_n 2.08525e-19 $X=0.475 $Y=0.135 $X2=0 $Y2=0
cc_280 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.837 $Y2=0.0405
cc_281 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.837 $Y2=0.0405
cc_282 VSS SI 0.00110314f $X=0.473 $Y=0.135 $X2=0 $Y2=0
cc_283 N_9_M6_g N_10_M8_g 2.82885e-19 $X=0.621 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_284 N_9_c_366_n N_10_c_410_n 5.29207e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_285 N_9_c_355_n N_10_c_411_n 0.00318254f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_286 N_9_c_350_n N_10_c_412_n 0.00128311f $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_287 N_9_M11_g N_11_M9_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_288 N_9_c_334_n N_11_c_485_n 2.98891e-19 $X=0.891 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_289 N_9_c_346_n N_11_c_453_n 3.24488e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_290 N_9_M6_g N_11_c_487_n 3.41974e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_291 N_9_c_346_n N_11_c_487_n 0.00102727f $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_292 N_9_c_342_n N_11_c_489_n 0.00133841f $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_293 N_9_c_351_n N_11_c_490_n 7.726e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_294 N_9_c_346_n N_11_c_460_n 8.63476e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_295 N_9_c_351_n N_11_c_460_n 5.92766e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_296 N_9_c_351_n N_11_c_472_n 3.70527e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_297 N_9_c_366_n N_11_c_473_n 3.70527e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_298 N_9_M11_g N_12_M12_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_299 N_9_M11_g N_13_c_570_n 3.18506e-19 $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_300 N_9_c_355_n N_13_c_570_n 4.09234e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_301 N_9_c_355_n N_13_c_590_n 0.00320381f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_302 N_9_c_355_n N_13_c_563_n 3.56772e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_303 N_9_c_350_n N_13_c_574_n 9.40125e-19 $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_304 N_9_c_335_n N_14_c_634_n 0.0010034f $X=0.16 $Y=0.216 $X2=0.081 $Y2=0.135
cc_305 N_9_c_344_n N_14_c_634_n 0.00105265f $X=0.189 $Y=0.153 $X2=0.081
+ $Y2=0.135
cc_306 N_9_c_351_n N_14_c_635_n 4.24134e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_307 N_9_c_337_n N_14_c_637_n 7.83928e-19 $X=0.18 $Y=0.234 $X2=0 $Y2=0
cc_308 VSS N_9_c_400_p 9.30745e-19 $X=0.16 $Y=0.054 $X2=0.081 $Y2=0.135
cc_309 N_10_M8_g N_11_M9_g 0.00268443f $X=0.729 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_310 N_10_c_418_n N_11_M9_g 3.7702e-19 $X=0.792 $Y=0.09 $X2=0.135 $Y2=0.054
cc_311 N_10_c_419_n N_11_c_480_n 2.46574e-19 $X=0.81 $Y=0.054 $X2=0 $Y2=0
cc_312 N_10_c_420_n N_11_c_498_n 0.00360624f $X=0.747 $Y=0.09 $X2=0 $Y2=0
cc_313 N_10_c_421_n N_11_c_458_n 3.99428e-19 $X=0.747 $Y=0.09 $X2=0.071
+ $Y2=0.054
cc_314 N_10_c_412_n N_11_c_490_n 2.22221e-19 $X=0.837 $Y=0.165 $X2=0.056
+ $Y2=0.216
cc_315 N_10_c_435_p N_11_c_466_n 2.22221e-19 $X=0.837 $Y=0.225 $X2=0.018
+ $Y2=0.045
cc_316 N_10_c_418_n N_11_c_471_n 0.00205899f $X=0.792 $Y=0.09 $X2=0.018
+ $Y2=0.198
cc_317 N_10_c_437_p N_11_c_471_n 7.38434e-19 $X=0.837 $Y=0.14 $X2=0.018
+ $Y2=0.198
cc_318 N_10_M8_g N_11_c_473_n 3.21351e-19 $X=0.729 $Y=0.0405 $X2=0.018 $Y2=0.216
cc_319 N_10_c_420_n N_11_c_473_n 0.00205899f $X=0.747 $Y=0.09 $X2=0.018
+ $Y2=0.216
cc_320 N_10_c_405_n N_13_c_556_n 0.00379158f $X=0.81 $Y=0.0405 $X2=0 $Y2=0
cc_321 N_10_c_419_n N_13_c_556_n 2.84891e-19 $X=0.81 $Y=0.054 $X2=0 $Y2=0
cc_322 N_10_c_416_n N_13_c_556_n 2.08929e-19 $X=0.837 $Y=0.09 $X2=0 $Y2=0
cc_323 N_10_c_408_n N_13_c_558_n 0.00222825f $X=0.866 $Y=0.2295 $X2=0 $Y2=0
cc_324 N_10_c_405_n N_13_c_569_n 3.41768e-19 $X=0.81 $Y=0.0405 $X2=0 $Y2=0
cc_325 N_10_c_416_n N_13_c_559_n 4.2911e-19 $X=0.837 $Y=0.09 $X2=0 $Y2=0
cc_326 N_10_c_414_n N_13_c_561_n 4.2911e-19 $X=0.837 $Y=0.207 $X2=0.056
+ $Y2=0.216
cc_327 N_10_c_408_n N_13_c_562_n 3.64454e-19 $X=0.866 $Y=0.2295 $X2=0.0505
+ $Y2=0.036
cc_328 N_10_c_410_n N_13_c_562_n 4.86017e-19 $X=0.828 $Y=0.234 $X2=0.0505
+ $Y2=0.036
cc_329 N_10_c_449_p N_13_c_563_n 4.2911e-19 $X=0.837 $Y=0.101 $X2=0.054
+ $Y2=0.234
cc_330 N_11_c_453_n N_14_c_635_n 0.00424458f $X=0.594 $Y=0.2025 $X2=0 $Y2=0
cc_331 N_11_c_455_n N_14_c_635_n 4.3429e-19 $X=0.595 $Y=0.234 $X2=0 $Y2=0
cc_332 N_11_c_455_n N_14_c_645_n 2.8677e-19 $X=0.595 $Y=0.234 $X2=0.837
+ $Y2=0.0405
cc_333 VSS N_11_c_453_n 0.0016174f $X=0.594 $Y=0.2025 $X2=0.567 $Y2=0.1355
cc_334 VSS N_11_c_477_n 0.00414127f $X=0.648 $Y=0.036 $X2=0.567 $Y2=0.1355
cc_335 VSS N_11_c_478_n 3.30384e-19 $X=0.649 $Y=0.036 $X2=0.567 $Y2=0.1355
cc_336 VSS N_11_c_477_n 2.79363e-19 $X=0.648 $Y=0.036 $X2=0.675 $Y2=0.0405
cc_337 VSS N_11_c_458_n 2.70508e-19 $X=0.693 $Y=0.081 $X2=0.675 $Y2=0.0405
cc_338 N_11_c_453_n N_19_c_701_n 0.00167238f $X=0.594 $Y=0.2025 $X2=0.567
+ $Y2=0.1355
cc_339 N_11_c_515_p N_19_c_701_n 0.00315491f $X=0.684 $Y=0.234 $X2=0.567
+ $Y2=0.1355
cc_340 N_11_c_487_n N_19_c_701_n 0.00111131f $X=0.649 $Y=0.234 $X2=0.567
+ $Y2=0.1355
cc_341 N_11_c_477_n N_19_c_701_n 5.67227e-19 $X=0.648 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_342 N_11_c_518_p N_19_c_701_n 4.0515e-19 $X=0.693 $Y=0.225 $X2=0.567
+ $Y2=0.1355
cc_343 N_11_c_519_p N_19_c_701_n 0.0409693f $X=0.693 $Y=0.216 $X2=0.567
+ $Y2=0.1355
cc_344 N_11_c_457_n N_22_M8_s 2.44135e-19 $X=0.684 $Y=0.036 $X2=0.135 $Y2=0.054
cc_345 N_11_c_480_n N_22_M8_s 3.62465e-19 $X=0.693 $Y=0.062 $X2=0.135 $Y2=0.054
cc_346 N_12_M12_g N_13_M13_g 0.00268443f $X=0.999 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_347 N_12_c_527_n N_13_M13_g 3.55314e-19 $X=1.062 $Y=0.036 $X2=0.135 $Y2=0.054
cc_348 N_12_c_525_n N_13_c_568_n 0.00136796f $X=1.008 $Y=0.036 $X2=0 $Y2=0
cc_349 N_12_c_523_n N_13_c_572_n 0.00136796f $X=0.999 $Y=0.105 $X2=0.056
+ $Y2=0.054
cc_350 N_12_c_544_p N_13_c_559_n 3.34766e-19 $X=0.999 $Y=0.1055 $X2=0 $Y2=0
cc_351 N_12_c_523_n N_13_c_559_n 0.00136796f $X=0.999 $Y=0.105 $X2=0 $Y2=0
cc_352 N_12_c_535_n N_13_c_561_n 5.28703e-19 $X=1.107 $Y=0.225 $X2=0.056
+ $Y2=0.216
cc_353 N_12_M12_g N_13_c_610_n 6.35734e-19 $X=0.999 $Y=0.0405 $X2=0.018
+ $Y2=0.045
cc_354 N_12_c_523_n N_13_c_610_n 7.99759e-19 $X=0.999 $Y=0.105 $X2=0.018
+ $Y2=0.045
cc_355 N_12_c_527_n N_13_c_612_n 2.75024e-19 $X=1.062 $Y=0.036 $X2=0.018
+ $Y2=0.164
cc_356 N_12_c_538_n N_13_c_612_n 0.00266503f $X=1.107 $Y=0.171 $X2=0.018
+ $Y2=0.164
cc_357 N_12_c_531_n N_13_c_574_n 2.19627e-19 $X=1.078 $Y=0.2295 $X2=0.135
+ $Y2=0.135
cc_358 N_12_c_538_n N_13_c_574_n 0.00106087f $X=1.107 $Y=0.171 $X2=0.135
+ $Y2=0.135
cc_359 N_12_c_553_p N_13_c_574_n 5.80975e-19 $X=1.098 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_360 N_12_c_525_n N_20_c_710_n 5.06067e-19 $X=1.008 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_361 N_13_c_566_n N_QN_M16_d 3.7444e-19 $X=1.323 $Y=0.136 $X2=0.135 $Y2=0.054
cc_362 N_13_c_566_n N_QN_M33_d 3.85232e-19 $X=1.323 $Y=0.136 $X2=0.135 $Y2=0.216
cc_363 N_13_c_566_n N_QN_c_685_n 8.43851e-19 $X=1.323 $Y=0.136 $X2=0.567
+ $Y2=0.1355
cc_364 N_13_c_577_n N_QN_c_685_n 0.00132451f $X=1.269 $Y=0.136 $X2=0.567
+ $Y2=0.1355
cc_365 N_13_M16_g N_QN_c_684_n 4.61823e-19 $X=1.323 $Y=0.0675 $X2=0 $Y2=0
cc_366 N_13_c_566_n N_QN_c_684_n 5.30021e-19 $X=1.323 $Y=0.136 $X2=0 $Y2=0
cc_367 N_13_c_566_n N_QN_c_686_n 7.60428e-19 $X=1.323 $Y=0.136 $X2=0 $Y2=0
cc_368 N_13_c_577_n N_QN_c_686_n 6.27401e-19 $X=1.269 $Y=0.136 $X2=0 $Y2=0
cc_369 N_13_M16_g N_QN_c_687_n 4.56718e-19 $X=1.323 $Y=0.0675 $X2=0.675
+ $Y2=0.0405
cc_370 N_13_c_566_n N_QN_c_687_n 5.38938e-19 $X=1.323 $Y=0.136 $X2=0.675
+ $Y2=0.0405
cc_371 N_13_c_566_n N_QN_c_698_n 3.64455e-19 $X=1.323 $Y=0.136 $X2=0 $Y2=0
cc_372 N_13_c_577_n N_QN_c_698_n 0.00122416f $X=1.269 $Y=0.136 $X2=0 $Y2=0
cc_373 N_13_c_556_n N_20_c_710_n 0.00210698f $X=0.864 $Y=0.0405 $X2=0.567
+ $Y2=0.1355
cc_374 N_13_c_568_n N_20_c_710_n 0.00203632f $X=0.936 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_375 N_13_c_571_n N_20_c_710_n 0.00129774f $X=0.92 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_376 N_13_c_572_n N_20_c_710_n 0.00104094f $X=0.945 $Y=0.081 $X2=0.567
+ $Y2=0.1355
cc_377 N_13_c_633_p N_20_c_710_n 2.5109e-19 $X=0.99 $Y=0.162 $X2=0.567
+ $Y2=0.1355
cc_378 VSS N_14_c_634_n 0.00156967f $X=0.272 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_379 VSS N_14_c_635_n 0.00145872f $X=0.542 $Y=0.2025 $X2=0.675 $Y2=0.178
cc_380 N_14_c_634_n N_16_c_677_n 0.003872f $X=0.272 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_381 N_14_c_642_n N_16_c_677_n 0.00248801f $X=0.447 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_382 N_14_c_635_n N_16_c_679_n 0.00434154f $X=0.542 $Y=0.2025 $X2=0.567
+ $Y2=0.1355
cc_383 N_14_c_642_n N_16_c_679_n 0.0025506f $X=0.447 $Y=0.234 $X2=0.567
+ $Y2=0.1355
cc_384 N_14_c_634_n N_16_c_663_n 3.19827e-19 $X=0.272 $Y=0.2025 $X2=0.567
+ $Y2=0.2025
cc_385 N_14_c_642_n N_16_c_663_n 0.0113176f $X=0.447 $Y=0.234 $X2=0.567
+ $Y2=0.2025
cc_386 VSS N_14_c_635_n 4.53012e-19 $X=0.542 $Y=0.2025 $X2=0.837 $Y2=0.178
cc_387 VSS N_16_c_679_n 0.00141703f $X=0.432 $Y=0.2025 $X2=0.135 $Y2=0.135

* END of "./SDFLx2_ASAP7_75t_SRAM.pex.sp.SDFLX2_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: SDFLx3_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 13:05:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "SDFLx3_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./SDFLx3_ASAP7_75t_SRAM.pex.sp.pex"
* File: SDFLx3_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 13:05:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_SDFLX3_ASAP7_75T_SRAM%CLK 2 5 7 11 16 VSS
c12 11 VSS 0.00713456f $X=0.081 $Y=0.135
c13 5 VSS 0.00188964f $X=0.081 $Y=0.135
c14 2 VSS 0.0628473f $X=0.081 $Y=0.054
r15 11 16 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.15
r16 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%4 2 5 7 10 13 16 19 22 25 28 31 45 48 50 57 58 65
+ 72 79 83 86 90 97 100 101 102 104 123 VSS
c122 134 VSS 7.0154e-20 $X=0.03 $Y=0.189
c123 133 VSS 5.9624e-19 $X=0.027 $Y=0.189
c124 123 VSS 6.49238e-19 $X=0.729 $Y=0.18
c125 104 VSS 0.00976003f $X=0.729 $Y=0.189
c126 102 VSS 0.00542037f $X=0.371 $Y=0.189
c127 101 VSS 0.00609885f $X=0.175 $Y=0.189
c128 100 VSS 0.0013748f $X=0.567 $Y=0.189
c129 97 VSS 0.00291011f $X=0.135 $Y=0.189
c130 93 VSS 5.52785e-19 $X=0.033 $Y=0.189
c131 90 VSS 9.61695e-20 $X=0.567 $Y=0.18
c132 86 VSS 5.76385e-19 $X=0.567 $Y=0.135
c133 83 VSS 1.05495e-19 $X=0.135 $Y=0.18
c134 79 VSS 6.50523e-19 $X=0.135 $Y=0.135
c135 75 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c136 74 VSS 0.00169428f $X=0.047 $Y=0.234
c137 72 VSS 0.0024557f $X=0.054 $Y=0.234
c138 70 VSS 0.00306385f $X=0.027 $Y=0.234
c139 68 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c140 67 VSS 0.00205521f $X=0.047 $Y=0.036
c141 65 VSS 0.00239525f $X=0.054 $Y=0.036
c142 63 VSS 0.00305101f $X=0.027 $Y=0.036
c143 62 VSS 3.84318e-19 $X=0.018 $Y=0.216
c144 61 VSS 3.30259e-19 $X=0.018 $Y=0.207
c145 60 VSS 3.64183e-19 $X=0.018 $Y=0.225
c146 58 VSS 0.0039492f $X=0.018 $Y=0.164
c147 57 VSS 0.00142827f $X=0.018 $Y=0.081
c148 56 VSS 8.21418e-19 $X=0.018 $Y=0.18
c149 53 VSS 0.00514186f $X=0.056 $Y=0.216
c150 50 VSS 2.98509e-19 $X=0.071 $Y=0.216
c151 48 VSS 0.00458629f $X=0.056 $Y=0.054
c152 45 VSS 2.98509e-19 $X=0.071 $Y=0.054
c153 28 VSS 0.108836f $X=0.945 $Y=0.178
c154 25 VSS 1.08457e-19 $X=0.837 $Y=0.178
c155 22 VSS 0.0600244f $X=0.837 $Y=0.0405
c156 19 VSS 2.24613e-19 $X=0.675 $Y=0.178
c157 16 VSS 0.0602569f $X=0.675 $Y=0.0405
c158 10 VSS 0.0660345f $X=0.567 $Y=0.1355
c159 5 VSS 0.00179729f $X=0.135 $Y=0.135
c160 2 VSS 0.0627664f $X=0.135 $Y=0.054
r161 133 134 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.03 $Y2=0.189
r162 130 133 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.027 $Y2=0.189
r163 122 123 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.729 $Y=0.18
+ $X2=0.729 $Y2=0.18
r164 104 123 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.729 $Y=0.189 $X2=0.729
+ $Y2=0.189
r165 101 102 13.3086 $w=1.8e-08 $l=1.96e-07 $layer=M2 $thickness=3.6e-08
+ $X=0.175 $Y=0.189 $X2=0.371 $Y2=0.189
r166 99 104 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.729 $Y2=0.189
r167 99 102 13.3086 $w=1.8e-08 $l=1.96e-07 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.371 $Y2=0.189
r168 99 100 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.567 $Y=0.189 $X2=0.567
+ $Y2=0.189
r169 96 101 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.175 $Y2=0.189
r170 96 97 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.135 $Y=0.189 $X2=0.135
+ $Y2=0.189
r171 93 134 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.03 $Y2=0.189
r172 92 96 6.92593 $w=1.8e-08 $l=1.02e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.135 $Y2=0.189
r173 92 93 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.189 $X2=0.033
+ $Y2=0.189
r174 90 100 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.18 $X2=0.567 $Y2=0.189
r175 89 90 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.171 $X2=0.567 $Y2=0.18
r176 86 89 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.171
r177 83 97 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.18 $X2=0.135 $Y2=0.189
r178 82 83 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.164 $X2=0.135 $Y2=0.18
r179 79 82 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.164
r180 74 75 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r181 72 75 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r182 70 74 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r183 67 68 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r184 65 68 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r185 63 67 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r186 61 62 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.207 $X2=0.018 $Y2=0.216
r187 60 70 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r188 60 62 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.216
r189 59 130 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.189
r190 59 61 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.207
r191 57 58 5.6358 $w=1.8e-08 $l=8.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.164
r192 56 130 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.189
r193 56 58 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.164
r194 55 63 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r195 55 57 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r196 53 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r197 50 53 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r198 48 65 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r199 45 48 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r200 28 31 192.945 $w=2e-08 $l=5.15e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.178 $X2=0.945 $Y2=0.2295
r201 25 28 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08 $X=0.837
+ $Y=0.178 $X2=0.945 $Y2=0.178
r202 25 122 86.044 $w=2.6e-08 $l=1.08e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.837 $Y=0.178 $X2=0.729 $Y2=0.178
r203 22 25 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0405 $X2=0.837 $Y2=0.178
r204 19 122 43.022 $w=2.6e-08 $l=5.4e-08 $layer=LISD $thickness=2.8e-08 $X=0.675
+ $Y=0.178 $X2=0.729 $Y2=0.178
r205 16 19 515.144 $w=2e-08 $l=1.375e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0405 $X2=0.675 $Y2=0.178
r206 10 86 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r207 10 13 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.1355 $X2=0.567 $Y2=0.2025
r208 5 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r209 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r210 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%SE 2 5 7 10 13 15 19 22 23 24 31 33 41 44 45 46 47
+ 54 58 59 62 63 VSS
c80 63 VSS 5.91978e-19 $X=1.215 $Y=0.113
c81 62 VSS 0.00226713f $X=1.215 $Y=0.09
c82 59 VSS 2.63823e-19 $X=0.225 $Y=0.099
c83 58 VSS 5.90201e-19 $X=0.225 $Y=0.081
c84 54 VSS 0.00209148f $X=1.215 $Y=0.136
c85 47 VSS 0.0381258f $X=1.175 $Y=0.045
c86 46 VSS 0.00642311f $X=0.337 $Y=0.045
c87 45 VSS 0.00700109f $X=1.215 $Y=0.045
c88 44 VSS 0.0031469f $X=1.215 $Y=0.045
c89 41 VSS 0.00531f $X=0.225 $Y=0.045
c90 31 VSS 0.00110873f $X=0.225 $Y=0.126
c91 24 VSS 2.51525e-19 $X=0.279 $Y=0.135
c92 23 VSS 1.48251e-19 $X=0.261 $Y=0.135
c93 22 VSS 6.38823e-20 $X=0.258 $Y=0.135
c94 21 VSS 0.00134071f $X=0.255 $Y=0.135
c95 19 VSS 6.89032e-19 $X=0.297 $Y=0.135
c96 13 VSS 0.0019468f $X=1.215 $Y=0.136
c97 10 VSS 0.0611074f $X=1.215 $Y=0.0675
c98 5 VSS 0.0031928f $X=0.297 $Y=0.135
c99 2 VSS 0.063344f $X=0.297 $Y=0.0675
r100 62 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.09 $X2=1.215 $Y2=0.113
r101 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.081 $X2=0.225 $Y2=0.099
r102 54 63 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.136 $X2=1.215 $Y2=0.113
r103 46 47 56.9012 $w=1.8e-08 $l=8.38e-07 $layer=M2 $thickness=3.6e-08 $X=0.337
+ $Y=0.045 $X2=1.175 $Y2=0.045
r104 45 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.215 $Y2=0.09
r105 44 47 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.215
+ $Y=0.045 $X2=1.175 $Y2=0.045
r106 44 45 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.215 $Y=0.045 $X2=1.215
+ $Y2=0.045
r107 41 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.081
r108 40 46 7.60494 $w=1.8e-08 $l=1.12e-07 $layer=M2 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.337 $Y2=0.045
r109 40 41 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.225 $Y=0.045 $X2=0.225
+ $Y2=0.045
r110 31 59 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.099
r111 31 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r112 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.135 $X2=0.279 $Y2=0.135
r113 22 23 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.258
+ $Y=0.135 $X2=0.261 $Y2=0.135
r114 21 22 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.255
+ $Y=0.135 $X2=0.258 $Y2=0.135
r115 19 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.279 $Y2=0.135
r116 17 33 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.225 $Y2=0.135
r117 17 21 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.255 $Y2=0.135
r118 13 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.215 $Y=0.136 $X2=1.215
+ $Y2=0.136
r119 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.136 $X2=1.215 $Y2=0.2025
r120 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.0675 $X2=1.215 $Y2=0.136
r121 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r122 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r123 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%6 2 5 7 9 12 14 17 23 26 28 29 33 36 38 39 43 51
+ 57 58 65 VSS
c72 65 VSS 6.55887e-20 $X=1.161 $Y=0.2125
c73 58 VSS 5.45782e-19 $X=0.351 $Y=0.126
c74 57 VSS 8.0335e-19 $X=0.351 $Y=0.099
c75 51 VSS 0.00278401f $X=1.161 $Y=0.049
c76 43 VSS 3.76741e-19 $X=0.351 $Y=0.135
c77 39 VSS 9.89222e-19 $X=0.936 $Y=0.081
c78 38 VSS 0.00685031f $X=0.9 $Y=0.081
c79 36 VSS 0.00203618f $X=1.161 $Y=0.081
c80 33 VSS 8.1122e-19 $X=0.351 $Y=0.081
c81 29 VSS 6.98259e-19 $X=1.179 $Y=0.234
c82 28 VSS 0.00240687f $X=1.17 $Y=0.234
c83 26 VSS 0.00313492f $X=1.188 $Y=0.234
c84 23 VSS 2.83663e-20 $X=1.161 $Y=0.225
c85 17 VSS 0.00673327f $X=1.19 $Y=0.2025
c86 14 VSS 3.02808e-19 $X=1.205 $Y=0.2025
c87 12 VSS 0.0657106f $X=1.19 $Y=0.0675
c88 9 VSS 3.25039e-19 $X=1.205 $Y=0.0675
c89 5 VSS 0.00125227f $X=0.351 $Y=0.135
c90 2 VSS 0.0585837f $X=0.351 $Y=0.0675
r91 64 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.2 $X2=1.161 $Y2=0.2125
r92 57 58 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.099 $X2=0.351 $Y2=0.126
r93 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.161 $Y=0.049 $X2=1.161
+ $Y2=0.049
r94 43 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.126
r95 38 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.9
+ $Y=0.081 $X2=0.936 $Y2=0.081
r96 37 64 8.08025 $w=1.8e-08 $l=1.19e-07 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.2
r97 37 51 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=1.161 $Y2=0.049
r98 36 39 15.2778 $w=1.8e-08 $l=2.25e-07 $layer=M2 $thickness=3.6e-08 $X=1.161
+ $Y=0.081 $X2=0.936 $Y2=0.081
r99 36 37 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.161 $Y=0.081 $X2=1.161
+ $Y2=0.081
r100 33 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.099
r101 32 38 37.2778 $w=1.8e-08 $l=5.49e-07 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.9 $Y2=0.081
r102 32 33 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.081 $X2=0.351
+ $Y2=0.081
r103 28 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.17
+ $Y=0.234 $X2=1.179 $Y2=0.234
r104 26 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.188
+ $Y=0.234 $X2=1.179 $Y2=0.234
r105 23 65 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.225 $X2=1.161 $Y2=0.2125
r106 22 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.17 $Y2=0.234
r107 22 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.234 $X2=1.161 $Y2=0.225
r108 17 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.188 $Y=0.234
+ $X2=1.188 $Y2=0.234
r109 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.2025 $X2=1.19 $Y2=0.2025
r110 12 50 7.35229 $w=8.1e-08 $l=2.9e-08 $layer=LISD $thickness=2.8e-08 $X=1.19
+ $Y=0.0675 $X2=1.161 $Y2=0.0675
r111 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.0675 $X2=1.19 $Y2=0.0675
r112 5 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r113 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r114 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%D 2 5 7 11 VSS
c18 11 VSS 0.00145113f $X=0.405 $Y=0.134
c19 5 VSS 0.00106786f $X=0.405 $Y=0.135
c20 2 VSS 0.0589243f $X=0.405 $Y=0.0675
r21 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%SI 2 7 11 14 VSS
c21 14 VSS 0.00329293f $X=0.475 $Y=0.135
c22 11 VSS 0.00333153f $X=0.473 $Y=0.135
c23 2 VSS 0.0640988f $X=0.459 $Y=0.0675
r24 11 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.475 $Y=0.135 $X2=0.475
+ $Y2=0.135
r25 5 14 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.475 $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%9 2 5 7 10 13 15 17 20 22 25 27 29 36 43 45 51 55
+ 56 57 59 61 62 69 79 80 81 82 84 85 VSS
c75 86 VSS 5.63033e-20 $X=0.189 $Y=0.216
c76 85 VSS 4.28571e-19 $X=0.189 $Y=0.207
c77 84 VSS 4.04265e-19 $X=0.189 $Y=0.189
c78 82 VSS 2.19344e-19 $X=0.189 $Y=0.1485
c79 81 VSS 3.0092e-19 $X=0.189 $Y=0.144
c80 80 VSS 4.92067e-19 $X=0.189 $Y=0.121
c81 79 VSS 8.32677e-19 $X=0.189 $Y=0.099
c82 69 VSS 0.001222f $X=0.891 $Y=0.135
c83 62 VSS 0.00209834f $X=0.817 $Y=0.153
c84 61 VSS 0.00277455f $X=0.743 $Y=0.153
c85 59 VSS 0.00277965f $X=0.891 $Y=0.153
c86 57 VSS 0.00120333f $X=0.337 $Y=0.153
c87 56 VSS 0.00116325f $X=0.211 $Y=0.153
c88 55 VSS 9.40943e-19 $X=0.621 $Y=0.153
c89 51 VSS 5.62309e-19 $X=0.189 $Y=0.153
c90 48 VSS 5.43917e-20 $X=0.189 $Y=0.225
c91 45 VSS 0.00373046f $X=0.18 $Y=0.036
c92 43 VSS 0.00194932f $X=0.189 $Y=0.036
c93 36 VSS 5.26559e-19 $X=0.621 $Y=0.135
c94 29 VSS 0.00311772f $X=0.162 $Y=0.234
c95 27 VSS 0.00522825f $X=0.18 $Y=0.234
c96 25 VSS 0.00583113f $X=0.16 $Y=0.216
c97 20 VSS 0.00576958f $X=0.16 $Y=0.054
c98 13 VSS 0.00216055f $X=0.891 $Y=0.135
c99 10 VSS 0.0585656f $X=0.891 $Y=0.0405
c100 5 VSS 0.00201785f $X=0.621 $Y=0.135
c101 2 VSS 0.0601628f $X=0.621 $Y=0.0675
r102 85 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.207 $X2=0.189 $Y2=0.216
r103 84 85 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.207
r104 83 84 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.189
r105 81 82 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.1485
r106 80 81 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.121 $X2=0.189 $Y2=0.144
r107 79 80 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.099 $X2=0.189 $Y2=0.121
r108 61 62 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.743
+ $Y=0.153 $X2=0.817 $Y2=0.153
r109 59 62 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.817 $Y2=0.153
r110 59 69 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.153 $X2=0.891
+ $Y2=0.153
r111 56 57 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M2 $thickness=3.6e-08 $X=0.211
+ $Y=0.153 $X2=0.337 $Y2=0.153
r112 54 61 8.28395 $w=1.8e-08 $l=1.22e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.743 $Y2=0.153
r113 54 57 19.284 $w=1.8e-08 $l=2.84e-07 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.337 $Y2=0.153
r114 54 55 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.621 $Y=0.153 $X2=0.621
+ $Y2=0.153
r115 51 83 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.164
r116 51 82 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.1485
r117 50 56 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.211 $Y2=0.153
r118 50 51 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.153 $X2=0.189
+ $Y2=0.153
r119 48 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.216
r120 45 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r121 44 79 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.099
r122 43 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r123 43 44 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r124 40 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r125 36 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.153
r126 27 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.234 $X2=0.189 $Y2=0.225
r127 27 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.162 $Y2=0.234
r128 25 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r129 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r130 20 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r131 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r132 13 69 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.135 $X2=0.891
+ $Y2=0.135
r133 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.135 $X2=0.891 $Y2=0.2295
r134 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.0405 $X2=0.891 $Y2=0.135
r135 5 36 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r136 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2295
r137 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%10 2 7 9 10 13 14 17 19 22 27 28 29 31 36 38 44 45
+ 46 47 48 49 50 54 VSS
c49 56 VSS 5.19568e-19 $X=0.828 $Y=0.09
c50 55 VSS 4.09996e-19 $X=0.819 $Y=0.09
c51 54 VSS 4.29e-19 $X=0.837 $Y=0.09
c52 50 VSS 5.92996e-19 $X=0.837 $Y=0.207
c53 49 VSS 1.19762e-19 $X=0.837 $Y=0.167
c54 48 VSS 1.59501e-19 $X=0.837 $Y=0.165
c55 47 VSS 3.13056e-19 $X=0.837 $Y=0.14
c56 46 VSS 5.61414e-19 $X=0.837 $Y=0.122
c57 45 VSS 1.91116e-19 $X=0.837 $Y=0.101
c58 44 VSS 4.02479e-19 $X=0.837 $Y=0.225
c59 42 VSS 3.58124e-20 $X=0.81 $Y=0.0715
c60 38 VSS 0.00112276f $X=0.81 $Y=0.054
c61 31 VSS 0.00670205f $X=0.828 $Y=0.234
c62 30 VSS 4.74851e-19 $X=0.7965 $Y=0.09
c63 29 VSS 0.00125276f $X=0.792 $Y=0.09
c64 28 VSS 0.00410211f $X=0.747 $Y=0.09
c65 27 VSS 4.49532e-19 $X=0.747 $Y=0.09
c66 24 VSS 1.65079e-19 $X=0.801 $Y=0.09
c67 22 VSS 0.0178177f $X=0.866 $Y=0.2295
c68 19 VSS 3.14771e-19 $X=0.881 $Y=0.2295
c69 17 VSS 2.67274e-19 $X=0.808 $Y=0.2295
c70 13 VSS 0.020153f $X=0.81 $Y=0.0405
c71 9 VSS 6.29543e-19 $X=0.827 $Y=0.0405
c72 2 VSS 0.0580179f $X=0.729 $Y=0.0405
r73 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.819
+ $Y=0.09 $X2=0.828 $Y2=0.09
r74 54 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.09 $X2=0.828 $Y2=0.09
r75 53 55 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.09 $X2=0.819 $Y2=0.09
r76 49 50 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.167 $X2=0.837 $Y2=0.207
r77 48 49 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.165 $X2=0.837 $Y2=0.167
r78 47 48 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.14 $X2=0.837 $Y2=0.165
r79 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.122 $X2=0.837 $Y2=0.14
r80 45 46 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.101 $X2=0.837 $Y2=0.122
r81 44 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.207
r82 43 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.09
r83 43 45 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.099 $X2=0.837 $Y2=0.101
r84 41 42 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.062 $X2=0.81 $Y2=0.0715
r85 38 41 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.054 $X2=0.81 $Y2=0.062
r86 36 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.09
r87 36 42 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.081 $X2=0.81 $Y2=0.0715
r88 31 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r89 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.81 $Y2=0.234
r90 29 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.792
+ $Y=0.09 $X2=0.7965 $Y2=0.09
r91 27 29 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.09 $X2=0.792 $Y2=0.09
r92 27 28 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.747 $Y=0.09 $X2=0.747
+ $Y2=0.09
r93 24 53 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.81 $Y2=0.09
r94 24 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.09 $X2=0.7965 $Y2=0.09
r95 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2295 $X2=0.866 $Y2=0.2295
r96 17 22 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.808
+ $Y=0.2295 $X2=0.866 $Y2=0.2295
r97 17 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.234 $X2=0.81
+ $Y2=0.234
r98 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2295 $X2=0.808 $Y2=0.2295
r99 13 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.054 $X2=0.81
+ $Y2=0.054
r100 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.0405 $X2=0.81 $Y2=0.0405
r101 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.0405 $X2=0.81 $Y2=0.0405
r102 5 28 16.3636 $w=2.2e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.09 $X2=0.747 $Y2=0.09
r103 5 7 522.637 $w=2e-08 $l=1.395e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.09 $X2=0.729 $Y2=0.2295
r104 2 5 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0405 $X2=0.729 $Y2=0.09
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%11 2 5 7 9 14 17 21 22 25 30 31 33 34 37 39 40 43
+ 44 45 46 48 50 51 52 53 54 55 56 59 61 62 64 VSS
c72 64 VSS 1.00092e-19 $X=0.693 $Y=0.131
c73 61 VSS 9.09188e-19 $X=0.72 $Y=0.131
c74 59 VSS 6.42979e-19 $X=0.783 $Y=0.131
c75 56 VSS 1.82087e-19 $X=0.693 $Y=0.216
c76 55 VSS 1.40959e-19 $X=0.693 $Y=0.207
c77 54 VSS 1.07888e-19 $X=0.693 $Y=0.189
c78 53 VSS 1.66071e-19 $X=0.693 $Y=0.171
c79 52 VSS 2.71272e-19 $X=0.693 $Y=0.165
c80 51 VSS 3.53682e-19 $X=0.693 $Y=0.153
c81 50 VSS 2.11704e-19 $X=0.693 $Y=0.225
c82 48 VSS 4.15228e-19 $X=0.693 $Y=0.114
c83 47 VSS 2.7378e-19 $X=0.693 $Y=0.106
c84 46 VSS 5.46003e-20 $X=0.693 $Y=0.099
c85 45 VSS 5.96385e-20 $X=0.693 $Y=0.081
c86 43 VSS 1.65771e-19 $X=0.693 $Y=0.062
c87 42 VSS 2.30403e-19 $X=0.693 $Y=0.122
c88 40 VSS 0.00145015f $X=0.6665 $Y=0.036
c89 39 VSS 0.00201121f $X=0.649 $Y=0.036
c90 37 VSS 0.00303728f $X=0.648 $Y=0.036
c91 34 VSS 0.00412969f $X=0.684 $Y=0.036
c92 33 VSS 0.00297725f $X=0.649 $Y=0.234
c93 32 VSS 2.2805e-19 $X=0.612 $Y=0.234
c94 31 VSS 0.00126734f $X=0.609 $Y=0.234
c95 30 VSS 0.0016591f $X=0.595 $Y=0.234
c96 25 VSS 0.00558865f $X=0.684 $Y=0.234
c97 24 VSS 5.62656e-19 $X=0.594 $Y=0.2295
c98 21 VSS 0.00254121f $X=0.594 $Y=0.2025
c99 18 VSS 1.02475e-19 $X=0.5895 $Y=0.216
c100 16 VSS 5.70081e-19 $X=0.648 $Y=0.0405
c101 10 VSS 7.61325e-20 $X=0.6435 $Y=0.054
c102 5 VSS 0.00241128f $X=0.783 $Y=0.131
c103 2 VSS 0.0591782f $X=0.783 $Y=0.0405
r104 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.131 $X2=0.738 $Y2=0.131
r105 59 62 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.131 $X2=0.738 $Y2=0.131
r106 57 64 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.693 $Y2=0.131
r107 57 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.131 $X2=0.72 $Y2=0.131
r108 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.207 $X2=0.693 $Y2=0.216
r109 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.189 $X2=0.693 $Y2=0.207
r110 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.171 $X2=0.693 $Y2=0.189
r111 52 53 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.165 $X2=0.693 $Y2=0.171
r112 51 52 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.153 $X2=0.693 $Y2=0.165
r113 50 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.225 $X2=0.693 $Y2=0.216
r114 49 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.131
r115 49 51 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.14 $X2=0.693 $Y2=0.153
r116 47 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.106 $X2=0.693 $Y2=0.114
r117 46 47 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.099 $X2=0.693 $Y2=0.106
r118 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.081 $X2=0.693 $Y2=0.099
r119 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.063 $X2=0.693 $Y2=0.081
r120 43 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.062 $X2=0.693 $Y2=0.063
r121 42 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.131
r122 42 48 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.122 $X2=0.693 $Y2=0.114
r123 41 43 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.045 $X2=0.693 $Y2=0.062
r124 39 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.649
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r125 36 39 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.649 $Y2=0.036
r126 36 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r127 34 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.036 $X2=0.693 $Y2=0.045
r128 34 40 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.036 $X2=0.6665 $Y2=0.036
r129 32 33 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.649 $Y2=0.234
r130 31 32 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.609
+ $Y=0.234 $X2=0.612 $Y2=0.234
r131 30 31 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.595
+ $Y=0.234 $X2=0.609 $Y2=0.234
r132 27 30 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.595 $Y2=0.234
r133 25 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.684 $Y=0.234 $X2=0.693 $Y2=0.225
r134 25 33 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.234 $X2=0.649 $Y2=0.234
r135 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2295 $X2=0.594 $Y2=0.2295
r136 21 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r137 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.594 $Y2=0.2295
r138 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.5895 $Y=0.216 $X2=0.5895 $Y2=0.189
r139 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.189 $X2=0.5895 $Y2=0.189
r140 14 16 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0405 $X2=0.648 $Y2=0.0405
r141 13 37 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r142 10 16 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.648 $Y2=0.0405
r143 10 13 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.6435 $Y=0.054 $X2=0.6435 $Y2=0.081
r144 9 13 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.081 $X2=0.6435 $Y2=0.081
r145 5 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.131 $X2=0.783
+ $Y2=0.131
r146 5 7 369.03 $w=2e-08 $l=9.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.131 $X2=0.783 $Y2=0.2295
r147 2 5 339.058 $w=2e-08 $l=9.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0405 $X2=0.783 $Y2=0.131
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%12 2 5 7 9 12 14 17 21 25 26 30 31 35 36 37 43 VSS
c33 43 VSS 0.00419842f $X=1.098 $Y=0.234
c34 42 VSS 0.00204425f $X=1.107 $Y=0.234
c35 37 VSS 0.00106107f $X=1.107 $Y=0.171
c36 36 VSS 0.00114275f $X=1.107 $Y=0.117
c37 35 VSS 0.00149546f $X=1.107 $Y=0.225
c38 33 VSS 7.70286e-19 $X=1.073 $Y=0.036
c39 32 VSS 4.41014e-19 $X=1.066 $Y=0.036
c40 31 VSS 0.00146362f $X=1.062 $Y=0.036
c41 30 VSS 0.00481311f $X=1.044 $Y=0.036
c42 26 VSS 0.00226308f $X=1.008 $Y=0.036
c43 25 VSS 0.00460331f $X=1.098 $Y=0.036
c44 21 VSS 7.16657e-19 $X=0.999 $Y=0.105
c45 17 VSS 0.00426839f $X=1.078 $Y=0.2295
c46 12 VSS 0.00485453f $X=1.078 $Y=0.0405
c47 5 VSS 0.00227106f $X=0.999 $Y=0.1055
c48 2 VSS 0.0590816f $X=0.999 $Y=0.0405
r49 43 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r50 42 44 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.234 $X2=1.1025 $Y2=0.234
r51 39 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.098 $Y2=0.234
r52 36 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.117 $X2=1.107 $Y2=0.171
r53 35 42 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.234
r54 35 37 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.225 $X2=1.107 $Y2=0.171
r55 34 36 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.107
+ $Y=0.045 $X2=1.107 $Y2=0.117
r56 32 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.066
+ $Y=0.036 $X2=1.073 $Y2=0.036
r57 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=1.062
+ $Y=0.036 $X2=1.066 $Y2=0.036
r58 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=1.062 $Y2=0.036
r59 28 33 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.036 $X2=1.073 $Y2=0.036
r60 26 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.008
+ $Y=0.036 $X2=1.044 $Y2=0.036
r61 25 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.098 $Y=0.036 $X2=1.107 $Y2=0.045
r62 25 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.036 $X2=1.08 $Y2=0.036
r63 19 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.999 $Y=0.045 $X2=1.008 $Y2=0.036
r64 19 21 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.045 $X2=0.999 $Y2=0.105
r65 17 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234 $X2=1.08
+ $Y2=0.234
r66 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2295 $X2=1.078 $Y2=0.2295
r67 12 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.036 $X2=1.08
+ $Y2=0.036
r68 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.0405 $X2=1.078 $Y2=0.0405
r69 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.999 $Y=0.105 $X2=0.999
+ $Y2=0.105
r70 5 7 464.566 $w=2e-08 $l=1.24e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.1055 $X2=0.999 $Y2=0.2295
r71 2 5 243.523 $w=2e-08 $l=6.5e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.0405 $X2=0.999 $Y2=0.1055
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%13 2 7 10 15 18 23 26 29 31 33 34 37 38 39 42 43
+ 48 49 51 54 55 56 57 59 62 63 66 76 81 84 86 87 94 VSS
c81 94 VSS 0.0032744f $X=1.269 $Y=0.136
c82 87 VSS 0.00159305f $X=1.229 $Y=0.153
c83 86 VSS 0.00790597f $X=1.175 $Y=0.153
c84 84 VSS 0.00437879f $X=1.269 $Y=0.153
c85 81 VSS 1.90327e-19 $X=0.945 $Y=0.153
c86 76 VSS 0.0033916f $X=0.936 $Y=0.234
c87 75 VSS 0.00253671f $X=0.945 $Y=0.234
c88 66 VSS 4.04001e-19 $X=1.053 $Y=0.14
c89 63 VSS 3.26354e-19 $X=1.008 $Y=0.162
c90 62 VSS 0.00199114f $X=0.99 $Y=0.162
c91 60 VSS 0.00235839f $X=1.044 $Y=0.162
c92 59 VSS 0.00104404f $X=0.945 $Y=0.225
c93 57 VSS 2.07499e-19 $X=0.945 $Y=0.136
c94 56 VSS 2.77769e-19 $X=0.945 $Y=0.119
c95 55 VSS 2.61356e-19 $X=0.945 $Y=0.101
c96 54 VSS 6.393e-19 $X=0.945 $Y=0.081
c97 53 VSS 3.04251e-19 $X=0.945 $Y=0.153
c98 51 VSS 0.00136569f $X=0.92 $Y=0.036
c99 50 VSS 4.8751e-19 $X=0.904 $Y=0.036
c100 49 VSS 0.00146362f $X=0.9 $Y=0.036
c101 48 VSS 0.00358427f $X=0.882 $Y=0.036
c102 43 VSS 0.00347893f $X=0.936 $Y=0.036
c103 42 VSS 0.00276615f $X=0.918 $Y=0.2295
c104 38 VSS 5.63046e-19 $X=0.935 $Y=0.2295
c105 37 VSS 0.0201056f $X=0.864 $Y=0.0405
c106 33 VSS 5.63046e-19 $X=0.881 $Y=0.0405
c107 29 VSS 0.0123941f $X=1.377 $Y=0.136
c108 26 VSS 0.0647964f $X=1.377 $Y=0.0675
c109 18 VSS 0.0615177f $X=1.323 $Y=0.0675
c110 10 VSS 0.0579453f $X=1.269 $Y=0.0675
c111 5 VSS 0.00302777f $X=1.053 $Y=0.14
c112 2 VSS 0.0627731f $X=1.053 $Y=0.0405
r113 86 87 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=1.175
+ $Y=0.153 $X2=1.229 $Y2=0.153
r114 84 87 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.269
+ $Y=0.153 $X2=1.229 $Y2=0.153
r115 84 94 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.269 $Y=0.153 $X2=1.269
+ $Y2=0.153
r116 80 86 15.6173 $w=1.8e-08 $l=2.3e-07 $layer=M2 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=1.175 $Y2=0.153
r117 80 81 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.945 $Y=0.153 $X2=0.945
+ $Y2=0.153
r118 76 77 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r119 75 77 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.234 $X2=0.9405 $Y2=0.234
r120 72 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.234 $X2=0.936 $Y2=0.234
r121 64 66 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.153 $X2=1.053 $Y2=0.14
r122 62 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.99
+ $Y=0.162 $X2=1.008 $Y2=0.162
r123 61 81 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.945 $Y2=0.162
r124 61 62 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.954
+ $Y=0.162 $X2=0.99 $Y2=0.162
r125 60 64 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.162 $X2=1.053 $Y2=0.153
r126 60 63 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.162 $X2=1.008 $Y2=0.162
r127 59 75 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.234
r128 58 81 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.162
r129 58 59 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.171 $X2=0.945 $Y2=0.225
r130 56 57 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.119 $X2=0.945 $Y2=0.136
r131 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.101 $X2=0.945 $Y2=0.119
r132 54 55 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.081 $X2=0.945 $Y2=0.101
r133 53 81 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.162
r134 53 57 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.153 $X2=0.945 $Y2=0.136
r135 52 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.081
r136 50 51 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.904
+ $Y=0.036 $X2=0.92 $Y2=0.036
r137 49 50 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.036 $X2=0.904 $Y2=0.036
r138 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.9 $Y2=0.036
r139 45 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.882 $Y2=0.036
r140 43 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r141 43 51 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.92 $Y2=0.036
r142 42 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.234
+ $X2=0.918 $Y2=0.234
r143 39 42 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.2295 $X2=0.918 $Y2=0.2295
r144 38 42 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.935 $Y=0.2295 $X2=0.918 $Y2=0.2295
r145 37 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036
+ $X2=0.864 $Y2=0.036
r146 34 37 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0405 $X2=0.864 $Y2=0.0405
r147 33 37 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0405 $X2=0.864 $Y2=0.0405
r148 29 31 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.377 $Y=0.136 $X2=1.377 $Y2=0.2025
r149 26 29 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.377 $Y=0.0675 $X2=1.377 $Y2=0.136
r150 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.323
+ $Y=0.136 $X2=1.377 $Y2=0.136
r151 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.136 $X2=1.323 $Y2=0.2025
r152 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.0675 $X2=1.323 $Y2=0.136
r153 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.269
+ $Y=0.136 $X2=1.323 $Y2=0.136
r154 13 94 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.269 $Y=0.136 $X2=1.269
+ $Y2=0.136
r155 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.136 $X2=1.269 $Y2=0.2025
r156 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.0675 $X2=1.269 $Y2=0.136
r157 5 66 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.053 $Y=0.14 $X2=1.053
+ $Y2=0.14
r158 5 7 335.312 $w=2e-08 $l=8.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.14 $X2=1.053 $Y2=0.2295
r159 2 5 372.777 $w=2e-08 $l=9.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.0405 $X2=1.053 $Y2=0.14
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%14 1 4 6 11 14 21 23 24 25 VSS
c29 26 VSS 0.00225833f $X=0.485 $Y=0.234
c30 25 VSS 0.00141737f $X=0.461 $Y=0.234
c31 24 VSS 0.0134342f $X=0.447 $Y=0.234
c32 23 VSS 0.00523898f $X=0.309 $Y=0.234
c33 21 VSS 0.00168783f $X=0.486 $Y=0.234
c34 14 VSS 0.0195485f $X=0.542 $Y=0.2025
c35 11 VSS 3.25039e-19 $X=0.557 $Y=0.2025
c36 9 VSS 4.57278e-19 $X=0.484 $Y=0.2025
c37 4 VSS 0.00250858f $X=0.272 $Y=0.2025
c38 1 VSS 3.31752e-19 $X=0.287 $Y=0.2025
r39 25 26 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.461
+ $Y=0.234 $X2=0.485 $Y2=0.234
r40 24 25 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.234 $X2=0.461 $Y2=0.234
r41 23 24 9.37037 $w=1.8e-08 $l=1.38e-07 $layer=M1 $thickness=3.6e-08 $X=0.309
+ $Y=0.234 $X2=0.447 $Y2=0.234
r42 21 26 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.485 $Y2=0.234
r43 17 23 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.309 $Y2=0.234
r44 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.542 $Y2=0.2025
r45 9 14 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.484
+ $Y=0.2025 $X2=0.542 $Y2=0.2025
r46 9 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r47 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.2025 $X2=0.484 $Y2=0.2025
r48 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r49 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.272 $Y2=0.2025
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%16 1 2 5 6 7 10 12 18 20 21 22 23 24 25 VSS
c21 25 VSS 3.8923e-20 $X=0.423 $Y=0.198
c22 24 VSS 8.46035e-21 $X=0.414 $Y=0.198
c23 23 VSS 0.00116854f $X=0.396 $Y=0.198
c24 22 VSS 0.00154511f $X=0.379 $Y=0.198
c25 21 VSS 8.46035e-21 $X=0.36 $Y=0.198
c26 20 VSS 2.61077e-19 $X=0.342 $Y=0.198
c27 18 VSS 3.31089e-19 $X=0.432 $Y=0.198
c28 12 VSS 5.32749e-19 $X=0.324 $Y=0.198
c29 10 VSS 0.00631853f $X=0.432 $Y=0.2025
c30 6 VSS 5.67296e-19 $X=0.449 $Y=0.2025
c31 5 VSS 0.00790786f $X=0.324 $Y=0.2025
c32 1 VSS 6.05629e-19 $X=0.341 $Y=0.2025
r33 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.198 $X2=0.423 $Y2=0.198
r34 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.414 $Y2=0.198
r35 22 23 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.198 $X2=0.396 $Y2=0.198
r36 21 22 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.198 $X2=0.379 $Y2=0.198
r37 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r38 18 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.423 $Y2=0.198
r39 12 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.342 $Y2=0.198
r40 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r41 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r42 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r43 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198 $X2=0.324
+ $Y2=0.198
r44 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
r45 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.324 $Y2=0.2025
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%QN 1 2 6 11 12 15 16 21 24 29 40 42 VSS
c18 42 VSS 0.00549964f $X=1.431 $Y=0.2
c19 41 VSS 0.00201603f $X=1.431 $Y=0.09
c20 40 VSS 0.00112176f $X=1.428 $Y=0.223
c21 29 VSS 0.019562f $X=1.422 $Y=0.234
c22 28 VSS 0.00635401f $X=1.404 $Y=0.036
c23 24 VSS 0.0096468f $X=1.296 $Y=0.036
c24 21 VSS 0.0193891f $X=1.422 $Y=0.036
c25 19 VSS 0.00662347f $X=1.402 $Y=0.2025
c26 15 VSS 0.010126f $X=1.296 $Y=0.2025
c27 11 VSS 5.72268e-19 $X=1.313 $Y=0.2025
c28 9 VSS 2.69461e-19 $X=1.402 $Y=0.0675
c29 1 VSS 5.72268e-19 $X=1.313 $Y=0.0675
r30 41 42 7.46914 $w=1.8e-08 $l=1.1e-07 $layer=M1 $thickness=3.6e-08 $X=1.431
+ $Y=0.09 $X2=1.431 $Y2=0.2
r31 40 42 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.431
+ $Y=0.223 $X2=1.431 $Y2=0.2
r32 38 40 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.431
+ $Y=0.225 $X2=1.431 $Y2=0.223
r33 37 41 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.431
+ $Y=0.045 $X2=1.431 $Y2=0.09
r34 31 35 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.234 $X2=1.404 $Y2=0.234
r35 29 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.422 $Y=0.234 $X2=1.431 $Y2=0.225
r36 29 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.422
+ $Y=0.234 $X2=1.404 $Y2=0.234
r37 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.404 $Y=0.036 $X2=1.404
+ $Y2=0.036
r38 23 27 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.036 $X2=1.404 $Y2=0.036
r39 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.036 $X2=1.296
+ $Y2=0.036
r40 21 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.422 $Y=0.036 $X2=1.431 $Y2=0.045
r41 21 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.422
+ $Y=0.036 $X2=1.404 $Y2=0.036
r42 19 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.404 $Y=0.234 $X2=1.404
+ $Y2=0.234
r43 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.387 $Y=0.2025 $X2=1.402 $Y2=0.2025
r44 15 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.234 $X2=1.296
+ $Y2=0.234
r45 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.279 $Y=0.2025 $X2=1.296 $Y2=0.2025
r46 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.313 $Y=0.2025 $X2=1.296 $Y2=0.2025
r47 9 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.404
+ $Y=0.0675 $X2=1.404 $Y2=0.036
r48 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.387
+ $Y=0.0675 $X2=1.402 $Y2=0.0675
r49 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.296
+ $Y=0.0675 $X2=1.296 $Y2=0.036
r50 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.279
+ $Y=0.0675 $X2=1.296 $Y2=0.0675
r51 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.313
+ $Y=0.0675 $X2=1.296 $Y2=0.0675
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%19 1 6 9 VSS
c10 9 VSS 0.0140217f $X=0.704 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.719 $Y=0.2295
c12 4 VSS 2.70811e-19 $X=0.646 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.646
+ $Y=0.2295 $X2=0.704 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.631
+ $Y=0.2295 $X2=0.646 $Y2=0.2295
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%20 1 6 9 VSS
c9 9 VSS 0.0145746f $X=0.974 $Y=0.0405
c10 6 VSS 3.14771e-19 $X=0.989 $Y=0.0405
c11 4 VSS 2.65708e-19 $X=0.916 $Y=0.0405
r12 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r13 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.916
+ $Y=0.0405 $X2=0.974 $Y2=0.0405
r14 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.901
+ $Y=0.0405 $X2=0.916 $Y2=0.0405
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%22 1 2 VSS
c2 1 VSS 0.00203573f $X=0.719 $Y=0.0405
r3 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0405 $X2=0.685 $Y2=0.0405
.ends

.subckt PM_SDFLX3_ASAP7_75T_SRAM%23 1 2 VSS
c0 1 VSS 0.00214045f $X=0.989 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.2295 $X2=0.955 $Y2=0.2295
.ends


* END of "./SDFLx3_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt SDFLx3_ASAP7_75t_SRAM  VSS VDD CLK SE D SI QN
* 
* QN	QN
* SI	SI
* D	D
* SE	SE
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_9_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_SE_M2_g noxref_15 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 noxref_21 N_6_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 noxref_17 N_D_M4_g noxref_21 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 noxref_15 N_SI_M5_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 N_11_M6_d N_9_M6_g noxref_17 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M7 N_22_M7_d N_4_M7_g N_11_M7_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M8 VSS N_10_M8_g N_22_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.027
M9 N_10_M9_d N_11_M9_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.027
M10 N_13_M10_d N_4_M10_g N_10_M10_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.827 $Y=0.027
M11 N_20_M11_d N_9_M11_g N_13_M11_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.027
M12 VSS N_12_M12_g N_20_M12_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.027
M13 N_12_M13_d N_13_M13_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.027
M14 VSS N_SE_M14_g N_6_M14_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.027
M15 N_QN_M15_d N_13_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M16 N_QN_M16_d N_13_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.027
M17 N_QN_M17_d N_13_M17_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.367
+ $Y=0.027
M18 VDD N_CLK_M18_g N_4_M18_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M19 N_9_M19_d N_4_M19_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M20 N_16_M20_d N_SE_M20_g N_14_M20_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M21 VDD N_6_M21_g N_16_M21_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M22 N_16_M22_d N_D_M22_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M23 N_14_M23_d N_SI_M23_g N_16_M23_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M24 N_11_M24_d N_4_M24_g N_14_M24_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M25 N_19_M25_d N_9_M25_g N_11_M25_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.611 $Y=0.216
M26 VDD N_10_M26_g N_19_M26_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719
+ $Y=0.216
M27 N_10_M27_d N_11_M27_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.773
+ $Y=0.216
M28 N_13_M28_d N_9_M28_g N_10_M28_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.216
M29 N_23_M29_d N_4_M29_g N_13_M29_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.935 $Y=0.216
M30 VDD N_12_M30_g N_23_M30_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.216
M31 N_12_M31_d N_13_M31_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.216
M32 VDD N_SE_M32_g N_6_M32_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.162
M33 N_QN_M33_d N_13_M33_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
M34 N_QN_M34_d N_13_M34_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.162
M35 N_QN_M35_d N_13_M35_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.367
+ $Y=0.162
*
* 
* .include "SDFLx3_ASAP7_75t_SRAM.pex.sp.SDFLX3_ASAP7_75T_SRAM.pxi"
* BEGIN of "./SDFLx3_ASAP7_75t_SRAM.pex.sp.SDFLX3_ASAP7_75T_SRAM.pxi"
* File: SDFLx3_ASAP7_75t_SRAM.pex.sp.SDFLX3_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 13:05:18 2017
* 
x_PM_SDFLX3_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M18_g N_CLK_c_3_p CLK
+ VSS PM_SDFLX3_ASAP7_75T_SRAM%CLK
x_PM_SDFLX3_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_14_n N_4_M19_g N_4_c_25_p N_4_M24_g
+ N_4_M7_g N_4_c_92_p N_4_M10_g N_4_c_76_p N_4_c_24_p N_4_M29_g N_4_M0_s
+ N_4_c_15_n N_4_M18_s N_4_c_16_n N_4_c_17_n N_4_c_18_n N_4_c_41_p N_4_c_19_n
+ N_4_c_59_p N_4_c_26_p N_4_c_27_p N_4_c_37_p N_4_c_28_p N_4_c_20_n N_4_c_21_p
+ N_4_c_29_p N_4_c_56_p VSS PM_SDFLX3_ASAP7_75T_SRAM%4
x_PM_SDFLX3_ASAP7_75T_SRAM%SE N_SE_M2_g N_SE_c_139_p N_SE_M20_g N_SE_M14_g
+ N_SE_c_177_p N_SE_M32_g N_SE_c_145_p N_SE_c_191_p N_SE_c_189_p N_SE_c_207_p
+ N_SE_c_136_n SE N_SE_c_135_n N_SE_c_140_p N_SE_c_141_p N_SE_c_137_n
+ N_SE_c_142_p N_SE_c_143_p N_SE_c_154_p N_SE_c_159_p N_SE_c_148_p N_SE_c_188_p
+ VSS PM_SDFLX3_ASAP7_75T_SRAM%SE
x_PM_SDFLX3_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_218_n N_6_M21_g N_6_M14_s N_6_c_219_n
+ N_6_M32_s N_6_c_222_n N_6_c_257_p N_6_c_267_p N_6_c_254_p N_6_c_263_p
+ N_6_c_271_p N_6_c_249_p N_6_c_215_n N_6_c_216_n N_6_c_224_n N_6_c_225_n
+ N_6_c_228_n N_6_c_229_n N_6_c_256_p VSS PM_SDFLX3_ASAP7_75T_SRAM%6
x_PM_SDFLX3_ASAP7_75T_SRAM%D N_D_M4_g N_D_c_289_n N_D_M22_g D VSS
+ PM_SDFLX3_ASAP7_75T_SRAM%D
x_PM_SDFLX3_ASAP7_75T_SRAM%SI N_SI_M5_g N_SI_M23_g SI N_SI_c_310_n VSS
+ PM_SDFLX3_ASAP7_75T_SRAM%SI
x_PM_SDFLX3_ASAP7_75T_SRAM%9 N_9_M6_g N_9_c_331_n N_9_M25_g N_9_M11_g N_9_c_334_n
+ N_9_M28_g N_9_M1_d N_9_c_400_p N_9_M19_d N_9_c_335_n N_9_c_337_n N_9_c_338_n
+ N_9_c_342_n N_9_c_361_n N_9_c_326_n N_9_c_344_n N_9_c_346_n N_9_c_347_n
+ N_9_c_349_n N_9_c_350_n N_9_c_351_n N_9_c_366_n N_9_c_355_n N_9_c_327_n
+ N_9_c_328_n N_9_c_356_n N_9_c_357_n N_9_c_358_n N_9_c_360_n VSS
+ PM_SDFLX3_ASAP7_75T_SRAM%9
x_PM_SDFLX3_ASAP7_75T_SRAM%10 N_10_M8_g N_10_M26_g N_10_M10_s N_10_M9_d
+ N_10_c_405_n N_10_M27_d N_10_c_406_n N_10_M28_s N_10_c_408_n N_10_c_420_n
+ N_10_c_421_n N_10_c_418_n N_10_c_410_n N_10_c_423_n N_10_c_419_n N_10_c_435_p
+ N_10_c_449_p N_10_c_411_n N_10_c_437_p N_10_c_412_n N_10_c_413_n N_10_c_414_n
+ N_10_c_416_n VSS PM_SDFLX3_ASAP7_75T_SRAM%10
x_PM_SDFLX3_ASAP7_75T_SRAM%11 N_11_M9_g N_11_c_485_n N_11_M27_g N_11_M6_d N_11_M7_s
+ N_11_M24_d N_11_c_453_n N_11_M25_s N_11_c_515_p N_11_c_455_n N_11_c_456_n
+ N_11_c_487_n N_11_c_457_n N_11_c_477_n N_11_c_478_n N_11_c_479_n N_11_c_480_n
+ N_11_c_498_n N_11_c_458_n N_11_c_459_n N_11_c_489_n N_11_c_518_p N_11_c_490_n
+ N_11_c_460_n N_11_c_461_n N_11_c_463_n N_11_c_466_n N_11_c_519_p N_11_c_471_n
+ N_11_c_472_n N_11_c_473_n N_11_c_475_n VSS PM_SDFLX3_ASAP7_75T_SRAM%11
x_PM_SDFLX3_ASAP7_75T_SRAM%12 N_12_M12_g N_12_c_544_p N_12_M30_g N_12_M13_d
+ N_12_c_529_n N_12_M31_d N_12_c_531_n N_12_c_523_n N_12_c_524_n N_12_c_525_n
+ N_12_c_526_n N_12_c_527_n N_12_c_535_n N_12_c_528_n N_12_c_538_n N_12_c_553_p
+ VSS PM_SDFLX3_ASAP7_75T_SRAM%12
x_PM_SDFLX3_ASAP7_75T_SRAM%13 N_13_M13_g N_13_M31_g N_13_M15_g N_13_M33_g
+ N_13_M16_g N_13_M34_g N_13_M17_g N_13_c_566_n N_13_M35_g N_13_M11_s N_13_M10_d
+ N_13_c_556_n N_13_M29_s N_13_M28_d N_13_c_558_n N_13_c_568_n N_13_c_569_n
+ N_13_c_570_n N_13_c_571_n N_13_c_572_n N_13_c_559_n N_13_c_590_n N_13_c_560_n
+ N_13_c_561_n N_13_c_635_p N_13_c_610_n N_13_c_612_n N_13_c_562_n N_13_c_563_n
+ N_13_c_573_n N_13_c_574_n N_13_c_575_n N_13_c_577_n VSS
+ PM_SDFLX3_ASAP7_75T_SRAM%13
x_PM_SDFLX3_ASAP7_75T_SRAM%14 N_14_M20_s N_14_c_636_n N_14_M23_d N_14_M24_s
+ N_14_c_637_n N_14_c_647_n N_14_c_639_n N_14_c_644_n N_14_c_640_n VSS
+ PM_SDFLX3_ASAP7_75T_SRAM%14
x_PM_SDFLX3_ASAP7_75T_SRAM%16 N_16_M21_s N_16_M20_d N_16_c_679_n N_16_M23_s
+ N_16_M22_d N_16_c_681_n N_16_c_665_n N_16_c_666_n N_16_c_667_n N_16_c_668_n
+ N_16_c_669_n N_16_c_670_n N_16_c_671_n N_16_c_672_n VSS
+ PM_SDFLX3_ASAP7_75T_SRAM%16
x_PM_SDFLX3_ASAP7_75T_SRAM%QN N_QN_M16_d N_QN_M15_d N_QN_M17_d N_QN_M34_d
+ N_QN_M33_d N_QN_c_687_n N_QN_M35_d N_QN_c_686_n N_QN_c_688_n N_QN_c_689_n QN
+ N_QN_c_702_n VSS PM_SDFLX3_ASAP7_75T_SRAM%QN
x_PM_SDFLX3_ASAP7_75T_SRAM%19 N_19_M25_d N_19_M26_s N_19_c_705_n VSS
+ PM_SDFLX3_ASAP7_75T_SRAM%19
x_PM_SDFLX3_ASAP7_75T_SRAM%20 N_20_M11_d N_20_M12_s N_20_c_714_n VSS
+ PM_SDFLX3_ASAP7_75T_SRAM%20
x_PM_SDFLX3_ASAP7_75T_SRAM%22 N_22_M8_s N_22_M7_d VSS PM_SDFLX3_ASAP7_75T_SRAM%22
x_PM_SDFLX3_ASAP7_75T_SRAM%23 N_23_M30_s N_23_M29_d VSS PM_SDFLX3_ASAP7_75T_SRAM%23
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_CLK_c_2_p N_4_c_14_n 9.79748e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_CLK_c_3_p N_4_c_15_n 2.66516e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.054
cc_4 N_CLK_c_3_p N_4_c_16_n 3.97017e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.081
cc_5 N_CLK_c_3_p N_4_c_17_n 0.00342695f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.164
cc_6 N_CLK_c_3_p N_4_c_18_n 4.97741e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.036
cc_7 N_CLK_c_3_p N_4_c_19_n 0.00171874f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_8 N_CLK_c_3_p N_4_c_20_n 8.1621e-19 $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.189
cc_9 N_CLK_c_3_p N_SE_c_135_n 2.45198e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_10 N_CLK_c_3_p N_9_c_326_n 6.32319e-19 $X=0.081 $Y=0.135 $X2=0.071 $Y2=0.054
cc_11 N_CLK_c_3_p N_9_c_327_n 0.00114506f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_12 N_CLK_c_3_p N_9_c_328_n 4.4946e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_13 N_4_c_21_p N_SE_c_136_n 4.53301e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_14 N_4_c_21_p N_SE_c_137_n 3.907e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_15 N_4_c_21_p N_6_c_215_n 0.0011956f $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_16 N_4_c_24_p N_6_c_216_n 3.37164e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_17 N_4_c_25_p N_SI_M5_g 2.94371e-19 $X=0.567 $Y=0.1355 $X2=0.081 $Y2=0.054
cc_18 N_4_c_26_p SI 0.00114959f $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.135
cc_19 N_4_c_27_p SI 0.00114959f $X=0.567 $Y=0.18 $X2=0.081 $Y2=0.135
cc_20 N_4_c_28_p SI 0.00239259f $X=0.567 $Y=0.189 $X2=0.081 $Y2=0.135
cc_21 N_4_c_29_p SI 0.00167124f $X=0.729 $Y=0.189 $X2=0.081 $Y2=0.135
cc_22 N_4_c_25_p N_SI_c_310_n 5.18435e-19 $X=0.567 $Y=0.1355 $X2=0 $Y2=0
cc_23 N_4_c_25_p N_9_M6_g 0.00365763f $X=0.567 $Y=0.1355 $X2=0.081 $Y2=0.054
cc_24 N_4_M7_g N_9_M6_g 0.00355599f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_25 N_4_c_25_p N_9_c_331_n 9.97803e-19 $X=0.567 $Y=0.1355 $X2=0.081 $Y2=0.135
cc_26 N_4_M10_g N_9_M11_g 0.00355599f $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_27 N_4_c_24_p N_9_M11_g 0.00605856f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.135
cc_28 N_4_c_24_p N_9_c_334_n 0.00180656f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_29 N_4_c_37_p N_9_c_335_n 3.29411e-19 $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_30 N_4_c_20_n N_9_c_335_n 3.38615e-19 $X=0.175 $Y=0.189 $X2=0 $Y2=0
cc_31 N_4_c_21_p N_9_c_337_n 2.67996e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_32 N_4_M1_g N_9_c_338_n 2.57258e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_33 N_4_c_41_p N_9_c_338_n 3.72764e-19 $X=0.054 $Y=0.234 $X2=0 $Y2=0
cc_34 N_4_c_37_p N_9_c_338_n 0.00209054f $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_35 N_4_c_20_n N_9_c_338_n 2.67996e-19 $X=0.175 $Y=0.189 $X2=0 $Y2=0
cc_36 N_4_c_26_p N_9_c_342_n 0.00279251f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_20_n N_9_c_326_n 2.60625e-19 $X=0.175 $Y=0.189 $X2=0 $Y2=0
cc_38 N_4_c_37_p N_9_c_344_n 9.44301e-19 $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_39 N_4_c_21_p N_9_c_344_n 2.46239e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_40 N_4_c_29_p N_9_c_346_n 3.80004e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_41 N_4_c_19_n N_9_c_347_n 3.53344e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_42 N_4_c_21_p N_9_c_347_n 0.0235609f $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_43 N_4_c_29_p N_9_c_349_n 0.0235609f $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_44 N_4_c_24_p N_9_c_350_n 5.51712e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_45 N_4_c_24_p N_9_c_351_n 0.00168667f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_46 N_4_c_26_p N_9_c_351_n 9.87747e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_47 N_4_c_28_p N_9_c_351_n 2.46239e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_48 N_4_c_56_p N_9_c_351_n 2.81643e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_49 N_4_c_24_p N_9_c_355_n 0.00123876f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_50 N_4_c_19_n N_9_c_356_n 9.44301e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_51 N_4_c_59_p N_9_c_357_n 9.44301e-19 $X=0.135 $Y=0.18 $X2=0 $Y2=0
cc_52 N_4_c_37_p N_9_c_358_n 0.00103771f $X=0.135 $Y=0.189 $X2=0 $Y2=0
cc_53 N_4_c_21_p N_9_c_358_n 5.9968e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_54 N_4_c_21_p N_9_c_360_n 4.92128e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_55 N_4_M7_g N_10_M8_g 0.00341068f $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_56 N_4_M10_g N_10_M8_g 2.13359e-19 $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_57 N_4_c_24_p N_10_M8_g 0.00205997f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_58 N_4_c_56_p N_10_M8_g 3.19768e-19 $X=0.729 $Y=0.18 $X2=0.081 $Y2=0.054
cc_59 N_4_c_24_p N_10_c_405_n 5.52012e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_60 N_4_c_24_p N_10_c_406_n 2.12581e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_61 N_4_c_24_p N_10_M28_s 2.50995e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_62 N_4_M10_g N_10_c_408_n 0.00200065f $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_63 N_4_c_24_p N_10_c_408_n 0.00322783f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_64 N_4_c_24_p N_10_c_410_n 3.41745e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_65 N_4_M10_g N_10_c_411_n 2.74825e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_66 N_4_M10_g N_10_c_412_n 2.10136e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_67 N_4_c_56_p N_10_c_413_n 6.73839e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_68 N_4_c_76_p N_10_c_414_n 0.00195059f $X=0.837 $Y=0.178 $X2=0 $Y2=0
cc_69 N_4_c_24_p N_10_c_414_n 0.00191847f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_70 N_4_M10_g N_10_c_416_n 3.61755e-19 $X=0.837 $Y=0.0405 $X2=0 $Y2=0
cc_71 N_4_M7_g N_11_M9_g 2.13359e-19 $X=0.675 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_72 N_4_M10_g N_11_M9_g 0.00341068f $X=0.837 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_73 N_4_c_24_p N_11_M9_g 0.00302156f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_74 N_4_c_26_p N_11_c_453_n 7.70794e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_75 N_4_c_28_p N_11_c_453_n 0.001307f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_76 N_4_c_28_p N_11_c_455_n 0.00138499f $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_77 N_4_c_29_p N_11_c_456_n 0.00160025f $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_78 N_4_M7_g N_11_c_457_n 4.38308e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_79 N_4_M7_g N_11_c_458_n 2.0845e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_80 N_4_M7_g N_11_c_459_n 2.27141e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_81 N_4_c_24_p N_11_c_460_n 0.0361494f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_82 N_4_c_24_p N_11_c_461_n 2.38252e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_83 N_4_c_56_p N_11_c_461_n 0.00386452f $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_84 N_4_c_92_p N_11_c_463_n 7.00743e-19 $X=0.675 $Y=0.178 $X2=0 $Y2=0
cc_85 N_4_c_24_p N_11_c_463_n 7.89771e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_86 N_4_c_29_p N_11_c_463_n 4.88732e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_87 N_4_M7_g N_11_c_466_n 2.5554e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_88 N_4_c_24_p N_11_c_466_n 3.47488e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_89 N_4_c_28_p N_11_c_466_n 2.13133e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_90 N_4_c_29_p N_11_c_466_n 4.32971e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_91 N_4_c_56_p N_11_c_466_n 2.60223e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_92 N_4_c_24_p N_11_c_471_n 4.26771e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_93 N_4_c_24_p N_11_c_472_n 4.41163e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_94 N_4_c_24_p N_11_c_473_n 3.33141e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_95 N_4_c_56_p N_11_c_473_n 9.1388e-19 $X=0.729 $Y=0.18 $X2=0 $Y2=0
cc_96 N_4_M7_g N_11_c_475_n 2.11651e-19 $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_97 N_4_c_24_p N_12_M12_g 0.00341068f $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_98 N_4_c_24_p N_13_M13_g 2.13359e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.054
cc_99 N_4_c_24_p N_13_c_556_n 8.27183e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_100 N_4_c_24_p N_13_M29_s 3.37661e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_101 N_4_c_24_p N_13_c_558_n 0.00145657f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_102 N_4_c_24_p N_13_c_559_n 3.13444e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_103 N_4_c_24_p N_13_c_560_n 2.6418e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_104 N_4_c_24_p N_13_c_561_n 0.00294656f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_105 N_4_c_24_p N_13_c_562_n 3.75802e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_106 N_4_c_24_p N_13_c_563_n 5.46321e-19 $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_107 N_4_c_21_p N_14_c_636_n 4.92298e-19 $X=0.371 $Y=0.189 $X2=0.081 $Y2=0.135
cc_108 N_4_c_26_p N_14_c_637_n 9.68946e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_109 N_4_c_29_p N_14_c_637_n 6.49405e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_110 N_4_c_21_p N_14_c_639_n 7.84624e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_111 N_4_c_29_p N_14_c_640_n 6.22262e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_112 N_4_c_21_p N_16_c_665_n 2.13751e-19 $X=0.371 $Y=0.189 $X2=0.081 $Y2=0.135
cc_113 N_4_c_29_p N_16_c_666_n 7.1298e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_114 N_4_c_21_p N_16_c_667_n 6.46208e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_115 N_4_c_21_p N_16_c_668_n 4.50553e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_116 N_4_c_21_p N_16_c_669_n 2.85141e-19 $X=0.371 $Y=0.189 $X2=0 $Y2=0
cc_117 N_4_c_29_p N_16_c_670_n 4.60071e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_118 N_4_c_29_p N_16_c_671_n 4.38038e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_119 N_4_c_29_p N_16_c_672_n 2.31538e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_120 VSS N_4_c_25_p 3.33061e-19 $X=0.567 $Y=0.1355 $X2=0 $Y2=0
cc_121 VSS N_4_c_26_p 0.00110314f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_122 N_4_c_24_p N_19_M26_s 2.33161e-19 $X=0.945 $Y=0.178 $X2=0.081 $Y2=0.216
cc_123 N_4_M7_g N_19_c_705_n 0.00248549f $X=0.675 $Y=0.0405 $X2=0 $Y2=0
cc_124 N_4_c_24_p N_19_c_705_n 0.00208457f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_125 N_4_c_29_p N_19_c_705_n 7.88525e-19 $X=0.729 $Y=0.189 $X2=0 $Y2=0
cc_126 N_4_c_24_p N_20_c_714_n 0.00250239f $X=0.945 $Y=0.178 $X2=0 $Y2=0
cc_127 N_SE_M2_g N_6_M3_g 0.00304756f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_128 N_SE_c_139_p N_6_c_218_n 0.00126421f $X=0.297 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_129 N_SE_c_140_p N_6_c_219_n 2.80156e-19 $X=1.215 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_130 N_SE_c_141_p N_6_c_219_n 0.00154788f $X=1.215 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_131 N_SE_c_142_p N_6_c_219_n 2.41437e-19 $X=1.175 $Y=0.045 $X2=0.081
+ $Y2=0.135
cc_132 N_SE_c_143_p N_6_c_222_n 0.00114532f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_133 N_SE_c_142_p N_6_c_215_n 0.0681088f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_134 N_SE_c_145_p N_6_c_224_n 8.79603e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_135 N_SE_c_141_p N_6_c_225_n 0.00603765f $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_136 N_SE_c_142_p N_6_c_225_n 0.00103045f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_137 N_SE_c_148_p N_6_c_225_n 3.73635e-19 $X=1.215 $Y=0.09 $X2=0 $Y2=0
cc_138 N_SE_c_142_p N_6_c_228_n 2.46239e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_139 N_SE_c_136_n N_6_c_229_n 3.24594e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_140 N_SE_M2_g N_D_M4_g 2.13359e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_141 N_SE_c_135_n N_9_c_361_n 0.00266639f $X=0.225 $Y=0.045 $X2=0 $Y2=0
cc_142 N_SE_c_137_n N_9_c_361_n 4.45368e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_143 N_SE_c_154_p N_9_c_361_n 2.64176e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_144 N_SE_c_136_n N_9_c_349_n 8.13669e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_145 N_SE_c_137_n N_9_c_349_n 0.00228623f $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_146 N_SE_c_142_p N_9_c_366_n 0.00228623f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_147 N_SE_c_154_p N_9_c_327_n 0.00292661f $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_148 N_SE_c_159_p N_9_c_328_n 0.00266639f $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_149 N_SE_c_136_n N_9_c_356_n 0.00266639f $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_150 N_SE_c_142_p N_10_c_405_n 4.38905e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_151 N_SE_c_142_p N_10_c_418_n 3.00479e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_152 N_SE_c_142_p N_10_c_419_n 7.16568e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_153 N_SE_c_142_p N_11_c_457_n 0.00113636f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_154 N_SE_c_142_p N_11_c_477_n 2.78297e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_155 N_SE_c_142_p N_11_c_478_n 5.99401e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_156 N_SE_c_142_p N_11_c_479_n 4.8504e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_157 N_SE_c_142_p N_11_c_480_n 4.65038e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_158 N_SE_c_142_p N_12_c_523_n 5.48108e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_159 N_SE_c_142_p N_12_c_524_n 0.00109158f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_160 N_SE_c_142_p N_12_c_525_n 5.50727e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_161 N_SE_c_142_p N_12_c_526_n 9.11285e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_162 N_SE_c_142_p N_12_c_527_n 4.62125e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_163 N_SE_c_142_p N_12_c_528_n 5.48546e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_164 N_SE_M14_g N_13_M15_g 0.00268443f $X=1.215 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_165 N_SE_M14_g N_13_M16_g 2.13359e-19 $X=1.215 $Y=0.0675 $X2=0 $Y2=0
cc_166 N_SE_c_177_p N_13_c_566_n 0.00112628f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_167 N_SE_c_142_p N_13_c_556_n 2.30689e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_168 N_SE_c_142_p N_13_c_568_n 9.08574e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_169 N_SE_c_142_p N_13_c_569_n 0.00124317f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_170 N_SE_c_142_p N_13_c_570_n 4.54245e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_171 N_SE_c_142_p N_13_c_571_n 4.39544e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_172 N_SE_c_142_p N_13_c_572_n 5.37888e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_173 N_SE_c_141_p N_13_c_573_n 3.26078e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_174 N_SE_c_142_p N_13_c_574_n 9.31342e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_175 N_SE_c_140_p N_13_c_575_n 9.31342e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_176 N_SE_c_143_p N_13_c_575_n 0.00114818f $X=1.215 $Y=0.136 $X2=0 $Y2=0
cc_177 N_SE_c_188_p N_13_c_577_n 0.00409622f $X=1.215 $Y=0.113 $X2=0 $Y2=0
cc_178 N_SE_c_189_p N_14_c_636_n 2.31793e-19 $X=0.261 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_179 N_SE_M2_g N_14_c_639_n 3.83731e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_180 N_SE_c_191_p N_14_c_639_n 6.51345e-19 $X=0.258 $Y=0.135 $X2=0 $Y2=0
cc_181 VSS N_SE_c_135_n 2.40719e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.135
cc_182 VSS N_SE_c_137_n 5.30841e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.135
cc_183 VSS N_SE_c_154_p 9.86432e-19 $X=0.225 $Y=0.081 $X2=0.081 $Y2=0.135
cc_184 VSS N_SE_c_145_p 0.00129447f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_185 VSS N_SE_c_137_n 7.061e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_186 VSS N_SE_c_154_p 7.68051e-19 $X=0.225 $Y=0.081 $X2=0 $Y2=0
cc_187 VSS N_SE_c_135_n 8.44602e-19 $X=0.225 $Y=0.045 $X2=0.081 $Y2=0.15
cc_188 VSS N_SE_c_137_n 5.36527e-19 $X=0.337 $Y=0.045 $X2=0.081 $Y2=0.15
cc_189 VSS N_SE_c_142_p 0.00141783f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_190 VSS N_SE_c_142_p 2.35788e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_191 VSS N_SE_c_137_n 6.93145e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_192 VSS N_SE_c_142_p 9.13621e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_193 VSS N_SE_c_142_p 4.6862e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_194 VSS N_SE_c_142_p 5.41611e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_195 VSS N_SE_c_142_p 8.51044e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_196 VSS N_SE_c_207_p 0.00129447f $X=0.279 $Y=0.135 $X2=0 $Y2=0
cc_197 VSS N_SE_c_137_n 3.48715e-19 $X=0.337 $Y=0.045 $X2=0 $Y2=0
cc_198 VSS N_SE_c_159_p 9.77595e-19 $X=0.225 $Y=0.099 $X2=0 $Y2=0
cc_199 VSS N_SE_c_142_p 2.40178e-19 $X=1.175 $Y=0.045 $X2=0.081 $Y2=0.135
cc_200 VSS N_SE_c_142_p 6.42719e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_201 VSS N_SE_c_142_p 0.00110738f $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_202 N_SE_c_141_p N_QN_c_686_n 8.3796e-19 $X=1.215 $Y=0.045 $X2=0 $Y2=0
cc_203 N_SE_c_142_p N_20_c_714_n 4.98441e-19 $X=1.175 $Y=0.045 $X2=0 $Y2=0
cc_204 N_6_M3_g N_D_M4_g 0.00304756f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_205 N_6_c_218_n N_D_c_289_n 9.71463e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_206 N_6_c_215_n D 3.33994e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_207 N_6_c_224_n D 0.00195518f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_208 N_6_c_229_n D 9.77589e-19 $X=0.351 $Y=0.126 $X2=0 $Y2=0
cc_209 N_6_M3_g N_SI_M5_g 2.48122e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_210 N_6_c_215_n SI 3.40688e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_211 N_6_c_215_n N_9_c_342_n 3.98881e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_212 N_6_c_215_n N_9_c_351_n 0.0176151f $X=0.9 $Y=0.081 $X2=0.018 $Y2=0.207
cc_213 N_6_c_224_n N_9_c_351_n 0.00113948f $X=0.351 $Y=0.135 $X2=0.018 $Y2=0.207
cc_214 N_6_c_215_n N_10_c_420_n 5.04077e-19 $X=0.9 $Y=0.081 $X2=0.945 $Y2=0.178
cc_215 N_6_c_215_n N_10_c_421_n 2.53924e-19 $X=0.9 $Y=0.081 $X2=0.945 $Y2=0.178
cc_216 N_6_c_215_n N_10_c_418_n 8.29294e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_217 N_6_c_215_n N_10_c_423_n 5.75824e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_218 N_6_c_215_n N_10_c_416_n 7.91051e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_219 N_6_c_215_n N_11_c_477_n 4.20387e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_220 N_6_c_215_n N_11_c_458_n 4.92006e-19 $X=0.9 $Y=0.081 $X2=0.071 $Y2=0.054
cc_221 N_6_c_215_n N_11_c_459_n 7.19039e-19 $X=0.9 $Y=0.081 $X2=0.056 $Y2=0.054
cc_222 N_6_c_219_n N_12_c_529_n 0.00122694f $X=1.19 $Y=0.0675 $X2=0.567
+ $Y2=0.2025
cc_223 N_6_c_249_p N_12_c_529_n 2.40393e-19 $X=1.161 $Y=0.081 $X2=0.567
+ $Y2=0.2025
cc_224 N_6_c_222_n N_12_c_531_n 4.63408e-19 $X=1.19 $Y=0.2025 $X2=0 $Y2=0
cc_225 N_6_c_249_p N_12_c_523_n 9.95523e-19 $X=1.161 $Y=0.081 $X2=0.837
+ $Y2=0.0405
cc_226 N_6_c_219_n N_12_c_524_n 9.66531e-19 $X=1.19 $Y=0.0675 $X2=0.837
+ $Y2=0.178
cc_227 N_6_c_225_n N_12_c_524_n 0.00241878f $X=1.161 $Y=0.049 $X2=0.837
+ $Y2=0.178
cc_228 N_6_c_254_p N_12_c_535_n 0.00241878f $X=1.17 $Y=0.234 $X2=0 $Y2=0
cc_229 N_6_c_249_p N_12_c_528_n 0.0012739f $X=1.161 $Y=0.081 $X2=0 $Y2=0
cc_230 N_6_c_256_p N_12_c_528_n 0.00241878f $X=1.161 $Y=0.2125 $X2=0 $Y2=0
cc_231 N_6_c_257_p N_12_c_538_n 0.00241878f $X=1.161 $Y=0.225 $X2=0 $Y2=0
cc_232 N_6_c_216_n N_13_c_569_n 6.23859e-19 $X=0.936 $Y=0.081 $X2=0.056
+ $Y2=0.054
cc_233 N_6_c_249_p N_13_c_572_n 3.66836e-19 $X=1.161 $Y=0.081 $X2=0 $Y2=0
cc_234 N_6_c_249_p N_13_c_559_n 5.24665e-19 $X=1.161 $Y=0.081 $X2=0.018
+ $Y2=0.045
cc_235 N_6_c_216_n N_13_c_562_n 3.12147e-19 $X=0.936 $Y=0.081 $X2=0 $Y2=0
cc_236 N_6_c_219_n N_13_c_574_n 2.31667e-19 $X=1.19 $Y=0.0675 $X2=0.567
+ $Y2=0.135
cc_237 N_6_c_263_p N_13_c_574_n 2.53206e-19 $X=1.179 $Y=0.234 $X2=0.567
+ $Y2=0.135
cc_238 N_6_c_249_p N_13_c_574_n 0.00813033f $X=1.161 $Y=0.081 $X2=0.567
+ $Y2=0.135
cc_239 N_6_c_225_n N_13_c_574_n 0.00109426f $X=1.161 $Y=0.049 $X2=0.567
+ $Y2=0.135
cc_240 N_6_c_222_n N_13_c_575_n 3.0124e-19 $X=1.19 $Y=0.2025 $X2=0.567 $Y2=0.135
cc_241 N_6_c_267_p N_13_c_575_n 2.53206e-19 $X=1.188 $Y=0.234 $X2=0.567
+ $Y2=0.135
cc_242 N_6_M3_g N_14_c_644_n 2.37298e-19 $X=0.351 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_243 VSS N_6_c_215_n 3.90811e-19 $X=0.9 $Y=0.081 $X2=0.567 $Y2=0.2025
cc_244 VSS N_6_c_228_n 7.35661e-19 $X=0.351 $Y=0.099 $X2=0.567 $Y2=0.2025
cc_245 VSS N_6_c_271_p 6.42252e-19 $X=0.351 $Y=0.081 $X2=0 $Y2=0
cc_246 VSS N_6_c_271_p 0.00369658f $X=0.351 $Y=0.081 $X2=0.837 $Y2=0.0405
cc_247 N_6_M3_g N_16_c_668_n 2.50526e-19 $X=0.351 $Y=0.0675 $X2=0.837 $Y2=0.0405
cc_248 N_6_c_224_n N_16_c_668_n 0.00110314f $X=0.351 $Y=0.135 $X2=0.837
+ $Y2=0.0405
cc_249 VSS N_6_c_228_n 2.30452e-19 $X=0.351 $Y=0.099 $X2=0.135 $Y2=0.135
cc_250 VSS N_6_c_215_n 7.92007e-19 $X=0.9 $Y=0.081 $X2=0.675 $Y2=0.0405
cc_251 VSS N_6_c_271_p 8.14481e-19 $X=0.351 $Y=0.081 $X2=0.675 $Y2=0.178
cc_252 VSS N_6_c_215_n 2.67459e-19 $X=0.9 $Y=0.081 $X2=0.675 $Y2=0.178
cc_253 VSS N_6_c_215_n 3.16736e-19 $X=0.9 $Y=0.081 $X2=0 $Y2=0
cc_254 VSS N_6_c_215_n 2.43408e-19 $X=0.9 $Y=0.081 $X2=0.837 $Y2=0.0405
cc_255 VSS N_6_c_215_n 5.19239e-19 $X=0.9 $Y=0.081 $X2=0.837 $Y2=0.178
cc_256 N_6_c_222_n N_QN_c_687_n 2.39643e-19 $X=1.19 $Y=0.2025 $X2=0.675
+ $Y2=0.0405
cc_257 N_6_c_219_n N_QN_c_688_n 2.66287e-19 $X=1.19 $Y=0.0675 $X2=0.837
+ $Y2=0.178
cc_258 N_6_c_267_p N_QN_c_689_n 2.75088e-19 $X=1.188 $Y=0.234 $X2=0 $Y2=0
cc_259 N_6_c_216_n N_20_c_714_n 5.02041e-19 $X=0.936 $Y=0.081 $X2=0.567
+ $Y2=0.1355
cc_260 VSS N_6_c_271_p 2.73492e-19 $X=0.351 $Y=0.081 $X2=0.135 $Y2=0.054
cc_261 N_D_M4_g N_SI_M5_g 0.00348334f $X=0.405 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_262 D SI 7.00288e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_263 N_D_c_289_n N_SI_c_310_n 0.00109838f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_264 D N_9_c_351_n 0.00102191f $X=0.405 $Y=0.134 $X2=0.018 $Y2=0.207
cc_265 N_D_M4_g N_14_c_644_n 2.37298e-19 $X=0.405 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_266 VSS N_D_M4_g 3.08888e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_267 VSS D 5.77345e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_268 N_D_M4_g N_16_c_671_n 2.43567e-19 $X=0.405 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_269 D N_16_c_671_n 0.00108212f $X=0.405 $Y=0.134 $X2=0.837 $Y2=0.178
cc_270 D N_16_c_672_n 3.4434e-19 $X=0.405 $Y=0.134 $X2=0.837 $Y2=0.178
cc_271 VSS D 8.86227e-19 $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.135
cc_272 VSS D 0.00161923f $X=0.405 $Y=0.134 $X2=0.675 $Y2=0.178
cc_273 SI N_9_c_351_n 0.00138386f $X=0.473 $Y=0.135 $X2=0.018 $Y2=0.207
cc_274 SI N_14_c_637_n 0.00560919f $X=0.473 $Y=0.135 $X2=0 $Y2=0
cc_275 SI N_14_c_647_n 0.00167456f $X=0.473 $Y=0.135 $X2=0.837 $Y2=0.0405
cc_276 N_SI_M5_g N_14_c_640_n 2.70361e-19 $X=0.459 $Y=0.0675 $X2=0.837 $Y2=0.178
cc_277 SI N_16_c_666_n 6.69571e-19 $X=0.473 $Y=0.135 $X2=0.675 $Y2=0.178
cc_278 VSS N_SI_M5_g 3.10987e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_279 VSS N_SI_c_310_n 2.08525e-19 $X=0.475 $Y=0.135 $X2=0 $Y2=0
cc_280 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.837 $Y2=0.0405
cc_281 VSS SI 5.41556e-19 $X=0.473 $Y=0.135 $X2=0.837 $Y2=0.0405
cc_282 VSS SI 0.00110314f $X=0.473 $Y=0.135 $X2=0 $Y2=0
cc_283 N_9_M6_g N_10_M8_g 2.82885e-19 $X=0.621 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_284 N_9_c_366_n N_10_c_410_n 5.29207e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_285 N_9_c_355_n N_10_c_411_n 0.00318254f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_286 N_9_c_350_n N_10_c_412_n 0.00128311f $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_287 N_9_M11_g N_11_M9_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_288 N_9_c_334_n N_11_c_485_n 2.98891e-19 $X=0.891 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_289 N_9_c_346_n N_11_c_453_n 3.24488e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_290 N_9_M6_g N_11_c_487_n 3.41974e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_291 N_9_c_346_n N_11_c_487_n 0.00102727f $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_292 N_9_c_342_n N_11_c_489_n 0.00133841f $X=0.621 $Y=0.135 $X2=0 $Y2=0
cc_293 N_9_c_351_n N_11_c_490_n 7.726e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_294 N_9_c_346_n N_11_c_460_n 8.63476e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_295 N_9_c_351_n N_11_c_460_n 5.92766e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_296 N_9_c_351_n N_11_c_472_n 3.70527e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_297 N_9_c_366_n N_11_c_473_n 3.70527e-19 $X=0.817 $Y=0.153 $X2=0 $Y2=0
cc_298 N_9_M11_g N_12_M12_g 2.82885e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_299 N_9_M11_g N_13_c_570_n 3.18506e-19 $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_300 N_9_c_355_n N_13_c_570_n 4.09234e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_301 N_9_c_355_n N_13_c_590_n 0.00320381f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_302 N_9_c_355_n N_13_c_563_n 3.56772e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_303 N_9_c_350_n N_13_c_574_n 9.40125e-19 $X=0.891 $Y=0.153 $X2=0 $Y2=0
cc_304 N_9_c_335_n N_14_c_636_n 0.0010034f $X=0.16 $Y=0.216 $X2=0.081 $Y2=0.135
cc_305 N_9_c_344_n N_14_c_636_n 0.00105265f $X=0.189 $Y=0.153 $X2=0.081
+ $Y2=0.135
cc_306 N_9_c_351_n N_14_c_637_n 4.24134e-19 $X=0.743 $Y=0.153 $X2=0 $Y2=0
cc_307 N_9_c_337_n N_14_c_639_n 7.83928e-19 $X=0.18 $Y=0.234 $X2=0 $Y2=0
cc_308 VSS N_9_c_400_p 9.30745e-19 $X=0.16 $Y=0.054 $X2=0.081 $Y2=0.135
cc_309 N_10_M8_g N_11_M9_g 0.00268443f $X=0.729 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_310 N_10_c_418_n N_11_M9_g 3.7702e-19 $X=0.792 $Y=0.09 $X2=0.135 $Y2=0.054
cc_311 N_10_c_419_n N_11_c_480_n 2.46574e-19 $X=0.81 $Y=0.054 $X2=0 $Y2=0
cc_312 N_10_c_420_n N_11_c_498_n 0.00360624f $X=0.747 $Y=0.09 $X2=0 $Y2=0
cc_313 N_10_c_421_n N_11_c_458_n 3.99428e-19 $X=0.747 $Y=0.09 $X2=0.071
+ $Y2=0.054
cc_314 N_10_c_412_n N_11_c_490_n 2.22221e-19 $X=0.837 $Y=0.165 $X2=0.056
+ $Y2=0.216
cc_315 N_10_c_435_p N_11_c_466_n 2.22221e-19 $X=0.837 $Y=0.225 $X2=0.018
+ $Y2=0.045
cc_316 N_10_c_418_n N_11_c_471_n 0.00205899f $X=0.792 $Y=0.09 $X2=0.018
+ $Y2=0.198
cc_317 N_10_c_437_p N_11_c_471_n 7.38434e-19 $X=0.837 $Y=0.14 $X2=0.018
+ $Y2=0.198
cc_318 N_10_M8_g N_11_c_473_n 3.21351e-19 $X=0.729 $Y=0.0405 $X2=0.018 $Y2=0.216
cc_319 N_10_c_420_n N_11_c_473_n 0.00205899f $X=0.747 $Y=0.09 $X2=0.018
+ $Y2=0.216
cc_320 N_10_c_405_n N_13_c_556_n 0.00379158f $X=0.81 $Y=0.0405 $X2=0 $Y2=0
cc_321 N_10_c_419_n N_13_c_556_n 2.84891e-19 $X=0.81 $Y=0.054 $X2=0 $Y2=0
cc_322 N_10_c_416_n N_13_c_556_n 2.08929e-19 $X=0.837 $Y=0.09 $X2=0 $Y2=0
cc_323 N_10_c_408_n N_13_c_558_n 0.00222825f $X=0.866 $Y=0.2295 $X2=0 $Y2=0
cc_324 N_10_c_405_n N_13_c_569_n 3.41768e-19 $X=0.81 $Y=0.0405 $X2=0.056
+ $Y2=0.054
cc_325 N_10_c_416_n N_13_c_559_n 4.2911e-19 $X=0.837 $Y=0.09 $X2=0.018 $Y2=0.045
cc_326 N_10_c_414_n N_13_c_561_n 4.2911e-19 $X=0.837 $Y=0.207 $X2=0.018
+ $Y2=0.198
cc_327 N_10_c_408_n N_13_c_562_n 3.64454e-19 $X=0.866 $Y=0.2295 $X2=0 $Y2=0
cc_328 N_10_c_410_n N_13_c_562_n 4.86017e-19 $X=0.828 $Y=0.234 $X2=0 $Y2=0
cc_329 N_10_c_449_p N_13_c_563_n 4.2911e-19 $X=0.837 $Y=0.101 $X2=0 $Y2=0
cc_330 N_11_c_453_n N_14_c_637_n 0.00424458f $X=0.594 $Y=0.2025 $X2=0 $Y2=0
cc_331 N_11_c_455_n N_14_c_637_n 4.3429e-19 $X=0.595 $Y=0.234 $X2=0 $Y2=0
cc_332 N_11_c_455_n N_14_c_647_n 2.8677e-19 $X=0.595 $Y=0.234 $X2=0.837
+ $Y2=0.0405
cc_333 VSS N_11_c_453_n 0.0016174f $X=0.594 $Y=0.2025 $X2=0.567 $Y2=0.1355
cc_334 VSS N_11_c_477_n 0.00414127f $X=0.648 $Y=0.036 $X2=0.567 $Y2=0.1355
cc_335 VSS N_11_c_478_n 3.30384e-19 $X=0.649 $Y=0.036 $X2=0.567 $Y2=0.1355
cc_336 VSS N_11_c_477_n 2.79363e-19 $X=0.648 $Y=0.036 $X2=0.675 $Y2=0.0405
cc_337 VSS N_11_c_458_n 2.70508e-19 $X=0.693 $Y=0.081 $X2=0.675 $Y2=0.0405
cc_338 N_11_c_453_n N_19_c_705_n 0.00167238f $X=0.594 $Y=0.2025 $X2=0.567
+ $Y2=0.1355
cc_339 N_11_c_515_p N_19_c_705_n 0.00315491f $X=0.684 $Y=0.234 $X2=0.567
+ $Y2=0.1355
cc_340 N_11_c_487_n N_19_c_705_n 0.00111131f $X=0.649 $Y=0.234 $X2=0.567
+ $Y2=0.1355
cc_341 N_11_c_477_n N_19_c_705_n 5.67227e-19 $X=0.648 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_342 N_11_c_518_p N_19_c_705_n 4.0515e-19 $X=0.693 $Y=0.225 $X2=0.567
+ $Y2=0.1355
cc_343 N_11_c_519_p N_19_c_705_n 0.0409693f $X=0.693 $Y=0.216 $X2=0.567
+ $Y2=0.1355
cc_344 N_11_c_457_n N_22_M8_s 2.44135e-19 $X=0.684 $Y=0.036 $X2=0.135 $Y2=0.054
cc_345 N_11_c_480_n N_22_M8_s 3.62465e-19 $X=0.693 $Y=0.062 $X2=0.135 $Y2=0.054
cc_346 N_12_M12_g N_13_M13_g 0.00268443f $X=0.999 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_347 N_12_c_527_n N_13_M13_g 3.55314e-19 $X=1.062 $Y=0.036 $X2=0.135 $Y2=0.054
cc_348 N_12_c_525_n N_13_c_568_n 0.00136796f $X=1.008 $Y=0.036 $X2=0 $Y2=0
cc_349 N_12_c_523_n N_13_c_572_n 0.00136796f $X=0.999 $Y=0.105 $X2=0 $Y2=0
cc_350 N_12_c_544_p N_13_c_559_n 3.34766e-19 $X=0.999 $Y=0.1055 $X2=0.018
+ $Y2=0.045
cc_351 N_12_c_523_n N_13_c_559_n 0.00136796f $X=0.999 $Y=0.105 $X2=0.018
+ $Y2=0.045
cc_352 N_12_c_535_n N_13_c_561_n 5.28703e-19 $X=1.107 $Y=0.225 $X2=0.018
+ $Y2=0.198
cc_353 N_12_M12_g N_13_c_610_n 6.35734e-19 $X=0.999 $Y=0.0405 $X2=0.027
+ $Y2=0.036
cc_354 N_12_c_523_n N_13_c_610_n 7.99759e-19 $X=0.999 $Y=0.105 $X2=0.027
+ $Y2=0.036
cc_355 N_12_c_527_n N_13_c_612_n 2.75024e-19 $X=1.062 $Y=0.036 $X2=0.054
+ $Y2=0.036
cc_356 N_12_c_538_n N_13_c_612_n 0.00266503f $X=1.107 $Y=0.171 $X2=0.054
+ $Y2=0.036
cc_357 N_12_c_531_n N_13_c_574_n 2.19627e-19 $X=1.078 $Y=0.2295 $X2=0.567
+ $Y2=0.135
cc_358 N_12_c_538_n N_13_c_574_n 0.00106087f $X=1.107 $Y=0.171 $X2=0.567
+ $Y2=0.135
cc_359 N_12_c_553_p N_13_c_574_n 5.80975e-19 $X=1.098 $Y=0.234 $X2=0.567
+ $Y2=0.135
cc_360 N_12_c_525_n N_20_c_714_n 5.06067e-19 $X=1.008 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_361 N_13_c_566_n N_QN_M16_d 3.7444e-19 $X=1.377 $Y=0.136 $X2=0.135 $Y2=0.054
cc_362 N_13_c_566_n N_QN_M34_d 3.85232e-19 $X=1.377 $Y=0.136 $X2=0 $Y2=0
cc_363 N_13_c_566_n N_QN_c_687_n 8.43851e-19 $X=1.377 $Y=0.136 $X2=0.675
+ $Y2=0.0405
cc_364 N_13_c_577_n N_QN_c_687_n 0.00133574f $X=1.269 $Y=0.136 $X2=0.675
+ $Y2=0.0405
cc_365 N_13_M16_g N_QN_c_686_n 4.61823e-19 $X=1.323 $Y=0.0675 $X2=0.837
+ $Y2=0.0405
cc_366 N_13_M17_g N_QN_c_686_n 4.61823e-19 $X=1.377 $Y=0.0675 $X2=0.837
+ $Y2=0.0405
cc_367 N_13_c_566_n N_QN_c_686_n 0.00131663f $X=1.377 $Y=0.136 $X2=0.837
+ $Y2=0.0405
cc_368 N_13_c_566_n N_QN_c_688_n 7.60428e-19 $X=1.377 $Y=0.136 $X2=0.837
+ $Y2=0.178
cc_369 N_13_c_577_n N_QN_c_688_n 6.32721e-19 $X=1.269 $Y=0.136 $X2=0.837
+ $Y2=0.178
cc_370 N_13_M16_g N_QN_c_689_n 4.56718e-19 $X=1.323 $Y=0.0675 $X2=0 $Y2=0
cc_371 N_13_M17_g N_QN_c_689_n 4.56718e-19 $X=1.377 $Y=0.0675 $X2=0 $Y2=0
cc_372 N_13_c_566_n N_QN_c_689_n 0.00134222f $X=1.377 $Y=0.136 $X2=0 $Y2=0
cc_373 N_13_c_566_n N_QN_c_702_n 3.65018e-19 $X=1.377 $Y=0.136 $X2=0 $Y2=0
cc_374 N_13_c_577_n N_QN_c_702_n 5.79504e-19 $X=1.269 $Y=0.136 $X2=0 $Y2=0
cc_375 N_13_c_556_n N_20_c_714_n 0.00210698f $X=0.864 $Y=0.0405 $X2=0.567
+ $Y2=0.1355
cc_376 N_13_c_568_n N_20_c_714_n 0.00203632f $X=0.936 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_377 N_13_c_571_n N_20_c_714_n 0.00129774f $X=0.92 $Y=0.036 $X2=0.567
+ $Y2=0.1355
cc_378 N_13_c_572_n N_20_c_714_n 0.00104094f $X=0.945 $Y=0.081 $X2=0.567
+ $Y2=0.1355
cc_379 N_13_c_635_p N_20_c_714_n 2.5109e-19 $X=0.99 $Y=0.162 $X2=0.567
+ $Y2=0.1355
cc_380 VSS N_14_c_636_n 0.00156967f $X=0.272 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_381 VSS N_14_c_637_n 0.00145872f $X=0.542 $Y=0.2025 $X2=0.675 $Y2=0.178
cc_382 N_14_c_636_n N_16_c_679_n 0.003872f $X=0.272 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_383 N_14_c_644_n N_16_c_679_n 0.00248801f $X=0.447 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_384 N_14_c_637_n N_16_c_681_n 0.00434154f $X=0.542 $Y=0.2025 $X2=0.567
+ $Y2=0.1355
cc_385 N_14_c_644_n N_16_c_681_n 0.0025506f $X=0.447 $Y=0.234 $X2=0.567
+ $Y2=0.1355
cc_386 N_14_c_636_n N_16_c_665_n 3.19827e-19 $X=0.272 $Y=0.2025 $X2=0.567
+ $Y2=0.2025
cc_387 N_14_c_644_n N_16_c_665_n 0.0113176f $X=0.447 $Y=0.234 $X2=0.567
+ $Y2=0.2025
cc_388 VSS N_14_c_637_n 4.53012e-19 $X=0.542 $Y=0.2025 $X2=0.837 $Y2=0.178
cc_389 VSS N_16_c_681_n 0.00141703f $X=0.432 $Y=0.2025 $X2=0.135 $Y2=0.135

* END of "./SDFLx3_ASAP7_75t_SRAM.pex.sp.SDFLX3_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: SDFLx4_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 13:05:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "SDFLx4_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./SDFLx4_ASAP7_75t_SRAM.pex.sp.pex"
* File: SDFLx4_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 13:05:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_SDFLX4_ASAP7_75T_SRAM%CLK 2 5 7 11 VSS
c13 11 VSS 0.00571615f $X=0.081 $Y=0.1345
c14 5 VSS 0.00203788f $X=0.081 $Y=0.135
c15 2 VSS 0.0654663f $X=0.081 $Y=0.0675
r16 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%4 2 5 7 10 13 15 18 21 23 25 30 33 36 38 41 45 46
+ 54 61 65 68 69 70 71 72 74 75 VSS
c84 114 VSS 1.06551e-19 $X=0.03 $Y=0.117
c85 113 VSS 6.89947e-19 $X=0.027 $Y=0.117
c86 75 VSS 0.00125248f $X=1.107 $Y=0.117
c87 74 VSS 0.0124661f $X=1.107 $Y=0.117
c88 72 VSS 0.00194293f $X=0.682 $Y=0.117
c89 71 VSS 0.00253628f $X=0.581 $Y=0.117
c90 70 VSS 0.00171031f $X=0.229 $Y=0.117
c91 69 VSS 0.00697398f $X=0.175 $Y=0.117
c92 68 VSS 7.51069e-19 $X=0.783 $Y=0.117
c93 65 VSS 0.00255826f $X=0.135 $Y=0.117
c94 61 VSS 6.34103e-19 $X=0.033 $Y=0.117
c95 57 VSS 2.97869e-19 $X=0.0505 $Y=0.234
c96 56 VSS 0.00199279f $X=0.047 $Y=0.234
c97 54 VSS 0.00251086f $X=0.054 $Y=0.234
c98 52 VSS 0.00305101f $X=0.027 $Y=0.234
c99 48 VSS 2.97869e-19 $X=0.0505 $Y=0.036
c100 47 VSS 0.00179897f $X=0.047 $Y=0.036
c101 46 VSS 0.00633992f $X=0.054 $Y=0.036
c102 45 VSS 0.00447521f $X=0.054 $Y=0.036
c103 43 VSS 0.00306551f $X=0.027 $Y=0.036
c104 42 VSS 5.16336e-19 $X=0.018 $Y=0.2125
c105 41 VSS 0.00321988f $X=0.018 $Y=0.2
c106 40 VSS 4.96914e-19 $X=0.018 $Y=0.225
c107 38 VSS 9.28596e-19 $X=0.018 $Y=0.0855
c108 37 VSS 7.23544e-19 $X=0.018 $Y=0.063
c109 36 VSS 9.58863e-19 $X=0.018 $Y=0.108
c110 33 VSS 0.00628074f $X=0.056 $Y=0.2025
c111 30 VSS 3.02808e-19 $X=0.071 $Y=0.2025
c112 25 VSS 2.55988e-19 $X=0.071 $Y=0.0675
c113 21 VSS 0.001261f $X=1.107 $Y=0.135
c114 18 VSS 0.0599455f $X=1.107 $Y=0.0675
c115 13 VSS 0.00144009f $X=0.783 $Y=0.135
c116 10 VSS 0.0633669f $X=0.783 $Y=0.0675
c117 5 VSS 0.00185078f $X=0.135 $Y=0.135
c118 2 VSS 0.0641982f $X=0.135 $Y=0.0675
r119 113 114 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.117 $X2=0.03 $Y2=0.117
r120 110 113 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.117 $X2=0.027 $Y2=0.117
r121 74 75 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.107 $Y=0.117 $X2=1.107
+ $Y2=0.117
r122 71 72 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M2 $thickness=3.6e-08 $X=0.581
+ $Y=0.117 $X2=0.682 $Y2=0.117
r123 70 71 23.9012 $w=1.8e-08 $l=3.52e-07 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.117 $X2=0.581 $Y2=0.117
r124 69 70 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.175
+ $Y=0.117 $X2=0.229 $Y2=0.117
r125 67 74 22 $w=1.8e-08 $l=3.24e-07 $layer=M2 $thickness=3.6e-08 $X=0.783
+ $Y=0.117 $X2=1.107 $Y2=0.117
r126 67 72 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M2 $thickness=3.6e-08 $X=0.783
+ $Y=0.117 $X2=0.682 $Y2=0.117
r127 67 68 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.783 $Y=0.117 $X2=0.783
+ $Y2=0.117
r128 64 69 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.117 $X2=0.175 $Y2=0.117
r129 64 65 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.135 $Y=0.117 $X2=0.135
+ $Y2=0.117
r130 61 114 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.117 $X2=0.03 $Y2=0.117
r131 60 64 6.92593 $w=1.8e-08 $l=1.02e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.117 $X2=0.135 $Y2=0.117
r132 60 61 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.117 $X2=0.033
+ $Y2=0.117
r133 56 57 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r134 54 57 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r135 52 56 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r136 47 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r137 45 48 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r138 45 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r139 43 47 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r140 41 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r141 40 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r142 40 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r143 39 110 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.117
r144 39 41 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.2
r145 37 38 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.0855
r146 36 110 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.108 $X2=0.018 $Y2=0.117
r147 36 38 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.108 $X2=0.018 $Y2=0.0855
r148 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r149 35 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r150 33 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r151 30 33 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r152 28 46 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.054 $Y=0.0675 $X2=0.054 $Y2=0.036
r153 25 28 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r154 21 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.107 $Y=0.135 $X2=1.107
+ $Y2=0.135
r155 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.135 $X2=1.107 $Y2=0.2025
r156 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.0675 $X2=1.107 $Y2=0.135
r157 13 68 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.135 $X2=0.783
+ $Y2=0.135
r158 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.135 $X2=0.783 $Y2=0.2025
r159 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.135
r160 5 65 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r161 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r162 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%SE 2 5 7 10 13 15 21 31 39 42 43 51 57 58 VSS
c56 58 VSS 6.15152e-20 $X=0.567 $Y=0.1205
c57 57 VSS 0.00112348f $X=0.567 $Y=0.106
c58 51 VSS 1.82947e-19 $X=0.567 $Y=0.135
c59 43 VSS 0.00116134f $X=0.567 $Y=0.081
c60 42 VSS 0.00971257f $X=0.567 $Y=0.081
c61 39 VSS 0.00947346f $X=0.243 $Y=0.081
c62 31 VSS 0.0100986f $X=0.243 $Y=0.135
c63 23 VSS 1.33806e-20 $X=0.2745 $Y=0.135
c64 22 VSS 0.00149043f $X=0.271 $Y=0.135
c65 21 VSS 1.85952e-19 $X=0.278 $Y=0.1345
c66 13 VSS 0.00121878f $X=0.567 $Y=0.135
c67 10 VSS 0.0587511f $X=0.567 $Y=0.0675
c68 5 VSS 0.00645728f $X=0.297 $Y=0.135
c69 2 VSS 0.070241f $X=0.297 $Y=0.0675
r70 57 58 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.106 $X2=0.567 $Y2=0.1205
r71 51 58 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.1205
r72 43 57 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.567 $Y2=0.106
r73 42 43 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.567 $Y=0.081 $X2=0.567
+ $Y2=0.081
r74 38 42 22 $w=1.8e-08 $l=3.24e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.081 $X2=0.567 $Y2=0.081
r75 38 39 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.081 $X2=0.243
+ $Y2=0.081
r76 30 39 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.081
r77 30 31 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.135
r78 22 23 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.271
+ $Y=0.135 $X2=0.2745 $Y2=0.135
r79 21 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.28 $Y=0.135 $X2=0.28
+ $Y2=0.135
r80 21 23 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.278
+ $Y=0.135 $X2=0.2745 $Y2=0.135
r81 19 31 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.243 $Y2=0.135
r82 19 22 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.271 $Y2=0.135
r83 13 51 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r84 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r85 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r86 5 25 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.28 $Y2=0.135
r87 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r88 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%D 2 5 7 24 VSS
c23 24 VSS 0.0118434f $X=0.459 $Y=0.1345
c24 5 VSS 0.00185098f $X=0.459 $Y=0.135
c25 2 VSS 0.0629574f $X=0.459 $Y=0.0675
r26 5 24 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r27 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r28 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%7 2 5 7 9 14 17 20 22 23 24 25 26 27 29 30 31 32
+ 35 37 38 42 44 45 52 53 56 VSS
c54 56 VSS 1.61802e-19 $X=0.351 $Y=0.072
c55 53 VSS 0.00367986f $X=0.342 $Y=0.234
c56 52 VSS 0.00194932f $X=0.351 $Y=0.234
c57 45 VSS 0.0036746f $X=0.342 $Y=0.036
c58 44 VSS 0.00199758f $X=0.351 $Y=0.036
c59 42 VSS 0.00774747f $X=0.324 $Y=0.036
c60 38 VSS 2.76819e-19 $X=0.513 $Y=0.117
c61 37 VSS 4.68887e-19 $X=0.513 $Y=0.099
c62 35 VSS 2.69498e-19 $X=0.513 $Y=0.135
c63 32 VSS 4.17962e-19 $X=0.486 $Y=0.072
c64 31 VSS 3.38584e-20 $X=0.468 $Y=0.072
c65 30 VSS 0.00175333f $X=0.418 $Y=0.072
c66 29 VSS 8.4059e-19 $X=0.378 $Y=0.072
c67 27 VSS 6.46578e-19 $X=0.504 $Y=0.072
c68 26 VSS 5.547e-19 $X=0.351 $Y=0.1845
c69 25 VSS 1.96258e-19 $X=0.351 $Y=0.144
c70 24 VSS 5.16212e-19 $X=0.351 $Y=0.126
c71 23 VSS 3.64391e-19 $X=0.351 $Y=0.099
c72 22 VSS 5.81348e-19 $X=0.351 $Y=0.225
c73 20 VSS 4.51561e-19 $X=0.351 $Y=0.063
c74 17 VSS 0.00759509f $X=0.322 $Y=0.2025
c75 12 VSS 3.78024e-19 $X=0.322 $Y=0.0675
c76 5 VSS 0.00134234f $X=0.513 $Y=0.135
c77 2 VSS 0.0585448f $X=0.513 $Y=0.0675
r78 53 54 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.3465 $Y2=0.234
r79 52 54 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.234 $X2=0.3465 $Y2=0.234
r80 49 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.342 $Y2=0.234
r81 45 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.3465 $Y2=0.036
r82 44 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.036 $X2=0.3465 $Y2=0.036
r83 41 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r84 41 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r85 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.099 $X2=0.513 $Y2=0.117
r86 35 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.117
r87 33 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.081 $X2=0.513 $Y2=0.099
r88 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.072 $X2=0.486 $Y2=0.072
r89 30 31 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.072 $X2=0.468 $Y2=0.072
r90 29 30 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.418 $Y2=0.072
r91 28 56 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.072 $X2=0.351 $Y2=0.072
r92 28 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.072 $X2=0.378 $Y2=0.072
r93 27 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.072 $X2=0.513 $Y2=0.081
r94 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.072 $X2=0.486 $Y2=0.072
r95 25 26 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.144 $X2=0.351 $Y2=0.1845
r96 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.144
r97 23 24 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.099 $X2=0.351 $Y2=0.126
r98 22 52 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.234
r99 22 26 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.1845
r100 21 56 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.072
r101 21 23 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.099
r102 20 56 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.063 $X2=0.351 $Y2=0.072
r103 19 44 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.036
r104 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.063
r105 17 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r106 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.322 $Y2=0.2025
r107 12 42 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r108 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.322 $Y2=0.0675
r109 5 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r110 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r111 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%SI 2 5 7 11 VSS
c26 11 VSS 0.0106807f $X=0.621 $Y=0.1345
c27 5 VSS 0.00120269f $X=0.621 $Y=0.135
c28 2 VSS 0.0596457f $X=0.621 $Y=0.0675
r29 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r30 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r31 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%9 2 8 11 14 17 20 23 25 30 33 35 37 38 47 48 54 66
+ 68 69 74 75 79 84 89 100 101 102 103 VSS
c124 105 VSS 1.0884e-19 $X=0.189 $Y=0.2125
c125 103 VSS 4.06956e-19 $X=0.189 $Y=0.128
c126 102 VSS 4.95407e-19 $X=0.189 $Y=0.103
c127 101 VSS 2.10509e-19 $X=0.189 $Y=0.081
c128 100 VSS 1.53051e-19 $X=0.189 $Y=0.063
c129 89 VSS 6.93139e-19 $X=1.161 $Y=0.135
c130 84 VSS 0.00122127f $X=1.053 $Y=0.135
c131 79 VSS 0.00146217f $X=0.837 $Y=0.135
c132 75 VSS 0.00122905f $X=0.693 $Y=0.135
c133 74 VSS 0.00324557f $X=0.693 $Y=0.135
c134 69 VSS 6.85269e-19 $X=1.141 $Y=0.153
c135 68 VSS 0.0221225f $X=1.121 $Y=0.153
c136 66 VSS 0.00121091f $X=1.161 $Y=0.153
c137 54 VSS 0.00100048f $X=0.189 $Y=0.153
c138 48 VSS 0.00383164f $X=0.18 $Y=0.234
c139 47 VSS 4.95331e-19 $X=0.189 $Y=0.225
c140 46 VSS 0.00196236f $X=0.189 $Y=0.234
c141 38 VSS 0.00853777f $X=0.162 $Y=0.036
c142 37 VSS 0.00301835f $X=0.162 $Y=0.036
c143 35 VSS 0.00516266f $X=0.18 $Y=0.036
c144 33 VSS 0.00868282f $X=0.16 $Y=0.2025
c145 28 VSS 2.55988e-19 $X=0.16 $Y=0.0675
c146 23 VSS 8.78735e-19 $X=1.161 $Y=0.135
c147 20 VSS 0.0586114f $X=1.161 $Y=0.0675
c148 14 VSS 0.0642113f $X=1.053 $Y=0.135
c149 8 VSS 0.0600934f $X=0.837 $Y=0.135
c150 2 VSS 0.0644358f $X=0.675 $Y=0.0675
r151 104 105 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.2 $X2=0.189 $Y2=0.2125
r152 102 103 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.103 $X2=0.189 $Y2=0.128
r153 101 102 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.081 $X2=0.189 $Y2=0.103
r154 100 101 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.063 $X2=0.189 $Y2=0.081
r155 74 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.693 $Y=0.135 $X2=0.693
+ $Y2=0.135
r156 68 69 1.35802 $w=1.8e-08 $l=2e-08 $layer=M2 $thickness=3.6e-08 $X=1.121
+ $Y=0.153 $X2=1.141 $Y2=0.153
r157 66 69 1.35802 $w=1.8e-08 $l=2e-08 $layer=M2 $thickness=3.6e-08 $X=1.161
+ $Y=0.153 $X2=1.141 $Y2=0.153
r158 66 89 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.161 $Y=0.153 $X2=1.161
+ $Y2=0.153
r159 63 68 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=1.053
+ $Y=0.153 $X2=1.121 $Y2=0.153
r160 63 84 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.053 $Y=0.153 $X2=1.053
+ $Y2=0.153
r161 60 63 14.6667 $w=1.8e-08 $l=2.16e-07 $layer=M2 $thickness=3.6e-08 $X=0.837
+ $Y=0.153 $X2=1.053 $Y2=0.153
r162 60 79 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.837 $Y=0.153 $X2=0.837
+ $Y2=0.153
r163 57 60 9.77778 $w=1.8e-08 $l=1.44e-07 $layer=M2 $thickness=3.6e-08 $X=0.693
+ $Y=0.153 $X2=0.837 $Y2=0.153
r164 57 75 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.693 $Y=0.153 $X2=0.693
+ $Y2=0.153
r165 54 104 3.19136 $w=1.8e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.2
r166 54 103 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.128
r167 53 57 34.2222 $w=1.8e-08 $l=5.04e-07 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.693 $Y2=0.153
r168 53 54 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.153 $X2=0.189
+ $Y2=0.153
r169 51 100 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r170 48 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r171 47 105 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.225 $X2=0.189 $Y2=0.2125
r172 46 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r173 46 47 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.189 $Y2=0.225
r174 43 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r175 37 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r176 35 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r177 35 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.162 $Y2=0.036
r178 33 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r179 30 33 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.16 $Y2=0.2025
r180 28 38 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.162 $Y=0.0675 $X2=0.162 $Y2=0.036
r181 25 28 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.16 $Y2=0.0675
r182 23 89 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.161 $Y=0.135 $X2=1.161
+ $Y2=0.135
r183 20 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.161 $Y=0.0675 $X2=1.161 $Y2=0.135
r184 14 84 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.053 $Y=0.135 $X2=1.053
+ $Y2=0.135
r185 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.135 $X2=1.053 $Y2=0.2025
r186 8 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.135 $X2=0.837
+ $Y2=0.135
r187 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.2025
r188 5 74 16.3636 $w=2.2e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.693 $Y2=0.135
r189 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0675 $X2=0.675 $Y2=0.135
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%10 4 7 9 11 16 19 21 26 29 33 36 38 40 42 43 49
+ VSS
c37 49 VSS 0.0362427f $X=0.999 $Y=0.162
c38 43 VSS 5.31938e-19 $X=0.954 $Y=0.072
c39 42 VSS 0.00378458f $X=0.936 $Y=0.072
c40 40 VSS 0.001558f $X=0.972 $Y=0.072
c41 38 VSS 8.97194e-19 $X=0.9 $Y=0.072
c42 36 VSS 6.15152e-20 $X=0.891 $Y=0.1205
c43 35 VSS 0.00121732f $X=0.891 $Y=0.106
c44 33 VSS 3.0794e-19 $X=0.891 $Y=0.135
c45 29 VSS 0.0225573f $X=1.028 $Y=0.2025
c46 26 VSS 3.25039e-19 $X=1.043 $Y=0.2025
c47 19 VSS 0.0555224f $X=1.082 $Y=0.0675
c48 16 VSS 3.25039e-19 $X=1.097 $Y=0.0675
c49 14 VSS 3.34937e-19 $X=0.97 $Y=0.0675
c50 7 VSS 0.00125164f $X=0.891 $Y=0.135
c51 4 VSS 0.0584835f $X=0.891 $Y=0.0675
r52 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.072 $X2=0.954 $Y2=0.072
r53 40 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.072 $X2=0.954 $Y2=0.072
r54 38 42 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.072 $X2=0.936 $Y2=0.072
r55 35 36 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.106 $X2=0.891 $Y2=0.1205
r56 33 36 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.135 $X2=0.891 $Y2=0.1205
r57 31 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.891 $Y=0.081 $X2=0.9 $Y2=0.072
r58 31 35 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.081 $X2=0.891 $Y2=0.106
r59 29 49 14.4321 $w=7.8e-08 $l=4.05e-08 $layer=LISD $thickness=2.8e-08 $X=0.999
+ $Y=0.2025 $X2=0.999 $Y2=0.162
r60 26 29 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.043 $Y=0.2025 $X2=1.028 $Y2=0.2025
r61 21 29 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.2025 $X2=0.97 $Y2=0.2025
r62 19 53 21.3536 $w=8.1e-08 $l=8.35e-08 $layer=LISD $thickness=2.8e-08 $X=1.082
+ $Y=0.0675 $X2=0.9985 $Y2=0.0675
r63 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.097 $Y=0.0675 $X2=1.082 $Y2=0.0675
r64 14 53 7.28836 $w=8.1e-08 $l=2.85e-08 $layer=LISD $thickness=2.8e-08 $X=0.97
+ $Y=0.0675 $X2=0.9985 $Y2=0.0675
r65 14 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.072 $X2=0.972
+ $Y2=0.072
r66 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.0675 $X2=0.97 $Y2=0.0675
r67 7 33 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.135 $X2=0.891
+ $Y2=0.135
r68 7 9 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.135 $X2=0.891 $Y2=0.2025
r69 4 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.0675 $X2=0.891 $Y2=0.135
r70 1 53 7.09296 $w=8.1e-08 $l=4.05e-08 $layer=LISD $thickness=2.8e-08 $X=0.9985
+ $Y=0.108 $X2=0.9985 $Y2=0.0675
r71 1 49 24.8571 $w=4.5e-08 $l=5.4e-08 $layer=LISD $thickness=2.8e-08 $X=0.9985
+ $Y=0.108 $X2=0.9985 $Y2=0.162
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%11 2 5 7 9 14 17 19 20 23 24 26 32 33 34 35 36 37
+ 38 40 46 47 49 50 51 54 59 VSS
c59 60 VSS 4.719e-19 $X=0.945 $Y=0.2
c60 59 VSS 0.00101748f $X=0.945 $Y=0.189
c61 58 VSS 1.48656e-19 $X=0.945 $Y=0.167
c62 54 VSS 2.26463e-19 $X=0.945 $Y=0.135
c63 52 VSS 0.00105105f $X=0.945 $Y=0.225
c64 51 VSS 0.00146362f $X=0.9 $Y=0.234
c65 50 VSS 0.00363455f $X=0.882 $Y=0.234
c66 49 VSS 0.0014995f $X=0.846 $Y=0.234
c67 48 VSS 0.00101201f $X=0.828 $Y=0.234
c68 47 VSS 0.0020447f $X=0.819 $Y=0.234
c69 46 VSS 0.00805618f $X=0.936 $Y=0.234
c70 40 VSS 5.31938e-19 $X=0.792 $Y=0.198
c71 39 VSS 2.07422e-19 $X=0.774 $Y=0.198
c72 38 VSS 4.09554e-20 $X=0.77 $Y=0.198
c73 37 VSS 8.20366e-20 $X=0.767 $Y=0.198
c74 36 VSS 6.34818e-19 $X=0.756 $Y=0.198
c75 35 VSS 5.99287e-19 $X=0.801 $Y=0.198
c76 34 VSS 2.66851e-19 $X=0.747 $Y=0.178
c77 33 VSS 1.28225e-19 $X=0.747 $Y=0.167
c78 32 VSS 9.95178e-19 $X=0.747 $Y=0.164
c79 26 VSS 4.68208e-19 $X=0.747 $Y=0.09
c80 24 VSS 2.54721e-19 $X=0.747 $Y=0.189
c81 23 VSS 0.00346721f $X=0.81 $Y=0.2025
c82 19 VSS 6.04398e-19 $X=0.827 $Y=0.2025
c83 17 VSS 0.0144192f $X=0.758 $Y=0.0675
c84 14 VSS 3.25039e-19 $X=0.773 $Y=0.0675
c85 12 VSS 6.23621e-19 $X=0.7 $Y=0.0675
c86 5 VSS 0.0014001f $X=0.945 $Y=0.135
c87 2 VSS 0.0619707f $X=0.945 $Y=0.0675
r88 59 60 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.189 $X2=0.945 $Y2=0.2
r89 58 59 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.167 $X2=0.945 $Y2=0.189
r90 57 58 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.164 $X2=0.945 $Y2=0.167
r91 54 57 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.135 $X2=0.945 $Y2=0.164
r92 52 60 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.2
r93 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.234 $X2=0.9 $Y2=0.234
r94 49 50 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.234 $X2=0.882 $Y2=0.234
r95 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.846 $Y2=0.234
r96 47 48 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.819
+ $Y=0.234 $X2=0.828 $Y2=0.234
r97 46 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r98 46 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.9 $Y2=0.234
r99 42 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.81 $Y=0.225 $X2=0.819 $Y2=0.234
r100 42 44 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.225 $X2=0.81 $Y2=0.216
r101 41 44 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.207 $X2=0.81 $Y2=0.216
r102 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.198 $X2=0.792 $Y2=0.198
r103 38 39 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.77
+ $Y=0.198 $X2=0.774 $Y2=0.198
r104 37 38 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.767
+ $Y=0.198 $X2=0.77 $Y2=0.198
r105 36 37 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.198 $X2=0.767 $Y2=0.198
r106 35 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.801 $Y=0.198 $X2=0.81 $Y2=0.207
r107 35 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.801
+ $Y=0.198 $X2=0.792 $Y2=0.198
r108 33 34 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.167 $X2=0.747 $Y2=0.178
r109 32 33 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.164 $X2=0.747 $Y2=0.167
r110 31 32 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.121 $X2=0.747 $Y2=0.164
r111 26 31 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.09 $X2=0.747 $Y2=0.121
r112 24 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.747 $Y=0.189 $X2=0.756 $Y2=0.198
r113 24 34 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.189 $X2=0.747 $Y2=0.178
r114 23 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.216 $X2=0.81
+ $Y2=0.216
r115 20 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2025 $X2=0.81 $Y2=0.2025
r116 19 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.2025 $X2=0.81 $Y2=0.2025
r117 17 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.747 $Y=0.09 $X2=0.747
+ $Y2=0.09
r118 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.758 $Y2=0.0675
r119 12 17 12.0194 $w=8.1e-08 $l=4.7e-08 $layer=LISD $thickness=2.8e-08 $X=0.7
+ $Y=0.0675 $X2=0.747 $Y2=0.0675
r120 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.0675 $X2=0.7 $Y2=0.0675
r121 5 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.945 $Y=0.135 $X2=0.945
+ $Y2=0.135
r122 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.945
+ $Y=0.135 $X2=0.945 $Y2=0.2025
r123 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.945
+ $Y=0.0675 $X2=0.945 $Y2=0.135
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%12 2 5 7 9 12 14 17 19 21 25 27 32 36 37 38 43 44
+ VSS
c31 44 VSS 2.89087e-19 $X=1.314 $Y=0.09
c32 43 VSS 1.16913e-19 $X=1.323 $Y=0.09
c33 38 VSS 1.92014e-19 $X=1.323 $Y=0.144
c34 37 VSS 2.83021e-19 $X=1.323 $Y=0.126
c35 36 VSS 4.65462e-19 $X=1.323 $Y=0.182
c36 34 VSS 1.81242e-20 $X=1.2915 $Y=0.191
c37 33 VSS 2.15286e-20 $X=1.287 $Y=0.191
c38 32 VSS 0.00127461f $X=1.283 $Y=0.191
c39 31 VSS 7.15474e-19 $X=1.242 $Y=0.191
c40 27 VSS 5.27395e-20 $X=1.224 $Y=0.191
c41 26 VSS 3.73006e-19 $X=1.314 $Y=0.191
c42 25 VSS 2.89178e-19 $X=1.215 $Y=0.163
c43 21 VSS 1.79849e-19 $X=1.215 $Y=0.135
c44 19 VSS 7.49026e-19 $X=1.215 $Y=0.182
c45 17 VSS 0.00885042f $X=1.294 $Y=0.2025
c46 12 VSS 0.0205477f $X=1.294 $Y=0.0675
c47 5 VSS 0.00122126f $X=1.215 $Y=0.135
c48 2 VSS 0.0583406f $X=1.215 $Y=0.0675
r49 44 45 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.314
+ $Y=0.09 $X2=1.3185 $Y2=0.09
r50 43 45 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.09 $X2=1.3185 $Y2=0.09
r51 40 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.09 $X2=1.314 $Y2=0.09
r52 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.126 $X2=1.323 $Y2=0.144
r53 36 38 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.182 $X2=1.323 $Y2=0.144
r54 35 43 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.099 $X2=1.323 $Y2=0.09
r55 35 37 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.099 $X2=1.323 $Y2=0.126
r56 33 34 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.287
+ $Y=0.191 $X2=1.2915 $Y2=0.191
r57 32 33 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=1.283
+ $Y=0.191 $X2=1.287 $Y2=0.191
r58 31 32 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.242
+ $Y=0.191 $X2=1.283 $Y2=0.191
r59 29 34 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.296
+ $Y=0.191 $X2=1.2915 $Y2=0.191
r60 27 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.224
+ $Y=0.191 $X2=1.242 $Y2=0.191
r61 26 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.314 $Y=0.191 $X2=1.323 $Y2=0.182
r62 26 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.314
+ $Y=0.191 $X2=1.296 $Y2=0.191
r63 24 25 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.144 $X2=1.215 $Y2=0.163
r64 21 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.135 $X2=1.215 $Y2=0.144
r65 19 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.215 $Y=0.182 $X2=1.224 $Y2=0.191
r66 19 25 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=1.215
+ $Y=0.182 $X2=1.215 $Y2=0.163
r67 17 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.191 $X2=1.296
+ $Y2=0.191
r68 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.279 $Y=0.2025 $X2=1.294 $Y2=0.2025
r69 12 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.09 $X2=1.296
+ $Y2=0.09
r70 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.279 $Y=0.0675 $X2=1.294 $Y2=0.0675
r71 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.215 $Y=0.135 $X2=1.215
+ $Y2=0.135
r72 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.215
+ $Y=0.135 $X2=1.215 $Y2=0.2025
r73 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.215
+ $Y=0.0675 $X2=1.215 $Y2=0.135
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%13 2 5 7 10 15 18 23 26 31 34 37 39 41 42 46 47 50
+ 51 53 59 60 61 62 63 66 67 72 73 74 77 80 81 82 83 86 87 90 91 92 94 105 107
+ 110 VSS
c67 110 VSS 2.79962e-19 $X=1.377 $Y=0.135
c68 108 VSS 4.98311e-20 $X=1.2645 $Y=0.135
c69 107 VSS 3.49116e-19 $X=1.26 $Y=0.135
c70 105 VSS 5.14517e-19 $X=1.269 $Y=0.135
c71 101 VSS 0.00253921f $X=1.251 $Y=0.036
c72 97 VSS 0.00331528f $X=1.431 $Y=0.135
c73 94 VSS 0.00474203f $X=1.377 $Y=0.225
c74 92 VSS 0.00144937f $X=1.377 $Y=0.1035
c75 91 VSS 0.00219086f $X=1.377 $Y=0.081
c76 90 VSS 0.00103511f $X=1.377 $Y=0.126
c77 88 VSS 0.00208651f $X=1.35 $Y=0.036
c78 87 VSS 0.00350381f $X=1.332 $Y=0.036
c79 86 VSS 3.87876e-19 $X=1.287 $Y=0.036
c80 85 VSS 0.00192765f $X=1.283 $Y=0.036
c81 83 VSS 0.00526264f $X=1.368 $Y=0.036
c82 82 VSS 4.91035e-19 $X=1.251 $Y=0.116
c83 81 VSS 2.41096e-19 $X=1.251 $Y=0.106
c84 80 VSS 7.80213e-19 $X=1.251 $Y=0.099
c85 79 VSS 4.80483e-19 $X=1.251 $Y=0.081
c86 78 VSS 4.9709e-19 $X=1.251 $Y=0.07
c87 77 VSS 0.00124273f $X=1.251 $Y=0.063
c88 76 VSS 1.26074e-19 $X=1.251 $Y=0.126
c89 74 VSS 0.00146362f $X=1.224 $Y=0.036
c90 73 VSS 0.00333697f $X=1.206 $Y=0.036
c91 72 VSS 0.00146362f $X=1.17 $Y=0.036
c92 71 VSS 0.00251494f $X=1.152 $Y=0.036
c93 67 VSS 0.0045992f $X=1.134 $Y=0.036
c94 66 VSS 0.00224226f $X=1.134 $Y=0.036
c95 64 VSS 0.00328022f $X=1.242 $Y=0.036
c96 63 VSS 0.0129562f $X=1.332 $Y=0.234
c97 62 VSS 0.00350786f $X=1.206 $Y=0.234
c98 61 VSS 0.00141253f $X=1.17 $Y=0.234
c99 60 VSS 0.00310297f $X=1.152 $Y=0.234
c100 59 VSS 0.00146362f $X=1.116 $Y=0.234
c101 58 VSS 0.00245593f $X=1.098 $Y=0.234
c102 53 VSS 0.00215392f $X=1.08 $Y=0.234
c103 51 VSS 0.00775972f $X=1.368 $Y=0.234
c104 50 VSS 0.00362692f $X=1.08 $Y=0.2025
c105 46 VSS 5.38922e-19 $X=1.097 $Y=0.2025
c106 41 VSS 5.38922e-19 $X=1.151 $Y=0.0675
c107 37 VSS 0.0148754f $X=1.593 $Y=0.135
c108 34 VSS 0.0645347f $X=1.593 $Y=0.0675
c109 26 VSS 0.0644226f $X=1.539 $Y=0.0675
c110 18 VSS 0.0644226f $X=1.485 $Y=0.0675
c111 10 VSS 0.0650932f $X=1.431 $Y=0.0675
c112 5 VSS 0.00193244f $X=1.269 $Y=0.135
c113 2 VSS 0.0615704f $X=1.269 $Y=0.0675
r114 107 108 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.26
+ $Y=0.135 $X2=1.2645 $Y2=0.135
r115 105 108 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.269 $Y=0.135 $X2=1.2645 $Y2=0.135
r116 102 107 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.135 $X2=1.26 $Y2=0.135
r117 95 110 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.386
+ $Y=0.135 $X2=1.377 $Y2=0.135
r118 95 97 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.386
+ $Y=0.135 $X2=1.431 $Y2=0.135
r119 93 110 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.144 $X2=1.377 $Y2=0.135
r120 93 94 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.144 $X2=1.377 $Y2=0.225
r121 91 92 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.081 $X2=1.377 $Y2=0.1035
r122 90 110 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.126 $X2=1.377 $Y2=0.135
r123 90 92 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.126 $X2=1.377 $Y2=0.1035
r124 89 91 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.045 $X2=1.377 $Y2=0.081
r125 87 88 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.332
+ $Y=0.036 $X2=1.35 $Y2=0.036
r126 86 87 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.287
+ $Y=0.036 $X2=1.332 $Y2=0.036
r127 85 86 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=1.283
+ $Y=0.036 $X2=1.287 $Y2=0.036
r128 84 101 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.26
+ $Y=0.036 $X2=1.251 $Y2=0.036
r129 84 85 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=1.26
+ $Y=0.036 $X2=1.283 $Y2=0.036
r130 83 89 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.368 $Y=0.036 $X2=1.377 $Y2=0.045
r131 83 88 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.368
+ $Y=0.036 $X2=1.35 $Y2=0.036
r132 81 82 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.106 $X2=1.251 $Y2=0.116
r133 80 81 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.099 $X2=1.251 $Y2=0.106
r134 79 80 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.081 $X2=1.251 $Y2=0.099
r135 78 79 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.07 $X2=1.251 $Y2=0.081
r136 77 78 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.063 $X2=1.251 $Y2=0.07
r137 76 102 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.126 $X2=1.251 $Y2=0.135
r138 76 82 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.126 $X2=1.251 $Y2=0.116
r139 75 101 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.045 $X2=1.251 $Y2=0.036
r140 75 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.251
+ $Y=0.045 $X2=1.251 $Y2=0.063
r141 73 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.206
+ $Y=0.036 $X2=1.224 $Y2=0.036
r142 72 73 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.17
+ $Y=0.036 $X2=1.206 $Y2=0.036
r143 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.152
+ $Y=0.036 $X2=1.17 $Y2=0.036
r144 66 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.134
+ $Y=0.036 $X2=1.152 $Y2=0.036
r145 66 67 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.134 $Y=0.036
+ $X2=1.134 $Y2=0.036
r146 64 101 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.242
+ $Y=0.036 $X2=1.251 $Y2=0.036
r147 64 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.242
+ $Y=0.036 $X2=1.224 $Y2=0.036
r148 62 63 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M1 $thickness=3.6e-08 $X=1.206
+ $Y=0.234 $X2=1.332 $Y2=0.234
r149 61 62 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.17
+ $Y=0.234 $X2=1.206 $Y2=0.234
r150 60 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.152
+ $Y=0.234 $X2=1.17 $Y2=0.234
r151 59 60 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.116
+ $Y=0.234 $X2=1.152 $Y2=0.234
r152 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.098
+ $Y=0.234 $X2=1.116 $Y2=0.234
r153 53 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.098 $Y2=0.234
r154 51 94 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.368 $Y=0.234 $X2=1.377 $Y2=0.225
r155 51 63 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.368
+ $Y=0.234 $X2=1.332 $Y2=0.234
r156 50 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234 $X2=1.08
+ $Y2=0.234
r157 47 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2025 $X2=1.08 $Y2=0.2025
r158 46 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.097 $Y=0.2025 $X2=1.08 $Y2=0.2025
r159 45 67 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=1.134 $Y=0.0675 $X2=1.134 $Y2=0.036
r160 42 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.117 $Y=0.0675 $X2=1.134 $Y2=0.0675
r161 41 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.151 $Y=0.0675 $X2=1.134 $Y2=0.0675
r162 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.593 $Y=0.135 $X2=1.593 $Y2=0.2025
r163 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.593 $Y=0.0675 $X2=1.593 $Y2=0.135
r164 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.539
+ $Y=0.135 $X2=1.593 $Y2=0.135
r165 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.539 $Y=0.135 $X2=1.539 $Y2=0.2025
r166 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.539 $Y=0.0675 $X2=1.539 $Y2=0.135
r167 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.485
+ $Y=0.135 $X2=1.539 $Y2=0.135
r168 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.485 $Y=0.135 $X2=1.485 $Y2=0.2025
r169 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.485 $Y=0.0675 $X2=1.485 $Y2=0.135
r170 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.431
+ $Y=0.135 $X2=1.485 $Y2=0.135
r171 13 97 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.431 $Y=0.135 $X2=1.431
+ $Y2=0.135
r172 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.431 $Y=0.135 $X2=1.431 $Y2=0.2025
r173 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.431 $Y=0.0675 $X2=1.431 $Y2=0.135
r174 5 105 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.269 $Y=0.135 $X2=1.269
+ $Y2=0.135
r175 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.269
+ $Y=0.135 $X2=1.269 $Y2=0.2025
r176 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.269
+ $Y=0.0675 $X2=1.269 $Y2=0.135
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%15 1 4 6 7 10 11 14 23 24 26 27 28 30 33 34 35 36
+ 37 VSS
c32 37 VSS 8.46035e-21 $X=0.63 $Y=0.198
c33 36 VSS 1.62375e-19 $X=0.612 $Y=0.198
c34 35 VSS 9.14524e-20 $X=0.599 $Y=0.198
c35 34 VSS 3.12342e-19 $X=0.58 $Y=0.198
c36 33 VSS 5.31938e-19 $X=0.576 $Y=0.198
c37 32 VSS 0.00134307f $X=0.558 $Y=0.198
c38 30 VSS 5.86427e-19 $X=0.648 $Y=0.198
c39 28 VSS 3.95078e-19 $X=0.531 $Y=0.198
c40 27 VSS 5.17397e-19 $X=0.522 $Y=0.198
c41 26 VSS 0.00400558f $X=0.504 $Y=0.198
c42 25 VSS 4.26131e-19 $X=0.468 $Y=0.198
c43 24 VSS 1.4604e-19 $X=0.459 $Y=0.198
c44 23 VSS 5.61374e-19 $X=0.45 $Y=0.198
c45 14 VSS 0.00375596f $X=0.646 $Y=0.2025
c46 10 VSS 0.00555436f $X=0.54 $Y=0.2025
c47 6 VSS 6.69874e-19 $X=0.557 $Y=0.2025
c48 4 VSS 0.00689207f $X=0.434 $Y=0.2025
c49 1 VSS 2.69461e-19 $X=0.449 $Y=0.2025
r50 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.198 $X2=0.63 $Y2=0.198
r51 35 36 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.599
+ $Y=0.198 $X2=0.612 $Y2=0.198
r52 34 35 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.58
+ $Y=0.198 $X2=0.599 $Y2=0.198
r53 33 34 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.198 $X2=0.58 $Y2=0.198
r54 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.198 $X2=0.576 $Y2=0.198
r55 30 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.198 $X2=0.63 $Y2=0.198
r56 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.198 $X2=0.531 $Y2=0.198
r57 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.198 $X2=0.522 $Y2=0.198
r58 25 26 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.198 $X2=0.504 $Y2=0.198
r59 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.198 $X2=0.468 $Y2=0.198
r60 23 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.198 $X2=0.459 $Y2=0.198
r61 21 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.198 $X2=0.558 $Y2=0.198
r62 21 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.198 $X2=0.531 $Y2=0.198
r63 17 23 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.45 $Y2=0.198
r64 14 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.198 $X2=0.648
+ $Y2=0.198
r65 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.646 $Y2=0.2025
r66 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.198 $X2=0.54
+ $Y2=0.198
r67 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r68 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r69 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r70 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.449
+ $Y=0.2025 $X2=0.434 $Y2=0.2025
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%16 1 2 5 6 9 16 18 19 20 21 23 VSS
c26 23 VSS 7.00634e-19 $X=0.747 $Y=0.234
c27 22 VSS 0.00298267f $X=0.738 $Y=0.234
c28 21 VSS 0.00103868f $X=0.711 $Y=0.234
c29 20 VSS 0.00157473f $X=0.702 $Y=0.234
c30 19 VSS 0.00206804f $X=0.684 $Y=0.234
c31 18 VSS 0.00706733f $X=0.662 $Y=0.234
c32 16 VSS 0.00225063f $X=0.756 $Y=0.234
c33 9 VSS 0.00345307f $X=0.758 $Y=0.2025
c34 6 VSS 7.37037e-19 $X=0.773 $Y=0.2025
c35 5 VSS 0.00358468f $X=0.594 $Y=0.2025
c36 1 VSS 6.32999e-19 $X=0.611 $Y=0.2025
r37 22 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.234 $X2=0.747 $Y2=0.234
r38 21 22 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.711
+ $Y=0.234 $X2=0.738 $Y2=0.234
r39 20 21 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.234 $X2=0.711 $Y2=0.234
r40 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.234 $X2=0.702 $Y2=0.234
r41 18 19 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.662
+ $Y=0.234 $X2=0.684 $Y2=0.234
r42 16 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.747 $Y2=0.234
r43 12 18 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.662 $Y2=0.234
r44 9 16 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234 $X2=0.756
+ $Y2=0.234
r45 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2025 $X2=0.758 $Y2=0.2025
r46 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r47 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.577
+ $Y=0.2025 $X2=0.594 $Y2=0.2025
r48 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.611
+ $Y=0.2025 $X2=0.594 $Y2=0.2025
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%QN 1 2 6 7 11 12 15 16 17 20 21 23 24 30 31 33 44
+ 45 VSS
c19 48 VSS 0.00300284f $X=1.6465 $Y=0.1845
c20 46 VSS 2.62283e-19 $X=1.6465 $Y=0.13025
c21 45 VSS 0.00548083f $X=1.6465 $Y=0.126
c22 44 VSS 6.00307e-19 $X=1.646 $Y=0.1345
c23 42 VSS 0.00247012f $X=1.6465 $Y=0.225
c24 33 VSS 0.00155282f $X=1.458 $Y=0.234
c25 31 VSS 0.0249971f $X=1.637 $Y=0.234
c26 30 VSS 0.00929647f $X=1.566 $Y=0.036
c27 24 VSS 0.00904424f $X=1.458 $Y=0.036
c28 23 VSS 0.00155282f $X=1.458 $Y=0.036
c29 21 VSS 0.0249971f $X=1.637 $Y=0.036
c30 20 VSS 0.00929647f $X=1.566 $Y=0.2025
c31 16 VSS 5.38922e-19 $X=1.583 $Y=0.2025
c32 15 VSS 0.00918054f $X=1.458 $Y=0.2025
c33 11 VSS 5.72268e-19 $X=1.475 $Y=0.2025
c34 6 VSS 5.38922e-19 $X=1.583 $Y=0.0675
c35 1 VSS 5.72268e-19 $X=1.475 $Y=0.0675
r36 47 48 2.57237 $w=1.9e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.144 $X2=1.6465 $Y2=0.1845
r37 45 46 0.26994 $w=1.9e-08 $l=4.25e-09 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.126 $X2=1.6465 $Y2=0.13025
r38 44 47 0.603395 $w=1.9e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.1345 $X2=1.6465 $Y2=0.144
r39 44 46 0.26994 $w=1.9e-08 $l=4.25e-09 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.1345 $X2=1.6465 $Y2=0.13025
r40 42 48 2.57237 $w=1.9e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.225 $X2=1.6465 $Y2=0.1845
r41 41 45 5.14474 $w=1.9e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.6465
+ $Y=0.045 $X2=1.6465 $Y2=0.126
r42 33 39 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.458
+ $Y=0.234 $X2=1.566 $Y2=0.234
r43 31 42 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.637 $Y=0.234 $X2=1.6465 $Y2=0.225
r44 31 39 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.637
+ $Y=0.234 $X2=1.566 $Y2=0.234
r45 29 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.566 $Y=0.036 $X2=1.566
+ $Y2=0.036
r46 23 29 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.458
+ $Y=0.036 $X2=1.566 $Y2=0.036
r47 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.458 $Y=0.036 $X2=1.458
+ $Y2=0.036
r48 21 41 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.637 $Y=0.036 $X2=1.6465 $Y2=0.045
r49 21 29 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.637
+ $Y=0.036 $X2=1.566 $Y2=0.036
r50 20 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.566 $Y=0.234 $X2=1.566
+ $Y2=0.234
r51 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.549 $Y=0.2025 $X2=1.566 $Y2=0.2025
r52 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.583 $Y=0.2025 $X2=1.566 $Y2=0.2025
r53 15 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.458 $Y=0.234 $X2=1.458
+ $Y2=0.234
r54 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.441 $Y=0.2025 $X2=1.458 $Y2=0.2025
r55 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.475 $Y=0.2025 $X2=1.458 $Y2=0.2025
r56 10 30 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.566
+ $Y=0.0675 $X2=1.566 $Y2=0.036
r57 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.549 $Y=0.0675 $X2=1.566 $Y2=0.0675
r58 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.583 $Y=0.0675 $X2=1.566 $Y2=0.0675
r59 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.458
+ $Y=0.0675 $X2=1.458 $Y2=0.036
r60 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.441
+ $Y=0.0675 $X2=1.458 $Y2=0.0675
r61 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=1.475
+ $Y=0.0675 $X2=1.458 $Y2=0.0675
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%18 1 6 9 VSS
c11 9 VSS 0.0194001f $X=0.866 $Y=0.0675
c12 6 VSS 3.25039e-19 $X=0.881 $Y=0.0675
c13 4 VSS 3.25039e-19 $X=0.808 $Y=0.0675
r14 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.881
+ $Y=0.0675 $X2=0.866 $Y2=0.0675
r15 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.808
+ $Y=0.0675 $X2=0.866 $Y2=0.0675
r16 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.793
+ $Y=0.0675 $X2=0.808 $Y2=0.0675
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%19 1 2 5 VSS
c5 5 VSS 0.00655974f $X=0.864 $Y=0.2025
c6 1 VSS 6.96227e-19 $X=0.881 $Y=0.2025
r7 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.847
+ $Y=0.2025 $X2=0.864 $Y2=0.2025
r8 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.881
+ $Y=0.2025 $X2=0.864 $Y2=0.2025
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%20 1 6 9 VSS
c13 9 VSS 0.0132338f $X=1.19 $Y=0.2025
c14 6 VSS 3.22787e-19 $X=1.205 $Y=0.2025
c15 4 VSS 3.14547e-19 $X=1.132 $Y=0.2025
r16 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=1.205
+ $Y=0.2025 $X2=1.19 $Y2=0.2025
r17 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=1.132
+ $Y=0.2025 $X2=1.19 $Y2=0.2025
r18 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=1.117
+ $Y=0.2025 $X2=1.132 $Y2=0.2025
.ends

.subckt PM_SDFLX4_ASAP7_75T_SRAM%23 1 2 VSS
c1 1 VSS 0.00183233f $X=1.205 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=1.205
+ $Y=0.0675 $X2=1.171 $Y2=0.0675
.ends


* END of "./SDFLx4_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt SDFLx4_ASAP7_75t_SRAM  VSS VDD CLK SE D SI QN
* 
* QN	QN
* SI	SI
* D	D
* SE	SE
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_9_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_7_M2_d N_SE_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 noxref_21 N_D_M3_g noxref_14 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M4 VSS N_7_M4_g noxref_21 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M5 noxref_22 N_SE_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M6 noxref_14 N_SI_M6_g noxref_22 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M7 N_11_M7_d N_9_M7_g noxref_14 VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M8 N_18_M8_d N_4_M8_g N_11_M8_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.027
M9 VSS N_10_M9_g N_18_M9_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.027
M10 N_10_M10_d N_11_M10_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.027
M11 N_13_M11_d N_4_M11_g N_10_M11_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=1.097 $Y=0.027
M12 N_23_M12_d N_9_M12_g N_13_M12_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=1.151 $Y=0.027
M13 VSS N_12_M13_g N_23_M13_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.027
M14 N_12_M14_d N_13_M14_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M15 N_QN_M15_d N_13_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.421
+ $Y=0.027
M16 N_QN_M16_d N_13_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.475
+ $Y=0.027
M17 N_QN_M17_d N_13_M17_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.529
+ $Y=0.027
M18 N_QN_M18_d N_13_M18_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.583
+ $Y=0.027
M19 VDD N_CLK_M19_g N_4_M19_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M20 N_9_M20_d N_4_M20_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M21 N_7_M21_d N_SE_M21_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M22 VDD N_D_M22_g N_15_M22_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M23 N_15_M23_d N_7_M23_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M24 N_16_M24_d N_SE_M24_g N_15_M24_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.557 $Y=0.162
M25 N_15_M25_d N_SI_M25_g N_16_M25_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.611 $Y=0.162
M26 N_11_M26_d N_4_M26_g N_16_M26_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.773 $Y=0.162
M27 N_19_M27_d N_9_M27_g N_11_M27_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.827 $Y=0.162
M28 VDD N_10_M28_g N_19_M28_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.162
M29 N_10_M29_d N_11_M29_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.162
M30 N_13_M30_d N_9_M30_g N_10_M30_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=1.043 $Y=0.162
M31 N_20_M31_d N_4_M31_g N_13_M31_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=1.097 $Y=0.162
M32 VDD N_12_M32_g N_20_M32_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.162
M33 N_12_M33_d N_13_M33_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
M34 N_QN_M34_d N_13_M34_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.421
+ $Y=0.162
M35 N_QN_M35_d N_13_M35_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.475
+ $Y=0.162
M36 N_QN_M36_d N_13_M36_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.529
+ $Y=0.162
M37 N_QN_M37_d N_13_M37_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.583
+ $Y=0.162
*
* 
* .include "SDFLx4_ASAP7_75t_SRAM.pex.sp.SDFLX4_ASAP7_75T_SRAM.pxi"
* BEGIN of "./SDFLx4_ASAP7_75t_SRAM.pex.sp.SDFLX4_ASAP7_75T_SRAM.pxi"
* File: SDFLx4_ASAP7_75t_SRAM.pex.sp.SDFLX4_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 13:05:41 2017
* 
x_PM_SDFLX4_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_2_p N_CLK_M19_g CLK VSS
+ PM_SDFLX4_ASAP7_75T_SRAM%CLK
x_PM_SDFLX4_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_15_n N_4_M20_g N_4_M8_g N_4_c_42_p
+ N_4_M26_g N_4_M11_g N_4_c_44_p N_4_M31_g N_4_M0_s N_4_M19_s N_4_c_16_n
+ N_4_c_17_n N_4_c_18_n N_4_c_19_n N_4_c_20_n N_4_c_22_n N_4_c_57_p N_4_c_23_n
+ N_4_c_24_n N_4_c_61_p N_4_c_25_n N_4_c_50_p N_4_c_27_p N_4_c_30_p N_4_c_39_p
+ N_4_c_63_p VSS PM_SDFLX4_ASAP7_75T_SRAM%4
x_PM_SDFLX4_ASAP7_75T_SRAM%SE N_SE_M2_g N_SE_c_98_n N_SE_M21_g N_SE_M5_g
+ N_SE_c_110_p N_SE_M24_g SE N_SE_c_114_p N_SE_c_100_n N_SE_c_101_n N_SE_c_102_n
+ N_SE_c_103_n N_SE_c_104_n N_SE_c_105_n VSS PM_SDFLX4_ASAP7_75T_SRAM%SE
x_PM_SDFLX4_ASAP7_75T_SRAM%D N_D_M3_g N_D_c_156_n N_D_M22_g D VSS
+ PM_SDFLX4_ASAP7_75T_SRAM%D
x_PM_SDFLX4_ASAP7_75T_SRAM%7 N_7_M4_g N_7_c_181_n N_7_M23_g N_7_M2_d N_7_M21_d
+ N_7_c_214_p N_7_c_182_n N_7_c_203_n N_7_c_183_n N_7_c_177_n N_7_c_184_n
+ N_7_c_185_n N_7_c_186_n N_7_c_188_n N_7_c_189_n N_7_c_190_n N_7_c_191_n
+ N_7_c_178_n N_7_c_193_n N_7_c_179_n N_7_c_196_n N_7_c_227_p N_7_c_197_n
+ N_7_c_212_n N_7_c_199_n N_7_c_200_n VSS PM_SDFLX4_ASAP7_75T_SRAM%7
x_PM_SDFLX4_ASAP7_75T_SRAM%SI N_SI_M6_g N_SI_c_234_n N_SI_M25_g SI VSS
+ PM_SDFLX4_ASAP7_75T_SRAM%SI
x_PM_SDFLX4_ASAP7_75T_SRAM%9 N_9_M7_g N_9_c_259_n N_9_M27_g N_9_c_261_n N_9_M30_g
+ N_9_M12_g N_9_c_264_n N_9_M1_d N_9_M20_d N_9_c_265_n N_9_c_268_n N_9_c_269_n
+ N_9_c_273_n N_9_c_294_n N_9_c_275_n N_9_c_277_n N_9_c_349_p N_9_c_278_n
+ N_9_c_357_p N_9_c_282_n N_9_c_283_n N_9_c_284_n N_9_c_286_n N_9_c_288_n
+ N_9_c_300_n N_9_c_257_n N_9_c_302_n N_9_c_290_n VSS PM_SDFLX4_ASAP7_75T_SRAM%9
x_PM_SDFLX4_ASAP7_75T_SRAM%10 N_10_M9_g N_10_c_390_n N_10_M28_g N_10_M10_d
+ N_10_M11_s N_10_c_382_n N_10_M29_d N_10_M30_s N_10_c_394_n N_10_c_384_n
+ N_10_c_385_n N_10_c_397_n N_10_c_386_n N_10_c_387_n N_10_c_401_p N_10_c_388_n
+ VSS PM_SDFLX4_ASAP7_75T_SRAM%10
x_PM_SDFLX4_ASAP7_75T_SRAM%11 N_11_M10_g N_11_c_431_n N_11_M29_g N_11_M7_d
+ N_11_M8_s N_11_c_418_n N_11_M27_s N_11_M26_d N_11_c_435_n N_11_c_463_p
+ N_11_c_420_n N_11_c_422_n N_11_c_438_n N_11_c_459_p N_11_c_439_n N_11_c_460_p
+ N_11_c_440_n N_11_c_468_p N_11_c_424_n N_11_c_441_n N_11_c_471_p N_11_c_442_n
+ N_11_c_444_n N_11_c_451_n N_11_c_426_n N_11_c_447_n VSS
+ PM_SDFLX4_ASAP7_75T_SRAM%11
x_PM_SDFLX4_ASAP7_75T_SRAM%12 N_12_M13_g N_12_c_479_n N_12_M32_g N_12_M14_d
+ N_12_c_489_p N_12_M33_d N_12_c_487_p N_12_c_480_n N_12_c_481_n N_12_c_482_n
+ N_12_c_488_p N_12_c_484_p N_12_c_502_p N_12_c_494_p N_12_c_503_p N_12_c_501_p
+ N_12_c_493_p VSS PM_SDFLX4_ASAP7_75T_SRAM%12
x_PM_SDFLX4_ASAP7_75T_SRAM%13 N_13_M14_g N_13_c_528_n N_13_M33_g N_13_M15_g
+ N_13_M34_g N_13_M16_g N_13_M35_g N_13_M17_g N_13_M36_g N_13_M18_g N_13_c_549_p
+ N_13_M37_g N_13_M12_s N_13_M11_d N_13_M31_s N_13_M30_d N_13_c_512_n
+ N_13_c_566_p N_13_c_514_n N_13_c_508_n N_13_c_516_n N_13_c_517_n N_13_c_571_p
+ N_13_c_529_n N_13_c_524_n N_13_c_510_n N_13_c_519_n N_13_c_573_p N_13_c_533_n
+ N_13_c_535_n N_13_c_536_n N_13_c_537_n N_13_c_538_n N_13_c_559_p N_13_c_539_n
+ N_13_c_540_n N_13_c_542_n N_13_c_543_n N_13_c_544_n N_13_c_545_n N_13_c_546_n
+ N_13_c_547_n N_13_c_548_n VSS PM_SDFLX4_ASAP7_75T_SRAM%13
x_PM_SDFLX4_ASAP7_75T_SRAM%15 N_15_M22_s N_15_c_578_n N_15_M24_s N_15_M23_d
+ N_15_c_588_n N_15_M25_d N_15_c_589_n N_15_c_579_n N_15_c_580_n N_15_c_591_n
+ N_15_c_582_n N_15_c_592_n N_15_c_584_n N_15_c_575_n N_15_c_594_n N_15_c_601_p
+ N_15_c_602_p N_15_c_585_n VSS PM_SDFLX4_ASAP7_75T_SRAM%15
x_PM_SDFLX4_ASAP7_75T_SRAM%16 N_16_M25_s N_16_M24_d N_16_c_608_n N_16_M26_s
+ N_16_c_613_n N_16_c_621_n N_16_c_607_n N_16_c_609_n N_16_c_611_n N_16_c_612_n
+ N_16_c_624_n VSS PM_SDFLX4_ASAP7_75T_SRAM%16
x_PM_SDFLX4_ASAP7_75T_SRAM%QN N_QN_M16_d N_QN_M15_d N_QN_M18_d N_QN_M17_d
+ N_QN_M35_d N_QN_M34_d N_QN_c_636_n N_QN_M37_d N_QN_M36_d N_QN_c_638_n
+ N_QN_c_639_n N_QN_c_642_n N_QN_c_644_n N_QN_c_645_n N_QN_c_646_n N_QN_c_649_n
+ QN N_QN_c_651_n VSS PM_SDFLX4_ASAP7_75T_SRAM%QN
x_PM_SDFLX4_ASAP7_75T_SRAM%18 N_18_M8_d N_18_M9_s N_18_c_652_n VSS
+ PM_SDFLX4_ASAP7_75T_SRAM%18
x_PM_SDFLX4_ASAP7_75T_SRAM%19 N_19_M28_s N_19_M27_d N_19_c_663_n VSS
+ PM_SDFLX4_ASAP7_75T_SRAM%19
x_PM_SDFLX4_ASAP7_75T_SRAM%20 N_20_M31_d N_20_M32_s N_20_c_668_n VSS
+ PM_SDFLX4_ASAP7_75T_SRAM%20
x_PM_SDFLX4_ASAP7_75T_SRAM%23 N_23_M13_s N_23_M12_d VSS PM_SDFLX4_ASAP7_75T_SRAM%23
cc_1 N_CLK_M0_g N_4_M1_g 0.00287079f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_CLK_c_2_p N_4_c_15_n 0.00101351f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 CLK N_4_c_16_n 0.00121601f $X=0.081 $Y=0.1345 $X2=0.056 $Y2=0.2025
cc_4 CLK N_4_c_17_n 5.67914e-19 $X=0.081 $Y=0.1345 $X2=0.018 $Y2=0.108
cc_5 CLK N_4_c_18_n 5.67914e-19 $X=0.081 $Y=0.1345 $X2=0.018 $Y2=0.0855
cc_6 CLK N_4_c_19_n 0.00221557f $X=0.081 $Y=0.1345 $X2=0.018 $Y2=0.2
cc_7 N_CLK_M0_g N_4_c_20_n 2.42151e-19 $X=0.081 $Y=0.0675 $X2=0.054 $Y2=0.036
cc_8 CLK N_4_c_20_n 0.00198278f $X=0.081 $Y=0.1345 $X2=0.054 $Y2=0.036
cc_9 CLK N_4_c_22_n 9.57337e-19 $X=0.081 $Y=0.1345 $X2=0.054 $Y2=0.036
cc_10 CLK N_4_c_23_n 0.00121787f $X=0.081 $Y=0.1345 $X2=0.033 $Y2=0.117
cc_11 CLK N_4_c_24_n 0.00368715f $X=0.081 $Y=0.1345 $X2=0.135 $Y2=0.117
cc_12 CLK N_4_c_25_n 8.02183e-19 $X=0.081 $Y=0.1345 $X2=0.175 $Y2=0.117
cc_13 CLK N_9_c_257_n 2.03179e-19 $X=0.081 $Y=0.1345 $X2=0 $Y2=0
cc_14 N_4_c_15_n N_SE_c_98_n 2.02054e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_15 N_4_c_27_p N_SE_c_98_n 2.65253e-19 $X=0.581 $Y=0.117 $X2=0.081 $Y2=0.135
cc_16 N_4_c_27_p N_SE_c_100_n 0.00116615f $X=0.581 $Y=0.117 $X2=0 $Y2=0
cc_17 N_4_c_27_p N_SE_c_101_n 0.0291792f $X=0.581 $Y=0.117 $X2=0 $Y2=0
cc_18 N_4_c_30_p N_SE_c_102_n 3.49768e-19 $X=0.682 $Y=0.117 $X2=0 $Y2=0
cc_19 N_4_c_27_p N_SE_c_103_n 3.29785e-19 $X=0.581 $Y=0.117 $X2=0 $Y2=0
cc_20 N_4_c_27_p N_SE_c_104_n 2.46239e-19 $X=0.581 $Y=0.117 $X2=0 $Y2=0
cc_21 N_4_c_27_p N_SE_c_105_n 5.96604e-19 $X=0.581 $Y=0.117 $X2=0 $Y2=0
cc_22 N_4_c_27_p D 0.0013631f $X=0.581 $Y=0.117 $X2=0 $Y2=0
cc_23 N_4_c_27_p N_7_c_177_n 0.0010068f $X=0.581 $Y=0.117 $X2=0 $Y2=0
cc_24 N_4_c_27_p N_7_c_178_n 4.55831e-19 $X=0.581 $Y=0.117 $X2=0 $Y2=0
cc_25 N_4_c_27_p N_7_c_179_n 4.65024e-19 $X=0.581 $Y=0.117 $X2=0 $Y2=0
cc_26 N_4_c_30_p SI 0.00138281f $X=0.682 $Y=0.117 $X2=0.081 $Y2=0.1345
cc_27 N_4_c_39_p SI 6.61251e-19 $X=1.107 $Y=0.117 $X2=0.081 $Y2=0.1345
cc_28 N_4_M8_g N_9_M7_g 2.94371e-19 $X=0.783 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_29 N_4_M8_g N_9_c_259_n 0.00355599f $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_4_c_42_p N_9_c_259_n 0.00105615f $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_31 N_4_M11_g N_9_c_261_n 0.00365763f $X=1.107 $Y=0.0675 $X2=0 $Y2=0
cc_32 N_4_c_44_p N_9_c_261_n 0.00104184f $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_33 N_4_M11_g N_9_M12_g 0.00355599f $X=1.107 $Y=0.0675 $X2=0 $Y2=0
cc_34 N_4_c_44_p N_9_c_264_n 9.99654e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_35 N_4_c_16_n N_9_c_265_n 2.58009e-19 $X=0.056 $Y=0.2025 $X2=0 $Y2=0
cc_36 N_4_c_24_n N_9_c_265_n 0.00114532f $X=0.135 $Y=0.117 $X2=0 $Y2=0
cc_37 N_4_c_25_n N_9_c_265_n 2.54113e-19 $X=0.175 $Y=0.117 $X2=0 $Y2=0
cc_38 N_4_c_50_p N_9_c_268_n 2.25982e-19 $X=0.229 $Y=0.117 $X2=0 $Y2=0
cc_39 N_4_M1_g N_9_c_269_n 3.53841e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_40 N_4_c_20_n N_9_c_269_n 6.34683e-19 $X=0.054 $Y=0.036 $X2=0 $Y2=0
cc_41 N_4_c_24_n N_9_c_269_n 5.44188e-19 $X=0.135 $Y=0.117 $X2=0 $Y2=0
cc_42 N_4_c_25_n N_9_c_269_n 2.25982e-19 $X=0.175 $Y=0.117 $X2=0 $Y2=0
cc_43 N_4_c_22_n N_9_c_273_n 2.56213e-19 $X=0.054 $Y=0.036 $X2=0 $Y2=0
cc_44 N_4_c_25_n N_9_c_273_n 3.0124e-19 $X=0.175 $Y=0.117 $X2=0 $Y2=0
cc_45 N_4_c_57_p N_9_c_275_n 2.66501e-19 $X=0.054 $Y=0.234 $X2=0 $Y2=0
cc_46 N_4_c_25_n N_9_c_275_n 3.28854e-19 $X=0.175 $Y=0.117 $X2=0 $Y2=0
cc_47 N_4_c_50_p N_9_c_277_n 2.46239e-19 $X=0.229 $Y=0.117 $X2=0 $Y2=0
cc_48 N_4_c_24_n N_9_c_278_n 3.53853e-19 $X=0.135 $Y=0.117 $X2=0 $Y2=0
cc_49 N_4_c_61_p N_9_c_278_n 9.64586e-19 $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_50 N_4_c_50_p N_9_c_278_n 0.0783963f $X=0.229 $Y=0.117 $X2=0 $Y2=0
cc_51 N_4_c_63_p N_9_c_278_n 0.00107275f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_52 N_4_c_42_p N_9_c_282_n 4.70423e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_53 N_4_c_39_p N_9_c_283_n 2.46239e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_54 N_4_c_61_p N_9_c_284_n 0.00403694f $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_55 N_4_c_39_p N_9_c_284_n 0.00115955f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_56 N_4_c_39_p N_9_c_286_n 0.00124223f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_57 N_4_c_63_p N_9_c_286_n 0.00262191f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_58 N_4_c_39_p N_9_c_288_n 3.53977e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_59 N_4_c_63_p N_9_c_288_n 0.00260528f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_60 N_4_c_24_n N_9_c_290_n 0.0038017f $X=0.135 $Y=0.117 $X2=0 $Y2=0
cc_61 N_4_c_50_p N_9_c_290_n 9.1421e-19 $X=0.229 $Y=0.117 $X2=0 $Y2=0
cc_62 N_4_M8_g N_10_M9_g 2.82885e-19 $X=0.783 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_63 N_4_c_39_p N_10_c_382_n 0.00134228f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_64 N_4_c_63_p N_10_c_382_n 0.00127195f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_65 N_4_c_39_p N_10_c_384_n 3.31762e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_66 N_4_c_39_p N_10_c_385_n 5.67404e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_67 N_4_c_39_p N_10_c_386_n 3.4734e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_68 N_4_c_39_p N_10_c_387_n 4.8206e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_69 N_4_c_39_p N_10_c_388_n 4.09721e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_70 N_4_c_61_p N_11_c_418_n 4.91424e-19 $X=0.783 $Y=0.117 $X2=0.081 $Y2=0.135
cc_71 N_4_c_39_p N_11_c_418_n 8.86983e-19 $X=1.107 $Y=0.117 $X2=0.081 $Y2=0.135
cc_72 N_4_c_61_p N_11_c_420_n 0.00811029f $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_73 N_4_c_39_p N_11_c_420_n 5.82789e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_74 N_4_c_61_p N_11_c_422_n 2.60223e-19 $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_75 N_4_c_39_p N_11_c_422_n 3.09845e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_76 N_4_M8_g N_11_c_424_n 3.61002e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_77 N_4_c_61_p N_11_c_424_n 0.001177f $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_78 N_4_c_39_p N_11_c_426_n 9.67845e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_79 N_4_M11_g N_12_M13_g 2.82885e-19 $X=1.107 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_80 N_4_M11_g N_13_c_508_n 3.47081e-19 $X=1.107 $Y=0.0675 $X2=0 $Y2=0
cc_81 N_4_c_63_p N_13_c_508_n 4.94366e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_82 N_4_c_63_p N_13_c_510_n 0.00130997f $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_83 VSS N_4_c_30_p 2.05877e-19 $X=0.682 $Y=0.117 $X2=0 $Y2=0
cc_84 N_4_c_61_p N_18_c_652_n 0.00102036f $X=0.783 $Y=0.117 $X2=0 $Y2=0
cc_85 N_4_c_39_p N_18_c_652_n 9.9685e-19 $X=1.107 $Y=0.117 $X2=0 $Y2=0
cc_86 N_SE_M5_g N_D_M3_g 2.13359e-19 $X=0.567 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_87 N_SE_c_98_n N_D_c_156_n 2.39808e-19 $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.135
cc_88 N_SE_c_101_n D 3.54801e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_89 N_SE_M5_g N_7_M4_g 0.00304756f $X=0.567 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_90 N_SE_c_110_p N_7_c_181_n 0.00105615f $X=0.567 $Y=0.135 $X2=0.135 $Y2=0.135
cc_91 N_SE_c_100_n N_7_c_182_n 6.84024e-19 $X=0.243 $Y=0.081 $X2=1.107 $Y2=0.135
cc_92 N_SE_c_101_n N_7_c_183_n 6.55402e-19 $X=0.567 $Y=0.081 $X2=1.107
+ $Y2=0.2025
cc_93 SE N_7_c_184_n 4.48296e-19 $X=0.278 $Y=0.1345 $X2=0.071 $Y2=0.0675
cc_94 N_SE_c_114_p N_7_c_185_n 6.16983e-19 $X=0.243 $Y=0.135 $X2=0.056
+ $Y2=0.0675
cc_95 N_SE_c_101_n N_7_c_186_n 9.88868e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_96 N_SE_c_102_n N_7_c_186_n 0.00105704f $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_97 N_SE_c_101_n N_7_c_188_n 4.38038e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_98 N_SE_c_101_n N_7_c_189_n 0.00100123f $X=0.567 $Y=0.081 $X2=0.071
+ $Y2=0.2025
cc_99 N_SE_c_101_n N_7_c_190_n 0.00123902f $X=0.567 $Y=0.081 $X2=0.056
+ $Y2=0.2025
cc_100 N_SE_c_101_n N_7_c_191_n 4.81197e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_101 N_SE_c_103_n N_7_c_178_n 0.00105704f $X=0.567 $Y=0.135 $X2=0.018
+ $Y2=0.045
cc_102 N_SE_c_101_n N_7_c_193_n 5.77999e-19 $X=0.567 $Y=0.081 $X2=0.018
+ $Y2=0.063
cc_103 N_SE_c_104_n N_7_c_193_n 0.00115045f $X=0.567 $Y=0.106 $X2=0.018
+ $Y2=0.063
cc_104 N_SE_c_105_n N_7_c_179_n 0.00105704f $X=0.567 $Y=0.1205 $X2=0.018
+ $Y2=0.0855
cc_105 N_SE_c_101_n N_7_c_196_n 3.53821e-19 $X=0.567 $Y=0.081 $X2=0.018
+ $Y2=0.2125
cc_106 N_SE_c_100_n N_7_c_197_n 6.58915e-19 $X=0.243 $Y=0.081 $X2=0.054
+ $Y2=0.036
cc_107 N_SE_c_101_n N_7_c_197_n 4.3742e-19 $X=0.567 $Y=0.081 $X2=0.054 $Y2=0.036
cc_108 N_SE_c_114_p N_7_c_199_n 6.58915e-19 $X=0.243 $Y=0.135 $X2=0.054
+ $Y2=0.234
cc_109 N_SE_c_101_n N_7_c_200_n 3.89571e-19 $X=0.567 $Y=0.081 $X2=0.047
+ $Y2=0.234
cc_110 N_SE_M5_g N_SI_M6_g 0.00348334f $X=0.567 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_111 N_SE_c_110_p N_SI_c_234_n 0.00105615f $X=0.567 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_112 N_SE_c_102_n SI 7.03144e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_113 N_SE_c_103_n SI 0.00123983f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_114 N_SE_c_104_n SI 5.30073e-19 $X=0.567 $Y=0.106 $X2=0 $Y2=0
cc_115 N_SE_c_105_n SI 0.00123983f $X=0.567 $Y=0.1205 $X2=0 $Y2=0
cc_116 N_SE_M5_g N_9_M7_g 2.88628e-19 $X=0.567 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_117 N_SE_c_100_n N_9_c_268_n 0.00211947f $X=0.243 $Y=0.081 $X2=0.018
+ $Y2=0.045
cc_118 N_SE_c_114_p N_9_c_294_n 0.00211947f $X=0.243 $Y=0.135 $X2=0.047
+ $Y2=0.036
cc_119 N_SE_c_114_p N_9_c_277_n 0.00221288f $X=0.243 $Y=0.135 $X2=0.054
+ $Y2=0.234
cc_120 N_SE_c_98_n N_9_c_278_n 2.61615e-19 $X=0.297 $Y=0.135 $X2=0.783 $Y2=0.117
cc_121 N_SE_c_114_p N_9_c_278_n 8.88734e-19 $X=0.243 $Y=0.135 $X2=0.783
+ $Y2=0.117
cc_122 N_SE_c_101_n N_9_c_278_n 0.00161941f $X=0.567 $Y=0.081 $X2=0.783
+ $Y2=0.117
cc_123 N_SE_c_103_n N_9_c_278_n 8.13099e-19 $X=0.567 $Y=0.135 $X2=0.783
+ $Y2=0.117
cc_124 N_SE_c_100_n N_9_c_300_n 0.00211947f $X=0.243 $Y=0.081 $X2=0 $Y2=0
cc_125 N_SE_c_101_n N_9_c_257_n 3.51588e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_126 N_SE_c_114_p N_9_c_302_n 0.00211947f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_127 VSS N_SE_c_101_n 2.01433e-19 $X=0.567 $Y=0.081 $X2=0.783 $Y2=0.135
cc_128 VSS N_SE_c_101_n 4.83825e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_129 VSS N_SE_M5_g 2.34002e-19 $X=0.567 $Y=0.0675 $X2=1.107 $Y2=0.135
cc_130 VSS N_SE_c_102_n 0.00426739f $X=0.567 $Y=0.081 $X2=1.107 $Y2=0.135
cc_131 N_SE_M5_g N_15_c_575_n 3.61002e-19 $X=0.567 $Y=0.0675 $X2=0.056
+ $Y2=0.2025
cc_132 N_SE_c_103_n N_15_c_575_n 0.00117826f $X=0.567 $Y=0.135 $X2=0.056
+ $Y2=0.2025
cc_133 VSS N_SE_c_102_n 3.06453e-19 $X=0.567 $Y=0.081 $X2=0.135 $Y2=0.0675
cc_134 N_D_M3_g N_7_M4_g 0.00304756f $X=0.459 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_135 N_D_c_156_n N_7_c_181_n 0.00105595f $X=0.459 $Y=0.135 $X2=0.135 $Y2=0.135
cc_136 D N_7_c_203_n 0.00251305f $X=0.459 $Y=0.1345 $X2=1.107 $Y2=0.2025
cc_137 D N_7_c_177_n 0.00251305f $X=0.459 $Y=0.1345 $X2=0 $Y2=0
cc_138 D N_7_c_184_n 0.00251305f $X=0.459 $Y=0.1345 $X2=0.071 $Y2=0.0675
cc_139 D N_7_c_185_n 0.00251305f $X=0.459 $Y=0.1345 $X2=0.056 $Y2=0.0675
cc_140 D N_7_c_189_n 0.00388774f $X=0.459 $Y=0.1345 $X2=0.071 $Y2=0.2025
cc_141 N_D_M3_g N_7_c_190_n 2.16728e-19 $X=0.459 $Y=0.0675 $X2=0.056 $Y2=0.2025
cc_142 D N_7_c_190_n 0.00388774f $X=0.459 $Y=0.1345 $X2=0.056 $Y2=0.2025
cc_143 D N_7_c_178_n 0.00141867f $X=0.459 $Y=0.1345 $X2=0.018 $Y2=0.045
cc_144 D N_7_c_179_n 0.00141867f $X=0.459 $Y=0.1345 $X2=0.018 $Y2=0.0855
cc_145 D N_7_c_212_n 0.00251305f $X=0.459 $Y=0.1345 $X2=0.027 $Y2=0.234
cc_146 D N_9_c_278_n 0.00217382f $X=0.459 $Y=0.1345 $X2=0.783 $Y2=0.117
cc_147 VSS D 0.00172965f $X=0.459 $Y=0.1345 $X2=0.783 $Y2=0.135
cc_148 VSS N_D_M3_g 2.37298e-19 $X=0.459 $Y=0.0675 $X2=1.107 $Y2=0.0675
cc_149 D N_15_M22_s 3.13248e-19 $X=0.459 $Y=0.1345 $X2=0.135 $Y2=0.0675
cc_150 D N_15_c_578_n 0.00310236f $X=0.459 $Y=0.1345 $X2=0.135 $Y2=0.135
cc_151 D N_15_c_579_n 0.00415606f $X=0.459 $Y=0.1345 $X2=1.107 $Y2=0.2025
cc_152 D N_15_c_580_n 0.00115405f $X=0.459 $Y=0.1345 $X2=0 $Y2=0
cc_153 N_7_M4_g N_SI_M6_g 2.48122e-19 $X=0.513 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_154 N_7_c_214_p N_9_c_265_n 2.28803e-19 $X=0.322 $Y=0.2025 $X2=0.056
+ $Y2=0.2025
cc_155 N_7_c_214_p N_9_c_278_n 3.0124e-19 $X=0.322 $Y=0.2025 $X2=0.783 $Y2=0.117
cc_156 N_7_c_185_n N_9_c_278_n 9.75625e-19 $X=0.351 $Y=0.1845 $X2=0.783
+ $Y2=0.117
cc_157 N_7_c_178_n N_9_c_278_n 8.02031e-19 $X=0.513 $Y=0.135 $X2=0.783 $Y2=0.117
cc_158 N_7_c_199_n N_9_c_278_n 3.70293e-19 $X=0.342 $Y=0.234 $X2=0.783 $Y2=0.117
cc_159 VSS N_7_c_190_n 3.22316e-19 $X=0.468 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_160 VSS N_7_c_182_n 2.68628e-19 $X=0.351 $Y=0.063 $X2=0.783 $Y2=0.135
cc_161 VSS N_7_c_183_n 2.08206e-19 $X=0.351 $Y=0.099 $X2=0.783 $Y2=0.135
cc_162 VSS N_7_c_190_n 0.00291153f $X=0.468 $Y=0.072 $X2=0.783 $Y2=0.135
cc_163 VSS N_7_c_193_n 2.08206e-19 $X=0.513 $Y=0.099 $X2=0.783 $Y2=0.135
cc_164 VSS N_7_c_196_n 0.00133246f $X=0.324 $Y=0.036 $X2=0.783 $Y2=0.135
cc_165 VSS N_7_M4_g 2.34002e-19 $X=0.513 $Y=0.0675 $X2=1.107 $Y2=0.0675
cc_166 VSS N_7_c_190_n 0.00904478f $X=0.468 $Y=0.072 $X2=1.107 $Y2=0.0675
cc_167 VSS N_7_c_227_p 6.34674e-19 $X=0.351 $Y=0.036 $X2=1.107 $Y2=0.0675
cc_168 N_7_c_214_p N_15_c_578_n 0.00134514f $X=0.322 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_169 N_7_M4_g N_15_c_582_n 3.50974e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_170 N_7_c_178_n N_15_c_582_n 0.00116301f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_171 N_SI_M6_g N_9_M7_g 0.00360681f $X=0.621 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_172 SI N_9_M7_g 4.66746e-19 $X=0.621 $Y=0.1345 $X2=0.135 $Y2=0.0675
cc_173 SI N_9_c_278_n 8.81805e-19 $X=0.621 $Y=0.1345 $X2=0.783 $Y2=0.117
cc_174 N_SI_c_234_n N_9_c_282_n 0.00113912f $X=0.621 $Y=0.135 $X2=1.107
+ $Y2=0.117
cc_175 SI N_9_c_282_n 2.86943e-19 $X=0.621 $Y=0.1345 $X2=1.107 $Y2=0.117
cc_176 SI N_9_c_283_n 0.00176948f $X=0.621 $Y=0.1345 $X2=1.107 $Y2=0.117
cc_177 SI N_11_c_418_n 0.0083394f $X=0.621 $Y=0.1345 $X2=1.107 $Y2=0.0675
cc_178 SI N_11_c_420_n 0.00227527f $X=0.621 $Y=0.1345 $X2=0.056 $Y2=0.0675
cc_179 VSS SI 0.00196285f $X=0.621 $Y=0.1345 $X2=0 $Y2=0
cc_180 VSS SI 0.00389367f $X=0.621 $Y=0.1345 $X2=1.107 $Y2=0.0675
cc_181 VSS N_SI_M6_g 3.5204e-19 $X=0.621 $Y=0.0675 $X2=1.107 $Y2=0.2025
cc_182 VSS SI 6.77952e-19 $X=0.621 $Y=0.1345 $X2=1.107 $Y2=0.2025
cc_183 VSS SI 0.0010238f $X=0.621 $Y=0.1345 $X2=1.107 $Y2=0.2025
cc_184 SI N_15_c_584_n 4.77922e-19 $X=0.621 $Y=0.1345 $X2=0.071 $Y2=0.2025
cc_185 N_SI_M6_g N_15_c_585_n 2.75159e-19 $X=0.621 $Y=0.0675 $X2=0.018 $Y2=0.063
cc_186 SI N_15_c_585_n 0.00116629f $X=0.621 $Y=0.1345 $X2=0.018 $Y2=0.063
cc_187 N_SI_M6_g N_16_c_607_n 2.38237e-19 $X=0.621 $Y=0.0675 $X2=1.107
+ $Y2=0.0675
cc_188 N_9_c_259_n N_10_M9_g 0.00341068f $X=0.837 $Y=0.135 $X2=0.081 $Y2=0.135
cc_189 N_9_c_259_n N_10_c_390_n 0.00105614f $X=0.837 $Y=0.135 $X2=0.081
+ $Y2=0.2025
cc_190 N_9_c_261_n N_10_c_382_n 0.00639681f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_191 N_9_c_278_n N_10_c_382_n 2.84796e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_192 N_9_c_286_n N_10_c_382_n 0.00138138f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_193 N_9_c_278_n N_10_c_394_n 7.48953e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_194 N_9_c_286_n N_10_c_394_n 0.00132074f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_195 N_9_c_278_n N_10_c_384_n 8.26567e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_196 N_9_c_284_n N_10_c_397_n 0.0037946f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_197 N_9_c_278_n N_10_c_388_n 4.07109e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_198 N_9_c_286_n N_10_c_388_n 0.00113688f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_199 N_9_c_259_n N_11_M10_g 2.13359e-19 $X=0.837 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_200 N_9_c_261_n N_11_M10_g 2.82885e-19 $X=1.053 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_201 N_9_c_261_n N_11_c_431_n 5.25211e-19 $X=1.053 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_202 N_9_c_278_n N_11_c_418_n 3.09707e-19 $X=1.121 $Y=0.153 $X2=0.081
+ $Y2=0.135
cc_203 N_9_c_282_n N_11_c_418_n 0.0010746f $X=0.693 $Y=0.135 $X2=0.081 $Y2=0.135
cc_204 N_9_c_283_n N_11_c_418_n 3.92611e-19 $X=0.693 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_205 N_9_c_278_n N_11_c_435_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_206 N_9_c_278_n N_11_c_422_n 8.09198e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_207 N_9_c_283_n N_11_c_422_n 0.00106879f $X=0.693 $Y=0.135 $X2=0 $Y2=0
cc_208 N_9_c_283_n N_11_c_438_n 0.00106879f $X=0.693 $Y=0.135 $X2=0 $Y2=0
cc_209 N_9_c_278_n N_11_c_439_n 3.46508e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_210 N_9_c_278_n N_11_c_440_n 2.42614e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_211 N_9_c_278_n N_11_c_441_n 4.07711e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_212 N_9_c_259_n N_11_c_442_n 3.51501e-19 $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_213 N_9_c_284_n N_11_c_442_n 5.11397e-19 $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_214 N_9_c_278_n N_11_c_444_n 5.75072e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_215 N_9_c_278_n N_11_c_426_n 0.00107683f $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_216 N_9_c_286_n N_11_c_426_n 4.32979e-19 $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_217 N_9_c_286_n N_11_c_447_n 4.15367e-19 $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_218 N_9_M12_g N_12_M13_g 0.00341068f $X=1.161 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_219 N_9_c_264_n N_12_c_479_n 9.22047e-19 $X=1.161 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_220 N_9_c_288_n N_12_c_480_n 0.00206054f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_221 N_9_c_288_n N_12_c_481_n 0.00206054f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_222 N_9_c_349_p N_12_c_482_n 3.53853e-19 $X=1.161 $Y=0.153 $X2=0 $Y2=0
cc_223 N_9_M12_g N_13_M14_g 2.13359e-19 $X=1.161 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_224 N_9_c_278_n N_13_c_512_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_225 N_9_c_286_n N_13_c_512_n 0.00130837f $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_226 N_9_c_261_n N_13_c_514_n 2.20599e-19 $X=1.053 $Y=0.135 $X2=0 $Y2=0
cc_227 N_9_c_278_n N_13_c_514_n 5.75548e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_228 N_9_c_278_n N_13_c_516_n 3.8246e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_229 N_9_c_288_n N_13_c_517_n 0.00102938f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_230 N_9_c_357_p N_13_c_510_n 2.51466e-19 $X=1.141 $Y=0.153 $X2=0 $Y2=0
cc_231 N_9_M12_g N_13_c_519_n 3.57114e-19 $X=1.161 $Y=0.0675 $X2=0 $Y2=0
cc_232 N_9_c_288_n N_13_c_519_n 5.22021e-19 $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_233 N_9_c_278_n N_15_c_578_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0.081 $Y2=0.135
cc_234 N_9_c_278_n N_15_c_588_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_235 N_9_c_278_n N_15_c_589_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_236 N_9_c_278_n N_15_c_579_n 3.10744e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_237 N_9_c_278_n N_15_c_591_n 4.72621e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_238 N_9_c_278_n N_15_c_592_n 4.8224e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_239 N_9_c_278_n N_15_c_584_n 3.65983e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_240 N_9_c_278_n N_15_c_594_n 4.66683e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_241 N_9_c_278_n N_16_c_608_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0.081 $Y2=0.135
cc_242 N_9_M7_g N_16_c_609_n 4.39425e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_243 N_9_c_278_n N_16_c_609_n 3.48349e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_244 N_9_c_283_n N_16_c_611_n 5.53288e-19 $X=0.693 $Y=0.135 $X2=0 $Y2=0
cc_245 N_9_c_278_n N_16_c_612_n 6.02073e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_246 N_9_c_259_n N_18_c_652_n 0.00639681f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_247 N_9_c_278_n N_18_c_652_n 2.4912e-19 $X=1.121 $Y=0.153 $X2=0 $Y2=0
cc_248 N_9_c_284_n N_18_c_652_n 0.00372445f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_249 N_9_c_278_n N_19_c_663_n 3.0124e-19 $X=1.121 $Y=0.153 $X2=0.081 $Y2=0.135
cc_250 N_9_M12_g N_20_c_668_n 0.00382563f $X=1.161 $Y=0.0675 $X2=0 $Y2=0
cc_251 N_9_c_264_n N_20_c_668_n 0.0019701f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_252 N_9_c_357_p N_20_c_668_n 4.50035e-19 $X=1.141 $Y=0.153 $X2=0 $Y2=0
cc_253 N_9_c_288_n N_20_c_668_n 0.00376163f $X=1.161 $Y=0.135 $X2=0 $Y2=0
cc_254 N_10_M9_g N_11_M10_g 0.00268443f $X=0.891 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_255 N_10_c_401_p N_11_M10_g 3.61002e-19 $X=0.954 $Y=0.072 $X2=0.135
+ $Y2=0.0675
cc_256 N_10_c_390_n N_11_c_431_n 0.00105598f $X=0.891 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_257 N_10_M9_g N_11_c_451_n 3.56998e-19 $X=0.891 $Y=0.0675 $X2=0 $Y2=0
cc_258 N_10_c_384_n N_11_c_451_n 4.80589e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_259 N_10_c_394_n N_11_c_426_n 0.00242354f $X=1.028 $Y=0.2025 $X2=0.054
+ $Y2=0.234
cc_260 N_10_c_385_n N_11_c_426_n 0.0021413f $X=0.891 $Y=0.1205 $X2=0.054
+ $Y2=0.234
cc_261 N_10_c_401_p N_11_c_426_n 0.00118287f $X=0.954 $Y=0.072 $X2=0.054
+ $Y2=0.234
cc_262 N_10_c_388_n N_11_c_426_n 0.00115834f $X=0.999 $Y=0.162 $X2=0.054
+ $Y2=0.234
cc_263 N_10_c_382_n N_13_c_512_n 0.00122411f $X=1.082 $Y=0.0675 $X2=0 $Y2=0
cc_264 N_10_c_394_n N_13_c_512_n 0.00270924f $X=1.028 $Y=0.2025 $X2=0 $Y2=0
cc_265 N_10_c_394_n N_13_c_514_n 5.74875e-19 $X=1.028 $Y=0.2025 $X2=0.054
+ $Y2=0.234
cc_266 N_10_c_382_n N_13_c_524_n 3.1278e-19 $X=1.082 $Y=0.0675 $X2=0.783
+ $Y2=0.117
cc_267 N_10_c_382_n N_13_c_510_n 0.00278091f $X=1.082 $Y=0.0675 $X2=0.783
+ $Y2=0.117
cc_268 N_10_c_382_n N_18_c_652_n 3.26365e-19 $X=1.082 $Y=0.0675 $X2=0.783
+ $Y2=0.0675
cc_269 N_10_c_397_n N_18_c_652_n 0.00127189f $X=0.9 $Y=0.072 $X2=0.783
+ $Y2=0.0675
cc_270 N_10_c_394_n N_19_c_663_n 2.12502e-19 $X=1.028 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_271 N_10_c_394_n N_20_c_668_n 3.11986e-19 $X=1.028 $Y=0.2025 $X2=0.783
+ $Y2=0.0675
cc_272 VSS N_11_c_418_n 2.62157e-19 $X=0.758 $Y=0.0675 $X2=0 $Y2=0
cc_273 VSS N_11_c_418_n 0.004062f $X=0.758 $Y=0.0675 $X2=1.107 $Y2=0.0675
cc_274 N_11_c_459_p N_15_c_589_n 2.93059e-19 $X=0.747 $Y=0.178 $X2=0.783
+ $Y2=0.2025
cc_275 N_11_c_460_p N_15_c_584_n 6.37567e-19 $X=0.756 $Y=0.198 $X2=0.071
+ $Y2=0.2025
cc_276 N_11_c_418_n N_16_c_613_n 0.00114234f $X=0.758 $Y=0.0675 $X2=0.783
+ $Y2=0.0675
cc_277 N_11_c_435_n N_16_c_613_n 0.00380633f $X=0.81 $Y=0.2025 $X2=0.783
+ $Y2=0.0675
cc_278 N_11_c_463_p N_16_c_613_n 3.87816e-19 $X=0.747 $Y=0.189 $X2=0.783
+ $Y2=0.0675
cc_279 N_11_c_422_n N_16_c_613_n 4.18661e-19 $X=0.747 $Y=0.164 $X2=0.783
+ $Y2=0.0675
cc_280 N_11_c_459_p N_16_c_613_n 4.06284e-19 $X=0.747 $Y=0.178 $X2=0.783
+ $Y2=0.0675
cc_281 N_11_c_460_p N_16_c_613_n 6.70593e-19 $X=0.756 $Y=0.198 $X2=0.783
+ $Y2=0.0675
cc_282 N_11_c_440_n N_16_c_613_n 7.05929e-19 $X=0.767 $Y=0.198 $X2=0.783
+ $Y2=0.0675
cc_283 N_11_c_468_p N_16_c_613_n 4.19603e-19 $X=0.77 $Y=0.198 $X2=0.783
+ $Y2=0.0675
cc_284 N_11_c_435_n N_16_c_621_n 2.42261e-19 $X=0.81 $Y=0.2025 $X2=0 $Y2=0
cc_285 N_11_c_440_n N_16_c_621_n 0.00137625f $X=0.767 $Y=0.198 $X2=0 $Y2=0
cc_286 N_11_c_471_p N_16_c_621_n 9.77254e-19 $X=0.819 $Y=0.234 $X2=0 $Y2=0
cc_287 N_11_c_460_p N_16_c_624_n 0.00137625f $X=0.756 $Y=0.198 $X2=1.107
+ $Y2=0.2025
cc_288 N_11_c_418_n N_18_c_652_n 0.00479956f $X=0.758 $Y=0.0675 $X2=0.783
+ $Y2=0.0675
cc_289 N_11_c_435_n N_18_c_652_n 0.00138279f $X=0.81 $Y=0.2025 $X2=0.783
+ $Y2=0.0675
cc_290 N_11_c_435_n N_19_c_663_n 0.00335562f $X=0.81 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_291 N_11_c_444_n N_19_c_663_n 0.00242949f $X=0.882 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_292 N_12_M13_g N_13_M14_g 0.00268443f $X=1.215 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_293 N_12_c_484_p N_13_M14_g 3.29607e-19 $X=1.283 $Y=0.191 $X2=0.135
+ $Y2=0.0675
cc_294 N_12_c_479_n N_13_c_528_n 0.00108446f $X=1.215 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_295 N_12_M13_g N_13_c_529_n 2.64276e-19 $X=1.215 $Y=0.0675 $X2=0.135
+ $Y2=0.117
cc_296 N_12_c_487_p N_13_c_529_n 0.00321328f $X=1.294 $Y=0.2025 $X2=0.135
+ $Y2=0.117
cc_297 N_12_c_488_p N_13_c_529_n 0.00838811f $X=1.224 $Y=0.191 $X2=0.135
+ $Y2=0.117
cc_298 N_12_c_489_p N_13_c_510_n 2.02397e-19 $X=1.294 $Y=0.0675 $X2=0.783
+ $Y2=0.117
cc_299 N_12_M13_g N_13_c_533_n 3.57119e-19 $X=1.215 $Y=0.0675 $X2=1.107
+ $Y2=0.117
cc_300 N_12_c_481_n N_13_c_533_n 5.37372e-19 $X=1.215 $Y=0.135 $X2=1.107
+ $Y2=0.117
cc_301 N_12_c_489_p N_13_c_535_n 0.00115323f $X=1.294 $Y=0.0675 $X2=0 $Y2=0
cc_302 N_12_c_493_p N_13_c_536_n 9.36593e-19 $X=1.314 $Y=0.09 $X2=0 $Y2=0
cc_303 N_12_c_494_p N_13_c_537_n 7.6566e-19 $X=1.323 $Y=0.126 $X2=0 $Y2=0
cc_304 N_12_c_481_n N_13_c_538_n 0.0030621f $X=1.215 $Y=0.135 $X2=0 $Y2=0
cc_305 N_12_c_489_p N_13_c_539_n 6.1907e-19 $X=1.294 $Y=0.0675 $X2=0 $Y2=0
cc_306 N_12_c_489_p N_13_c_540_n 0.003475f $X=1.294 $Y=0.0675 $X2=0 $Y2=0
cc_307 N_12_c_493_p N_13_c_540_n 0.00207793f $X=1.314 $Y=0.09 $X2=0 $Y2=0
cc_308 N_12_c_494_p N_13_c_542_n 0.00149664f $X=1.323 $Y=0.126 $X2=0 $Y2=0
cc_309 N_12_c_489_p N_13_c_543_n 3.63761e-19 $X=1.294 $Y=0.0675 $X2=0 $Y2=0
cc_310 N_12_c_501_p N_13_c_544_n 0.00149664f $X=1.323 $Y=0.09 $X2=0 $Y2=0
cc_311 N_12_c_502_p N_13_c_545_n 0.00149664f $X=1.323 $Y=0.182 $X2=0 $Y2=0
cc_312 N_12_c_503_p N_13_c_546_n 9.53904e-19 $X=1.323 $Y=0.144 $X2=0 $Y2=0
cc_313 N_12_c_484_p N_13_c_547_n 0.00190954f $X=1.283 $Y=0.191 $X2=0 $Y2=0
cc_314 N_12_c_503_p N_13_c_548_n 0.00149664f $X=1.323 $Y=0.144 $X2=0.018
+ $Y2=0.117
cc_315 N_12_c_487_p N_20_c_668_n 2.83378e-19 $X=1.294 $Y=0.2025 $X2=0.783
+ $Y2=0.0675
cc_316 N_12_c_482_n N_20_c_668_n 0.00102083f $X=1.215 $Y=0.163 $X2=0.783
+ $Y2=0.0675
cc_317 N_13_c_549_p N_QN_M16_d 3.8044e-19 $X=1.593 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_318 N_13_c_549_p N_QN_M18_d 3.80663e-19 $X=1.593 $Y=0.135 $X2=0.135
+ $Y2=0.2025
cc_319 N_13_c_549_p N_QN_M35_d 3.8044e-19 $X=1.593 $Y=0.135 $X2=0 $Y2=0
cc_320 N_13_c_549_p N_QN_c_636_n 7.78051e-19 $X=1.593 $Y=0.135 $X2=0.783
+ $Y2=0.2025
cc_321 N_13_c_549_p N_QN_M37_d 3.80663e-19 $X=1.593 $Y=0.135 $X2=0 $Y2=0
cc_322 N_13_c_549_p N_QN_c_638_n 8.00061e-19 $X=1.593 $Y=0.135 $X2=1.107
+ $Y2=0.135
cc_323 N_13_M16_g N_QN_c_639_n 4.59284e-19 $X=1.485 $Y=0.0675 $X2=1.107
+ $Y2=0.135
cc_324 N_13_M17_g N_QN_c_639_n 4.59284e-19 $X=1.539 $Y=0.0675 $X2=1.107
+ $Y2=0.135
cc_325 N_13_M18_g N_QN_c_639_n 4.59284e-19 $X=1.593 $Y=0.0675 $X2=1.107
+ $Y2=0.135
cc_326 N_13_c_549_p N_QN_c_642_n 0.00187443f $X=1.593 $Y=0.135 $X2=1.107
+ $Y2=0.2025
cc_327 N_13_c_559_p N_QN_c_642_n 4.23911e-19 $X=1.368 $Y=0.036 $X2=1.107
+ $Y2=0.2025
cc_328 N_13_c_549_p N_QN_c_644_n 7.78051e-19 $X=1.593 $Y=0.135 $X2=0 $Y2=0
cc_329 N_13_c_549_p N_QN_c_645_n 8.00061e-19 $X=1.593 $Y=0.135 $X2=0.071
+ $Y2=0.2025
cc_330 N_13_M16_g N_QN_c_646_n 4.59284e-19 $X=1.485 $Y=0.0675 $X2=0.056
+ $Y2=0.2025
cc_331 N_13_M17_g N_QN_c_646_n 4.59284e-19 $X=1.539 $Y=0.0675 $X2=0.056
+ $Y2=0.2025
cc_332 N_13_M18_g N_QN_c_646_n 4.59284e-19 $X=1.593 $Y=0.0675 $X2=0.056
+ $Y2=0.2025
cc_333 N_13_c_549_p N_QN_c_649_n 0.00187443f $X=1.593 $Y=0.135 $X2=0.056
+ $Y2=0.2025
cc_334 N_13_c_566_p N_QN_c_649_n 4.26942e-19 $X=1.368 $Y=0.234 $X2=0.056
+ $Y2=0.2025
cc_335 N_13_c_549_p N_QN_c_651_n 5.09179e-19 $X=1.593 $Y=0.135 $X2=0.054
+ $Y2=0.036
cc_336 N_13_c_512_n N_20_c_668_n 0.00412407f $X=1.08 $Y=0.2025 $X2=0.783
+ $Y2=0.0675
cc_337 N_13_c_516_n N_20_c_668_n 0.00284013f $X=1.152 $Y=0.234 $X2=0.783
+ $Y2=0.0675
cc_338 N_13_c_517_n N_20_c_668_n 0.00111255f $X=1.17 $Y=0.234 $X2=0.783
+ $Y2=0.0675
cc_339 N_13_c_571_p N_20_c_668_n 0.00302676f $X=1.206 $Y=0.234 $X2=0.783
+ $Y2=0.0675
cc_340 N_13_c_510_n N_20_c_668_n 0.00114658f $X=1.134 $Y=0.036 $X2=0.783
+ $Y2=0.0675
cc_341 N_13_c_573_p N_20_c_668_n 2.10553e-19 $X=1.206 $Y=0.036 $X2=0.783
+ $Y2=0.0675
cc_342 N_13_c_573_p N_23_M13_s 4.40115e-19 $X=1.206 $Y=0.036 $X2=0.135
+ $Y2=0.0675
cc_343 VSS N_15_c_578_n 0.00124679f $X=0.432 $Y=0.036 $X2=0.135 $Y2=0.135
cc_344 VSS N_15_c_589_n 0.0012783f $X=0.648 $Y=0.036 $X2=0.783 $Y2=0.2025
cc_345 VSS N_18_c_652_n 3.09059e-19 $X=0.648 $Y=0.036 $X2=0.783 $Y2=0.0675
cc_346 N_15_c_588_n N_16_c_608_n 0.00323532f $X=0.54 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_347 N_15_c_589_n N_16_c_608_n 0.00352176f $X=0.646 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_348 N_15_c_601_p N_16_c_608_n 0.00145268f $X=0.599 $Y=0.198 $X2=0.135
+ $Y2=0.135
cc_349 N_15_c_602_p N_16_c_608_n 8.58362e-19 $X=0.612 $Y=0.198 $X2=0.135
+ $Y2=0.135
cc_350 N_15_c_589_n N_16_c_613_n 0.00122215f $X=0.646 $Y=0.2025 $X2=0.783
+ $Y2=0.0675
cc_351 N_15_c_588_n N_16_c_607_n 5.00576e-19 $X=0.54 $Y=0.2025 $X2=1.107
+ $Y2=0.0675
cc_352 N_15_c_589_n N_16_c_607_n 0.0030897f $X=0.646 $Y=0.2025 $X2=1.107
+ $Y2=0.0675
cc_353 N_15_c_601_p N_16_c_607_n 0.00701208f $X=0.599 $Y=0.198 $X2=1.107
+ $Y2=0.0675
cc_354 N_18_c_652_n N_19_c_663_n 0.00138279f $X=0.866 $Y=0.0675 $X2=0.135
+ $Y2=0.135

* END of "./SDFLx4_ASAP7_75t_SRAM.pex.sp.SDFLX4_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: ASYNC_DFFHx1_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:17:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "ASYNC_DFFHx1_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./ASYNC_DFFHx1_ASAP7_75t_SRAM.pex.sp.pex"
* File: ASYNC_DFFHx1_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:17:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%CLK 2 5 7 12 16 VSS
c21 16 VSS 0.00662527f $X=0.081 $Y=0.135
c22 12 VSS 0.00676076f $X=0.082 $Y=0.119
c23 5 VSS 0.00165173f $X=0.081 $Y=0.135
c24 2 VSS 0.0629053f $X=0.081 $Y=0.054
r25 12 16 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.135
r26 5 16 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%4 2 7 10 13 16 19 22 25 27 29 32 34 40 41 42
+ 45 46 49 56 63 71 72 76 77 79 81 82 87 88 92 97 103 VSS
c85 133 VSS 1.06551e-19 $X=0.03 $Y=0.153
c86 132 VSS 6.89947e-19 $X=0.027 $Y=0.153
c87 103 VSS 9.20776e-19 $X=0.838 $Y=0.113
c88 97 VSS 5.70978e-19 $X=0.459 $Y=0.135
c89 92 VSS 0.00108052f $X=0.351 $Y=0.135
c90 88 VSS 0.0011617f $X=0.151 $Y=0.135
c91 87 VSS 0.00317449f $X=0.151 $Y=0.135
c92 82 VSS 7.14075e-19 $X=0.735 $Y=0.153
c93 81 VSS 0.00151903f $X=0.632 $Y=0.153
c94 79 VSS 0.0010088f $X=0.838 $Y=0.153
c95 77 VSS 3.20221e-19 $X=0.4115 $Y=0.153
c96 76 VSS 0.0031123f $X=0.364 $Y=0.153
c97 72 VSS 0.00253309f $X=0.263 $Y=0.153
c98 71 VSS 0.00604304f $X=0.175 $Y=0.153
c99 63 VSS 6.74716e-19 $X=0.033 $Y=0.153
c100 59 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c101 58 VSS 0.00180216f $X=0.047 $Y=0.234
c102 56 VSS 0.00250119f $X=0.054 $Y=0.234
c103 54 VSS 0.00305101f $X=0.027 $Y=0.234
c104 52 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c105 51 VSS 0.00199699f $X=0.047 $Y=0.036
c106 49 VSS 0.00250119f $X=0.054 $Y=0.036
c107 47 VSS 0.00305101f $X=0.027 $Y=0.036
c108 46 VSS 4.88707e-19 $X=0.018 $Y=0.2125
c109 45 VSS 0.00180363f $X=0.018 $Y=0.2
c110 44 VSS 4.69158e-19 $X=0.018 $Y=0.225
c111 42 VSS 0.00173342f $X=0.018 $Y=0.107
c112 41 VSS 9.57865e-19 $X=0.018 $Y=0.07
c113 40 VSS 0.00183429f $X=0.018 $Y=0.144
c114 37 VSS 0.00509483f $X=0.056 $Y=0.216
c115 34 VSS 2.98509e-19 $X=0.071 $Y=0.216
c116 32 VSS 0.00497933f $X=0.056 $Y=0.054
c117 29 VSS 2.98509e-19 $X=0.071 $Y=0.054
c118 25 VSS 0.00158412f $X=0.837 $Y=0.111
c119 22 VSS 0.0608155f $X=0.837 $Y=0.054
c120 16 VSS 0.0648216f $X=0.459 $Y=0.135
c121 13 VSS 0.00144498f $X=0.351 $Y=0.135
c122 10 VSS 0.0593284f $X=0.351 $Y=0.0675
c123 2 VSS 0.0616396f $X=0.135 $Y=0.054
r124 132 133 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r125 129 132 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r126 87 88 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.151 $Y=0.135 $X2=0.151
+ $Y2=0.135
r127 81 82 6.99383 $w=1.8e-08 $l=1.03e-07 $layer=M2 $thickness=3.6e-08 $X=0.632
+ $Y=0.153 $X2=0.735 $Y2=0.153
r128 80 103 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.838
+ $Y=0.153 $X2=0.838 $Y2=0.113
r129 79 82 6.99383 $w=1.8e-08 $l=1.03e-07 $layer=M2 $thickness=3.6e-08 $X=0.838
+ $Y=0.153 $X2=0.735 $Y2=0.153
r130 79 80 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.838 $Y=0.153 $X2=0.838
+ $Y2=0.153
r131 76 77 3.22531 $w=1.8e-08 $l=4.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.364
+ $Y=0.153 $X2=0.4115 $Y2=0.153
r132 74 81 11.7469 $w=1.8e-08 $l=1.73e-07 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.632 $Y2=0.153
r133 74 77 3.22531 $w=1.8e-08 $l=4.75e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.4115 $Y2=0.153
r134 74 97 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.459 $Y=0.153 $X2=0.459
+ $Y2=0.153
r135 71 72 5.97531 $w=1.8e-08 $l=8.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.175
+ $Y=0.153 $X2=0.263 $Y2=0.153
r136 69 76 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.153 $X2=0.364 $Y2=0.153
r137 69 72 5.97531 $w=1.8e-08 $l=8.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.153 $X2=0.263 $Y2=0.153
r138 69 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.153 $X2=0.351
+ $Y2=0.153
r139 66 71 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.151
+ $Y=0.153 $X2=0.175 $Y2=0.153
r140 66 88 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.151 $Y=0.153 $X2=0.151
+ $Y2=0.153
r141 63 133 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r142 62 66 8.01235 $w=1.8e-08 $l=1.18e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.151 $Y2=0.153
r143 62 63 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r144 58 59 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r145 56 59 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r146 54 58 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r147 51 52 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r148 49 52 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r149 47 51 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r150 45 46 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r151 44 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r152 44 46 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r153 43 129 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r154 43 45 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.2
r155 41 42 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.107
r156 40 129 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r157 40 42 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.107
r158 39 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r159 39 41 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r160 37 56 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r161 34 37 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r162 32 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r163 29 32 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r164 25 103 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.838 $Y=0.113
+ $X2=0.838 $Y2=0.113
r165 25 27 443.961 $w=2e-08 $l=1.185e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.111 $X2=0.837 $Y2=0.2295
r166 22 25 213.551 $w=2e-08 $l=5.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.054 $X2=0.837 $Y2=0.111
r167 16 97 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r168 16 19 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2295
r169 13 92 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r170 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r171 5 87 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.151 $Y2=0.135
r172 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r173 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%D 2 5 7 10 12 18 25 27 28 32 VSS
c20 32 VSS 0.00973151f $X=0.243 $Y=0.135
c21 28 VSS 2.45662e-20 $X=0.276 $Y=0.135
c22 27 VSS 7.4587e-19 $X=0.271 $Y=0.135
c23 25 VSS 2.67956e-19 $X=0.281 $Y=0.135
c24 18 VSS 1.8908e-19 $X=0.243 $Y=0.123
c25 16 VSS 7.25127e-19 $X=0.243 $Y=0.119
c26 12 VSS 0.0088416f $X=0.244 $Y=0.082
c27 10 VSS 1.58648e-20 $X=0.243 $Y=0.126
c28 5 VSS 0.0044978f $X=0.297 $Y=0.135
c29 2 VSS 0.0630445f $X=0.297 $Y=0.0675
r30 27 28 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.271
+ $Y=0.135 $X2=0.276 $Y2=0.135
r31 25 28 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.281
+ $Y=0.135 $X2=0.276 $Y2=0.135
r32 25 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.281 $Y=0.135 $X2=0.281
+ $Y2=0.135
r33 23 32 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.243 $Y2=0.135
r34 23 27 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.271 $Y2=0.135
r35 17 18 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.12 $X2=0.243 $Y2=0.123
r36 16 17 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.119 $X2=0.243 $Y2=0.12
r37 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.101 $X2=0.243 $Y2=0.119
r38 12 15 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.082 $X2=0.243 $Y2=0.101
r39 10 32 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.135
r40 10 18 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.123
r41 5 26 14.5455 $w=2.2e-08 $l=1.6e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.281 $Y2=0.135
r42 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r43 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%6 2 5 7 10 13 15 17 22 28 33 35 39 44 45 46
+ 55 57 58 59 60 64 69 79 80 81 82 87 95 VSS
c88 95 VSS 1.18012e-19 $X=0.891 $Y=0.173
c89 87 VSS 1.14917e-19 $X=0.405 $Y=0.178
c90 82 VSS 2.91958e-19 $X=0.189 $Y=0.182
c91 81 VSS 6.57126e-19 $X=0.189 $Y=0.167
c92 80 VSS 3.57675e-19 $X=0.189 $Y=0.106
c93 79 VSS 6.66951e-19 $X=0.189 $Y=0.088
c94 69 VSS 4.80366e-19 $X=0.891 $Y=0.111
c95 64 VSS 6.02738e-19 $X=0.405 $Y=0.135
c96 60 VSS 6.08738e-19 $X=0.852 $Y=0.189
c97 59 VSS 0.0164984f $X=0.741 $Y=0.189
c98 58 VSS 9.11862e-19 $X=0.891 $Y=0.189
c99 57 VSS 8.85234e-19 $X=0.891 $Y=0.189
c100 55 VSS 6.83354e-19 $X=0.405 $Y=0.189
c101 46 VSS 0.00169555f $X=0.18 $Y=0.234
c102 45 VSS 7.95076e-19 $X=0.189 $Y=0.225
c103 44 VSS 0.00196236f $X=0.189 $Y=0.234
c104 39 VSS 0.00193333f $X=0.162 $Y=0.234
c105 35 VSS 0.00170883f $X=0.18 $Y=0.036
c106 33 VSS 0.00196236f $X=0.189 $Y=0.036
c107 28 VSS 0.00193426f $X=0.162 $Y=0.036
c108 25 VSS 0.0072389f $X=0.16 $Y=0.216
c109 20 VSS 0.00719538f $X=0.16 $Y=0.054
c110 13 VSS 0.00184946f $X=0.891 $Y=0.111
c111 10 VSS 0.0589399f $X=0.891 $Y=0.0405
c112 5 VSS 0.00171178f $X=0.405 $Y=0.135
c113 2 VSS 0.0598132f $X=0.405 $Y=0.054
r114 94 95 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.167 $X2=0.891 $Y2=0.173
r115 86 87 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.167 $X2=0.405 $Y2=0.178
r116 81 82 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.167 $X2=0.189 $Y2=0.182
r117 80 81 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.106 $X2=0.189 $Y2=0.167
r118 79 80 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.088 $X2=0.189 $Y2=0.106
r119 69 94 3.80247 $w=1.8e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.111 $X2=0.891 $Y2=0.167
r120 64 86 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.167
r121 59 60 7.53704 $w=1.8e-08 $l=1.11e-07 $layer=M2 $thickness=3.6e-08 $X=0.741
+ $Y=0.189 $X2=0.852 $Y2=0.189
r122 58 95 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.189 $X2=0.891 $Y2=0.173
r123 57 60 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M2 $thickness=3.6e-08 $X=0.891
+ $Y=0.189 $X2=0.852 $Y2=0.189
r124 57 58 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.891 $Y=0.189 $X2=0.891
+ $Y2=0.189
r125 55 87 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.178
r126 54 59 22.8148 $w=1.8e-08 $l=3.36e-07 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.741 $Y2=0.189
r127 54 55 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.189 $X2=0.405
+ $Y2=0.189
r128 51 82 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.182
r129 50 54 14.6667 $w=1.8e-08 $l=2.16e-07 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.405 $Y2=0.189
r130 50 51 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.189 $X2=0.189
+ $Y2=0.189
r131 46 47 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r132 45 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.189
r133 44 47 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r134 44 45 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.189 $Y2=0.225
r135 39 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r136 35 36 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r137 34 79 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.088
r138 33 36 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r139 33 34 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.189 $Y2=0.045
r140 28 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r141 25 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r142 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r143 20 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r144 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r145 13 69 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.111 $X2=0.891
+ $Y2=0.111
r146 13 15 393.383 $w=2e-08 $l=1.05e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.111 $X2=0.891 $Y2=0.216
r147 10 13 264.128 $w=2e-08 $l=7.05e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.0405 $X2=0.891 $Y2=0.111
r148 5 64 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r149 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r150 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.054 $X2=0.405 $Y2=0.135
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%7 2 5 7 9 10 13 14 19 22 24 27 29 32 34 36
+ 40 42 43 45 46 47 49 55 56 57 58 59 60 61 62 64 68 69 70 75 78 79 80 81 101
+ 102 107 108 VSS
c95 108 VSS 5.17586e-19 $X=0.9875 $Y=0.225
c96 107 VSS 0.00158131f $X=0.981 $Y=0.225
c97 102 VSS 0.0012042f $X=0.747 $Y=0.225
c98 101 VSS 0.00156761f $X=0.729 $Y=0.225
c99 81 VSS 4.0314e-19 $X=0.913 $Y=0.225
c100 80 VSS 0.00639706f $X=0.905 $Y=0.225
c101 79 VSS 0.00308534f $X=0.994 $Y=0.225
c102 78 VSS 0.00374447f $X=0.994 $Y=0.225
c103 75 VSS 0.00219963f $X=0.755 $Y=0.225
c104 72 VSS 0.001396f $X=0.702 $Y=0.225
c105 70 VSS 8.62592e-19 $X=0.972 $Y=0.192
c106 69 VSS 7.48816e-19 $X=0.972 $Y=0.168
c107 68 VSS 2.49198e-19 $X=0.972 $Y=0.103
c108 64 VSS 0.00136128f $X=0.972 $Y=0.045
c109 62 VSS 9.10211e-19 $X=0.972 $Y=0.216
c110 61 VSS 2.46855e-19 $X=0.702 $Y=0.203
c111 60 VSS 1.8406e-19 $X=0.702 $Y=0.198
c112 59 VSS 3.59086e-19 $X=0.702 $Y=0.18
c113 58 VSS 4.7981e-19 $X=0.702 $Y=0.173
c114 57 VSS 4.05265e-19 $X=0.702 $Y=0.133
c115 56 VSS 2.16238e-19 $X=0.702 $Y=0.126
c116 55 VSS 8.40434e-19 $X=0.702 $Y=0.108
c117 49 VSS 0.0016703f $X=0.702 $Y=0.072
c118 47 VSS 3.37877e-19 $X=0.702 $Y=0.216
c119 46 VSS 9.74819e-19 $X=0.6805 $Y=0.225
c120 45 VSS 0.00610521f $X=0.668 $Y=0.225
c121 44 VSS 3.32809e-19 $X=0.612 $Y=0.225
c122 43 VSS 0.00243626f $X=0.608 $Y=0.225
c123 42 VSS 0.00160765f $X=0.576 $Y=0.225
c124 41 VSS 8.65354e-19 $X=0.693 $Y=0.225
c125 40 VSS 1.62557e-19 $X=0.567 $Y=0.207
c126 36 VSS 2.41699e-19 $X=0.567 $Y=0.18
c127 34 VSS 1.53526e-19 $X=0.567 $Y=0.216
c128 32 VSS 0.0152717f $X=0.812 $Y=0.2295
c129 29 VSS 3.14771e-19 $X=0.827 $Y=0.2295
c130 27 VSS 3.29654e-19 $X=0.754 $Y=0.216
c131 22 VSS 0.0152898f $X=0.974 $Y=0.0405
c132 19 VSS 3.14771e-19 $X=0.989 $Y=0.0405
c133 17 VSS 3.52885e-19 $X=0.916 $Y=0.0405
c134 13 VSS 0.0084744f $X=0.702 $Y=0.0405
c135 9 VSS 6.29543e-19 $X=0.719 $Y=0.0405
c136 5 VSS 0.00205979f $X=0.567 $Y=0.18
c137 2 VSS 0.0609977f $X=0.567 $Y=0.054
r138 107 108 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.981 $Y=0.225 $X2=0.9875 $Y2=0.225
r139 104 107 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.225 $X2=0.981 $Y2=0.225
r140 101 102 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.225 $X2=0.747 $Y2=0.225
r141 80 81 0.54321 $w=1.8e-08 $l=8e-09 $layer=M2 $thickness=3.6e-08 $X=0.905
+ $Y=0.225 $X2=0.913 $Y2=0.225
r142 79 108 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.994
+ $Y=0.225 $X2=0.9875 $Y2=0.225
r143 78 81 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.994
+ $Y=0.225 $X2=0.913 $Y2=0.225
r144 78 79 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.994 $Y=0.225 $X2=0.994
+ $Y2=0.225
r145 75 102 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.755
+ $Y=0.225 $X2=0.747 $Y2=0.225
r146 74 80 10.1852 $w=1.8e-08 $l=1.5e-07 $layer=M2 $thickness=3.6e-08 $X=0.755
+ $Y=0.225 $X2=0.905 $Y2=0.225
r147 74 75 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.755 $Y=0.225 $X2=0.755
+ $Y2=0.225
r148 71 101 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.711
+ $Y=0.225 $X2=0.729 $Y2=0.225
r149 71 72 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.711
+ $Y=0.225 $X2=0.702 $Y2=0.225
r150 69 70 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.168 $X2=0.972 $Y2=0.192
r151 68 69 4.41358 $w=1.8e-08 $l=6.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.103 $X2=0.972 $Y2=0.168
r152 67 68 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.054 $X2=0.972 $Y2=0.103
r153 64 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.045 $X2=0.972 $Y2=0.054
r154 62 104 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.216 $X2=0.972 $Y2=0.225
r155 62 70 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.216 $X2=0.972 $Y2=0.192
r156 60 61 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.198 $X2=0.702 $Y2=0.203
r157 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.18 $X2=0.702 $Y2=0.198
r158 58 59 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.173 $X2=0.702 $Y2=0.18
r159 57 58 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.133 $X2=0.702 $Y2=0.173
r160 56 57 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.126 $X2=0.702 $Y2=0.133
r161 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.108 $X2=0.702 $Y2=0.126
r162 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.09 $X2=0.702 $Y2=0.108
r163 49 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.072 $X2=0.702 $Y2=0.09
r164 49 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.072
+ $X2=0.702 $Y2=0.072
r165 47 72 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.216 $X2=0.702 $Y2=0.225
r166 47 61 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.216 $X2=0.702 $Y2=0.203
r167 45 46 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.668
+ $Y=0.225 $X2=0.6805 $Y2=0.225
r168 44 45 3.80247 $w=1.8e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.225 $X2=0.668 $Y2=0.225
r169 43 44 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.608
+ $Y=0.225 $X2=0.612 $Y2=0.225
r170 42 43 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.225 $X2=0.608 $Y2=0.225
r171 41 72 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.225 $X2=0.702 $Y2=0.225
r172 41 46 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.693
+ $Y=0.225 $X2=0.6805 $Y2=0.225
r173 39 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.198 $X2=0.567 $Y2=0.207
r174 36 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.18 $X2=0.567 $Y2=0.198
r175 34 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.567 $Y=0.216 $X2=0.576 $Y2=0.225
r176 34 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.216 $X2=0.567 $Y2=0.207
r177 29 32 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.2295 $X2=0.812 $Y2=0.2295
r178 27 32 22.2487 $w=5.4e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.754
+ $Y=0.216 $X2=0.812 $Y2=0.216
r179 27 75 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.225
+ $X2=0.756 $Y2=0.225
r180 24 27 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.216 $X2=0.754 $Y2=0.216
r181 22 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.045
+ $X2=0.972 $Y2=0.045
r182 19 22 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.989 $Y=0.0405 $X2=0.974 $Y2=0.0405
r183 17 22 42.963 $w=2.7e-08 $l=5.6e-08 $layer=LISD $thickness=2.8e-08 $X=0.916
+ $Y=0.0405 $X2=0.972 $Y2=0.0405
r184 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.0405 $X2=0.916 $Y2=0.0405
r185 13 50 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.702 $Y=0.0405 $X2=0.702 $Y2=0.072
r186 10 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.0405 $X2=0.702 $Y2=0.0405
r187 9 13 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.0405 $X2=0.702 $Y2=0.0405
r188 5 36 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.18 $X2=0.567
+ $Y2=0.18
r189 5 7 185.452 $w=2e-08 $l=4.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.18 $X2=0.567 $Y2=0.2295
r190 2 5 472.059 $w=2e-08 $l=1.26e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.054 $X2=0.567 $Y2=0.18
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%RESET 2 5 7 10 13 15 20 23 25 31 34 35 36 37
+ 38 39 40 41 57 58 VSS
c56 58 VSS 2.39249e-19 $X=0.638 $Y=0.117
c57 57 VSS 4.47202e-19 $X=0.63 $Y=0.117
c58 41 VSS 4.67084e-19 $X=0.983 $Y=0.117
c59 40 VSS 1.0352e-19 $X=0.913 $Y=0.117
c60 39 VSS 5.31777e-19 $X=0.905 $Y=0.117
c61 38 VSS 6.29272e-19 $X=0.852 $Y=0.117
c62 37 VSS 0.00107354f $X=0.778 $Y=0.117
c63 36 VSS 0.00121746f $X=0.752 $Y=0.117
c64 35 VSS 0.00103588f $X=1.053 $Y=0.117
c65 34 VSS 8.22015e-19 $X=1.053 $Y=0.117
c66 31 VSS 0.00106328f $X=0.646 $Y=0.117
c67 25 VSS 2.01705e-20 $X=0.621 $Y=0.167
c68 23 VSS 0.0024511f $X=0.622 $Y=0.17
c69 20 VSS 2.25553e-19 $X=0.621 $Y=0.159
c70 13 VSS 0.00202958f $X=1.053 $Y=0.135
c71 10 VSS 0.0568294f $X=1.053 $Y=0.0405
c72 5 VSS 0.00219384f $X=0.621 $Y=0.159
c73 2 VSS 0.0576659f $X=0.621 $Y=0.054
r74 57 58 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.117 $X2=0.638 $Y2=0.117
r75 54 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.117 $X2=0.63 $Y2=0.117
r76 40 41 4.75309 $w=1.8e-08 $l=7e-08 $layer=M2 $thickness=3.6e-08 $X=0.913
+ $Y=0.117 $X2=0.983 $Y2=0.117
r77 39 40 0.54321 $w=1.8e-08 $l=8e-09 $layer=M2 $thickness=3.6e-08 $X=0.905
+ $Y=0.117 $X2=0.913 $Y2=0.117
r78 38 39 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.852
+ $Y=0.117 $X2=0.905 $Y2=0.117
r79 37 38 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.778
+ $Y=0.117 $X2=0.852 $Y2=0.117
r80 36 37 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.752
+ $Y=0.117 $X2=0.778 $Y2=0.117
r81 34 41 4.75309 $w=1.8e-08 $l=7e-08 $layer=M2 $thickness=3.6e-08 $X=1.053
+ $Y=0.117 $X2=0.983 $Y2=0.117
r82 34 35 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.053 $Y=0.117 $X2=1.053
+ $Y2=0.117
r83 31 58 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.646
+ $Y=0.117 $X2=0.638 $Y2=0.117
r84 30 36 7.19753 $w=1.8e-08 $l=1.06e-07 $layer=M2 $thickness=3.6e-08 $X=0.646
+ $Y=0.117 $X2=0.752 $Y2=0.117
r85 30 31 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.646 $Y=0.117 $X2=0.646
+ $Y2=0.117
r86 24 25 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.164 $X2=0.621 $Y2=0.167
r87 23 25 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.17 $X2=0.621 $Y2=0.167
r88 20 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.159 $X2=0.621 $Y2=0.164
r89 17 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.126 $X2=0.621 $Y2=0.117
r90 17 20 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.126 $X2=0.621 $Y2=0.159
r91 13 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.053 $Y=0.135 $X2=1.053
+ $Y2=0.135
r92 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.135 $X2=1.053 $Y2=0.216
r93 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.053
+ $Y=0.0405 $X2=1.053 $Y2=0.135
r94 5 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.159 $X2=0.621
+ $Y2=0.159
r95 5 7 264.128 $w=2e-08 $l=7.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.159 $X2=0.621 $Y2=0.2295
r96 2 5 393.383 $w=2e-08 $l=1.05e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.054 $X2=0.621 $Y2=0.159
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%9 2 5 7 10 11 17 18 22 23 26 31 32 34 37 38
+ 39 40 41 44 48 50 51 52 53 VSS
c62 53 VSS 0.00185157f $X=0.685 $Y=0.081
c63 52 VSS 0.00634256f $X=0.632 $Y=0.081
c64 51 VSS 0.00165917f $X=0.738 $Y=0.081
c65 50 VSS 0.00295505f $X=0.738 $Y=0.081
c66 48 VSS 0.00318414f $X=0.521 $Y=0.081
c67 44 VSS 0.00164955f $X=0.378 $Y=0.081
c68 41 VSS 4.60428e-19 $X=0.504 $Y=0.081
c69 40 VSS 6.90371e-19 $X=0.495 $Y=0.203
c70 39 VSS 4.15852e-20 $X=0.495 $Y=0.167
c71 38 VSS 0.00129811f $X=0.495 $Y=0.164
c72 37 VSS 6.61901e-19 $X=0.495 $Y=0.119
c73 36 VSS 3.1486e-19 $X=0.495 $Y=0.108
c74 35 VSS 4.96683e-19 $X=0.495 $Y=0.101
c75 34 VSS 4.03342e-19 $X=0.495 $Y=0.225
c76 32 VSS 0.00146362f $X=0.468 $Y=0.234
c77 31 VSS 0.00343063f $X=0.45 $Y=0.234
c78 26 VSS 0.00404036f $X=0.486 $Y=0.234
c79 25 VSS 5.70081e-19 $X=0.432 $Y=0.2295
c80 22 VSS 0.00247374f $X=0.432 $Y=0.2025
c81 19 VSS 7.52159e-20 $X=0.4275 $Y=0.216
c82 17 VSS 0.0030948f $X=0.378 $Y=0.0675
c83 12 VSS 6.4484e-19 $X=0.378 $Y=0.0455
c84 5 VSS 0.00448045f $X=0.729 $Y=0.11
c85 2 VSS 0.058429f $X=0.729 $Y=0.0405
r86 52 53 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.632
+ $Y=0.081 $X2=0.685 $Y2=0.081
r87 51 58 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.081 $X2=0.738 $Y2=0.11
r88 50 53 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.738
+ $Y=0.081 $X2=0.685 $Y2=0.081
r89 50 51 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.738 $Y=0.081 $X2=0.738
+ $Y2=0.081
r90 47 52 7.53704 $w=1.8e-08 $l=1.11e-07 $layer=M2 $thickness=3.6e-08 $X=0.521
+ $Y=0.081 $X2=0.632 $Y2=0.081
r91 47 48 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.521 $Y=0.081 $X2=0.521
+ $Y2=0.081
r92 43 47 9.70988 $w=1.8e-08 $l=1.43e-07 $layer=M2 $thickness=3.6e-08 $X=0.378
+ $Y=0.081 $X2=0.521 $Y2=0.081
r93 43 44 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.378 $Y=0.081 $X2=0.378
+ $Y2=0.081
r94 41 48 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.081 $X2=0.521 $Y2=0.081
r95 39 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.167 $X2=0.495 $Y2=0.203
r96 38 39 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.164 $X2=0.495 $Y2=0.167
r97 37 38 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.119 $X2=0.495 $Y2=0.164
r98 36 37 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.108 $X2=0.495 $Y2=0.119
r99 35 36 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.101 $X2=0.495 $Y2=0.108
r100 34 40 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.225 $X2=0.495 $Y2=0.203
r101 33 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.495 $Y=0.09 $X2=0.504 $Y2=0.081
r102 33 35 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.09 $X2=0.495 $Y2=0.101
r103 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r104 28 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.45 $Y2=0.234
r105 26 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.486 $Y=0.234 $X2=0.495 $Y2=0.225
r106 26 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.468 $Y2=0.234
r107 23 25 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2295 $X2=0.432 $Y2=0.2295
r108 22 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r109 19 25 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.216 $X2=0.432 $Y2=0.2295
r110 19 22 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.216 $X2=0.4275 $Y2=0.189
r111 18 22 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.189 $X2=0.4275 $Y2=0.189
r112 17 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.085
+ $X2=0.378 $Y2=0.085
r113 11 12 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0455 $X2=0.378 $Y2=0.0455
r114 10 12 15.7779 $w=3.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.0455 $X2=0.378 $Y2=0.0455
r115 9 17 3.12934 $w=6.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.378 $Y=0.064 $X2=0.361 $Y2=0.064
r116 9 12 5.40574 $w=7.4e-08 $l=1.85e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.378 $Y=0.064 $X2=0.378 $Y2=0.0455
r117 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.738 $Y=0.11 $X2=0.738
+ $Y2=0.11
r118 5 7 397.129 $w=2e-08 $l=1.06e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.11 $X2=0.729 $Y2=0.216
r119 2 5 260.382 $w=2e-08 $l=6.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0405 $X2=0.729 $Y2=0.11
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%SET 2 7 10 16 19 21 34 38 41 VSS
c64 41 VSS 2.82896e-19 $X=0.783 $Y=0.146
c65 38 VSS 4.04314e-19 $X=0.783 $Y=0.159
c66 34 VSS 0.00148115f $X=0.782 $Y=0.132
c67 26 VSS 1.2365e-19 $X=0.6755 $Y=0.159
c68 19 VSS 0.0245757f $X=0.999 $Y=0.159
c69 16 VSS 0.0586646f $X=0.999 $Y=0.0405
c70 13 VSS 1.08403e-20 $X=0.783 $Y=0.159
c71 10 VSS 0.0586794f $X=0.783 $Y=0.054
c72 2 VSS 0.0585363f $X=0.675 $Y=0.0405
r73 40 41 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.133 $X2=0.783 $Y2=0.146
r74 38 41 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.159 $X2=0.783 $Y2=0.146
r75 34 40 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.132 $X2=0.783 $Y2=0.133
r76 19 21 213.551 $w=2e-08 $l=5.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.159 $X2=0.999 $Y2=0.216
r77 16 19 443.961 $w=2e-08 $l=1.185e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0405 $X2=0.999 $Y2=0.159
r78 13 19 186.429 $w=2.4e-08 $l=2.16e-07 $layer=LISD $thickness=2.8e-08 $X=0.783
+ $Y=0.159 $X2=0.999 $Y2=0.159
r79 13 26 92.7827 $w=2.4e-08 $l=1.075e-07 $layer=LISD $thickness=2.8e-08
+ $X=0.783 $Y=0.159 $X2=0.6755 $Y2=0.159
r80 13 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.783 $Y=0.159 $X2=0.783
+ $Y2=0.159
r81 13 38 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.159 $X2=0.783
+ $Y2=0.159
r82 10 13 393.383 $w=2e-08 $l=1.05e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.054 $X2=0.783 $Y2=0.159
r83 5 26 0.416667 $w=2.4e-08 $l=5e-10 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.159 $X2=0.6755 $Y2=0.159
r84 5 7 213.551 $w=2e-08 $l=5.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.159 $X2=0.675 $Y2=0.216
r85 2 5 443.961 $w=2e-08 $l=1.185e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0405 $X2=0.675 $Y2=0.159
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%11 2 5 7 10 13 15 17 18 21 22 23 26 27 32 33
+ 37 42 43 45 47 52 57 68 69 72 73 74 76 77 VSS
c70 77 VSS 3.97453e-19 $X=0.927 $Y=0.097
c71 76 VSS 4.37533e-19 $X=0.927 $Y=0.09
c72 75 VSS 1.24394e-19 $X=0.927 $Y=0.072
c73 74 VSS 8.64013e-20 $X=0.927 $Y=0.067
c74 73 VSS 4.06594e-20 $X=0.927 $Y=0.058
c75 72 VSS 2.92134e-20 $X=0.927 $Y=0.054
c76 69 VSS 0.00136895f $X=0.927 $Y=0.201
c77 68 VSS 0.00390486f $X=0.927 $Y=0.201
c78 57 VSS 0.00268841f $X=1.323 $Y=0.135
c79 52 VSS 0.00104826f $X=1.107 $Y=0.135
c80 48 VSS 0.00415682f $X=1.2605 $Y=0.153
c81 47 VSS 0.00496673f $X=1.198 $Y=0.153
c82 45 VSS 0.00598828f $X=1.323 $Y=0.153
c83 43 VSS 0.00259454f $X=1.067 $Y=0.153
c84 42 VSS 7.50229e-19 $X=1.008 $Y=0.153
c85 37 VSS 5.84953e-19 $X=0.927 $Y=0.153
c86 33 VSS 0.00126587f $X=0.9 $Y=0.039
c87 32 VSS 0.0025837f $X=0.882 $Y=0.039
c88 27 VSS 0.00357014f $X=0.918 $Y=0.039
c89 26 VSS 0.00314137f $X=0.864 $Y=0.216
c90 22 VSS 8.61759e-19 $X=0.881 $Y=0.216
c91 21 VSS 0.00159741f $X=0.864 $Y=0.054
c92 17 VSS 7.24097e-19 $X=0.881 $Y=0.0405
c93 13 VSS 0.00296536f $X=1.323 $Y=0.135
c94 10 VSS 0.0656672f $X=1.323 $Y=0.0675
c95 5 VSS 0.00193028f $X=1.107 $Y=0.135
c96 2 VSS 0.0575145f $X=1.107 $Y=0.0405
r97 76 77 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.927
+ $Y=0.09 $X2=0.927 $Y2=0.097
r98 75 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.927
+ $Y=0.072 $X2=0.927 $Y2=0.09
r99 74 75 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.927
+ $Y=0.067 $X2=0.927 $Y2=0.072
r100 73 74 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.927
+ $Y=0.058 $X2=0.927 $Y2=0.067
r101 72 73 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.927
+ $Y=0.054 $X2=0.927 $Y2=0.058
r102 68 69 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.927 $Y=0.201
+ $X2=0.927 $Y2=0.201
r103 61 68 44.0179 $w=2.4e-08 $l=5.1e-08 $layer=LISD $thickness=2.8e-08 $X=0.876
+ $Y=0.201 $X2=0.927 $Y2=0.201
r104 47 48 4.24383 $w=1.8e-08 $l=6.25e-08 $layer=M2 $thickness=3.6e-08 $X=1.198
+ $Y=0.153 $X2=1.2605 $Y2=0.153
r105 45 48 4.24383 $w=1.8e-08 $l=6.25e-08 $layer=M2 $thickness=3.6e-08 $X=1.323
+ $Y=0.153 $X2=1.2605 $Y2=0.153
r106 45 57 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.323 $Y=0.153 $X2=1.323
+ $Y2=0.153
r107 42 43 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M2 $thickness=3.6e-08 $X=1.008
+ $Y=0.153 $X2=1.067 $Y2=0.153
r108 40 47 6.17901 $w=1.8e-08 $l=9.1e-08 $layer=M2 $thickness=3.6e-08 $X=1.107
+ $Y=0.153 $X2=1.198 $Y2=0.153
r109 40 43 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=1.107
+ $Y=0.153 $X2=1.067 $Y2=0.153
r110 40 52 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.107 $Y=0.153 $X2=1.107
+ $Y2=0.153
r111 37 69 3.25926 $w=1.8e-08 $l=4.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.927
+ $Y=0.153 $X2=0.927 $Y2=0.201
r112 37 77 3.80247 $w=1.8e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.927
+ $Y=0.153 $X2=0.927 $Y2=0.097
r113 36 42 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.927
+ $Y=0.153 $X2=1.008 $Y2=0.153
r114 36 37 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.927 $Y=0.153 $X2=0.927
+ $Y2=0.153
r115 34 72 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.927
+ $Y=0.048 $X2=0.927 $Y2=0.054
r116 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.039 $X2=0.9 $Y2=0.039
r117 29 32 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.867
+ $Y=0.039 $X2=0.882 $Y2=0.039
r118 27 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.918 $Y=0.039 $X2=0.927 $Y2=0.048
r119 27 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.039 $X2=0.9 $Y2=0.039
r120 26 61 1.21653 $w=2.4e-08 $l=1.2e-08 $layer=LISD $thickness=2.8e-08 $X=0.864
+ $Y=0.201 $X2=0.876 $Y2=0.201
r121 23 26 21.6244 $w=4.675e-08 $l=2.27706e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2295 $X2=0.864 $Y2=0.216
r122 22 26 13.4224 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.216 $X2=0.864 $Y2=0.216
r123 21 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.867 $Y=0.039
+ $X2=0.867 $Y2=0.039
r124 18 21 13.4224 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.054 $X2=0.864 $Y2=0.054
r125 17 21 21.6244 $w=4.675e-08 $l=2.27706e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0405 $X2=0.864 $Y2=0.054
r126 13 57 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.323 $Y=0.135 $X2=1.323
+ $Y2=0.135
r127 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.135 $X2=1.323 $Y2=0.2025
r128 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.0675 $X2=1.323 $Y2=0.135
r129 5 52 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.107 $Y=0.135 $X2=1.107
+ $Y2=0.135
r130 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.107
+ $Y=0.135 $X2=1.107 $Y2=0.216
r131 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=1.107
+ $Y=0.0405 $X2=1.107 $Y2=0.135
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%12 1 3 5 9 15 18 21 24 33 34 37 38 VSS
c34 41 VSS 3.19801e-19 $X=1.132 $Y=0.216
c35 37 VSS 0.0335604f $X=1.08 $Y=0.0405
c36 33 VSS 6.29543e-19 $X=1.097 $Y=0.0405
c37 24 VSS 0.00969151f $X=1.161 $Y=0.2
c38 21 VSS 0.0625575f $X=1.161 $Y=0.0405
c39 15 VSS 0.0609503f $X=0.945 $Y=0.096
c40 13 VSS 0.0217413f $X=1.08 $Y=0.096
c41 9 VSS 0.0416987f $X=1.1605 $Y=0.189
c42 5 VSS 0.0128386f $X=1.146 $Y=0.096
c43 3 VSS 4.73091e-19 $X=0.9455 $Y=0.096
c44 1 VSS 0.00605869f $X=1.068 $Y=0.096
r45 38 41 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.117 $Y=0.216 $X2=1.132 $Y2=0.216
r46 34 37 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.0405 $X2=1.08 $Y2=0.0405
r47 33 37 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.097 $Y=0.0405 $X2=1.08 $Y2=0.0405
r48 24 41 9.33602 $w=3.55e-08 $l=1.6e-08 $layer=LISD $thickness=2.8e-08 $X=1.146
+ $Y=0.2 $X2=1.146 $Y2=0.216
r49 21 24 597.567 $w=2e-08 $l=1.595e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.161 $Y=0.0405 $X2=1.161 $Y2=0.2
r50 15 18 449.58 $w=2e-08 $l=1.2e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.945
+ $Y=0.096 $X2=0.945 $Y2=0.216
r51 12 37 37.5446 $w=2.4e-08 $l=4.35e-08 $layer=LISD $thickness=2.8e-08 $X=1.08
+ $Y=0.084 $X2=1.08 $Y2=0.0405
r52 12 13 2.27953 $w=4.8e-08 $l=1.2e-08 $layer=LISD $thickness=2.8e-08 $X=1.08
+ $Y=0.084 $X2=1.08 $Y2=0.096
r53 9 24 7.94115 $w=3.55e-08 $l=1.76635e-08 $layer=LISD $thickness=2.8e-08
+ $X=1.159 $Y=0.189 $X2=1.146 $Y2=0.2
r54 9 24 9.56522 $w=2.3e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=1.1605
+ $Y=0.189 $X2=1.1605 $Y2=0.2
r55 7 9 36.6696 $w=4.9e-08 $l=8.1e-08 $layer=LISD $thickness=2.8e-08 $X=1.159
+ $Y=0.108 $X2=1.159 $Y2=0.189
r56 6 13 8.77136 $w=2.4e-08 $l=1.2e-08 $layer=LISD $thickness=2.8e-08 $X=1.092
+ $Y=0.096 $X2=1.08 $Y2=0.096
r57 5 7 11.5978 $w=2.6e-08 $l=1.80278e-08 $layer=LISD $thickness=2.8e-08
+ $X=1.146 $Y=0.096 $X2=1.159 $Y2=0.108
r58 5 6 46.6071 $w=2.4e-08 $l=5.4e-08 $layer=LISD $thickness=2.8e-08 $X=1.146
+ $Y=0.096 $X2=1.092 $Y2=0.096
r59 3 15 0.416667 $w=2.4e-08 $l=5e-10 $layer=LIG $thickness=5e-08 $X=0.9455
+ $Y=0.096 $X2=0.945 $Y2=0.096
r60 1 13 8.77136 $w=2.4e-08 $l=1.2e-08 $layer=LISD $thickness=2.8e-08 $X=1.068
+ $Y=0.096 $X2=1.08 $Y2=0.096
r61 1 3 105.729 $w=2.4e-08 $l=1.225e-07 $layer=LISD $thickness=2.8e-08 $X=1.068
+ $Y=0.096 $X2=0.9455 $Y2=0.096
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%13 1 4 6 7 10 12 21 23 24 25 VSS
c12 25 VSS 0.00167049f $X=0.576 $Y=0.036
c13 24 VSS 0.00179001f $X=0.558 $Y=0.036
c14 23 VSS 0.00773487f $X=0.547 $Y=0.036
c15 22 VSS 0.00173283f $X=0.486 $Y=0.036
c16 21 VSS 0.00147791f $X=0.468 $Y=0.036
c17 20 VSS 0.00229295f $X=0.45 $Y=0.036
c18 18 VSS 0.00408509f $X=0.594 $Y=0.036
c19 12 VSS 0.0017807f $X=0.432 $Y=0.036
c20 10 VSS 0.00821636f $X=0.594 $Y=0.054
c21 6 VSS 5.65078e-19 $X=0.611 $Y=0.054
c22 4 VSS 0.00359891f $X=0.43 $Y=0.054
r23 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.576 $Y2=0.036
r24 23 24 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.547
+ $Y=0.036 $X2=0.558 $Y2=0.036
r25 22 23 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.547 $Y2=0.036
r26 21 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.486 $Y2=0.036
r27 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r28 18 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.576 $Y2=0.036
r29 12 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r30 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036 $X2=0.594
+ $Y2=0.036
r31 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.054 $X2=0.594 $Y2=0.054
r32 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.054 $X2=0.594 $Y2=0.054
r33 4 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r34 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.054 $X2=0.43 $Y2=0.054
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%14 1 2 5 6 13 16 17 18 19 VSS
c26 19 VSS 0.00272102f $X=1.1255 $Y=0.045
c27 18 VSS 0.0119822f $X=1.067 $Y=0.045
c28 17 VSS 0.00427953f $X=1.184 $Y=0.045
c29 16 VSS 0.00293942f $X=1.184 $Y=0.045
c30 13 VSS 0.00389734f $X=0.792 $Y=0.045
c31 9 VSS 0.00326847f $X=1.186 $Y=0.0405
c32 5 VSS 0.00361464f $X=0.81 $Y=0.054
c33 1 VSS 7.0838e-19 $X=0.827 $Y=0.054
r34 18 19 3.97222 $w=1.8e-08 $l=5.85e-08 $layer=M2 $thickness=3.6e-08 $X=1.067
+ $Y=0.045 $X2=1.1255 $Y2=0.045
r35 16 19 3.97222 $w=1.8e-08 $l=5.85e-08 $layer=M2 $thickness=3.6e-08 $X=1.184
+ $Y=0.045 $X2=1.1255 $Y2=0.045
r36 16 17 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=1.184 $Y=0.045 $X2=1.184
+ $Y2=0.045
r37 12 18 18.6728 $w=1.8e-08 $l=2.75e-07 $layer=M2 $thickness=3.6e-08 $X=0.792
+ $Y=0.045 $X2=1.067 $Y2=0.045
r38 12 13 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.792 $Y=0.045 $X2=0.792
+ $Y2=0.045
r39 9 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.188 $Y=0.045 $X2=1.188
+ $Y2=0.045
r40 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.171
+ $Y=0.0405 $X2=1.186 $Y2=0.0405
r41 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.045 $X2=0.81
+ $Y2=0.045
r42 2 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.793
+ $Y=0.054 $X2=0.81 $Y2=0.054
r43 1 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.827
+ $Y=0.054 $X2=0.81 $Y2=0.054
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%QN 1 6 14 21 VSS
c4 32 VSS 0.00447704f $X=1.368 $Y=0.234
c5 31 VSS 0.00278493f $X=1.377 $Y=0.234
c6 24 VSS 0.0044068f $X=1.368 $Y=0.036
c7 23 VSS 0.00278493f $X=1.377 $Y=0.036
c8 21 VSS 0.00646566f $X=1.35 $Y=0.036
c9 18 VSS 9.37071e-21 $X=1.377 $Y=0.168
c10 16 VSS 0.00135133f $X=1.377 $Y=0.09
c11 15 VSS 8.61213e-19 $X=1.377 $Y=0.054
c12 14 VSS 0.00347148f $X=1.377 $Y=0.15
c13 12 VSS 0.00258899f $X=1.377 $Y=0.225
c14 9 VSS 0.00695944f $X=1.348 $Y=0.2025
c15 4 VSS 3.7894e-19 $X=1.348 $Y=0.0675
r16 32 33 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.368
+ $Y=0.234 $X2=1.3725 $Y2=0.234
r17 31 33 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.234 $X2=1.3725 $Y2=0.234
r18 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.35
+ $Y=0.234 $X2=1.368 $Y2=0.234
r19 24 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.368
+ $Y=0.036 $X2=1.3725 $Y2=0.036
r20 23 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.036 $X2=1.3725 $Y2=0.036
r21 20 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.35
+ $Y=0.036 $X2=1.368 $Y2=0.036
r22 20 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.35 $Y=0.036 $X2=1.35
+ $Y2=0.036
r23 17 18 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.167 $X2=1.377 $Y2=0.168
r24 15 16 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.054 $X2=1.377 $Y2=0.09
r25 14 17 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.15 $X2=1.377 $Y2=0.167
r26 14 16 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.15 $X2=1.377 $Y2=0.09
r27 12 31 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.225 $X2=1.377 $Y2=0.234
r28 12 18 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.225 $X2=1.377 $Y2=0.168
r29 11 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.045 $X2=1.377 $Y2=0.036
r30 11 15 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.377
+ $Y=0.045 $X2=1.377 $Y2=0.054
r31 9 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.35 $Y=0.234 $X2=1.35
+ $Y2=0.234
r32 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=1.333
+ $Y=0.2025 $X2=1.348 $Y2=0.2025
r33 4 21 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.35
+ $Y=0.0675 $X2=1.35 $Y2=0.036
r34 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.333
+ $Y=0.0675 $X2=1.348 $Y2=0.0675
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%16 1 6 9 VSS
c9 9 VSS 0.0197342f $X=0.38 $Y=0.2025
c10 6 VSS 3.25039e-19 $X=0.395 $Y=0.2025
c11 4 VSS 3.25039e-19 $X=0.322 $Y=0.2025
r12 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.2025 $X2=0.38 $Y2=0.2025
r13 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.2025 $X2=0.38 $Y2=0.2025
r14 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2025 $X2=0.322 $Y2=0.2025
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%17 1 6 9 VSS
c5 9 VSS 0.0212112f $X=0.542 $Y=0.2295
c6 6 VSS 3.14771e-19 $X=0.557 $Y=0.2295
c7 4 VSS 2.84146e-19 $X=0.484 $Y=0.2295
r8 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.557
+ $Y=0.2295 $X2=0.542 $Y2=0.2295
r9 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.484
+ $Y=0.2295 $X2=0.542 $Y2=0.2295
r10 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.2295 $X2=0.484 $Y2=0.2295
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%18 1 2 VSS
c0 1 VSS 0.00221026f $X=0.341 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.0675 $X2=0.307 $Y2=0.0675
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%19 1 2 VSS
c1 1 VSS 0.00225397f $X=0.611 $Y=0.2295
r2 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.611
+ $Y=0.2295 $X2=0.577 $Y2=0.2295
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%20 1 2 VSS
c3 1 VSS 0.00265637f $X=0.719 $Y=0.216
r4 1 2 25.1852 $w=5.4e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.216 $X2=0.685 $Y2=0.216
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%21 1 2 VSS
c1 1 VSS 0.00245075f $X=0.935 $Y=0.216
r2 1 2 25.1852 $w=5.4e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.935
+ $Y=0.216 $X2=0.901 $Y2=0.216
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%22 1 2 VSS
c4 1 VSS 0.00228377f $X=0.989 $Y=0.216
r5 1 2 25.1852 $w=5.4e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.216 $X2=0.955 $Y2=0.216
.ends

.subckt PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%23 1 2 VSS
c0 1 VSS 0.00217465f $X=1.097 $Y=0.216
r1 1 2 25.1852 $w=5.4e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=1.097
+ $Y=0.216 $X2=1.063 $Y2=0.216
.ends


* END of "./ASYNC_DFFHx1_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt ASYNC_DFFHx1_ASAP7_75t_SRAM  VSS VDD CLK D RESET SET QN
* 
* QN	QN
* SET	SET
* RESET	RESET
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_18_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_9_M3_d N_4_M3_g N_18_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 N_13_M4_d N_6_M4_g N_9_M4_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.395
+ $Y=0.027
M5 N_13_M5_d N_7_M5_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.557
+ $Y=0.027
M6 VSS N_RESET_M6_g N_13_M6_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.611
+ $Y=0.027
M7 N_7_M7_d N_SET_M7_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.665
+ $Y=0.027
M8 VSS N_9_M8_g N_7_M8_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.719 $Y=0.027
M9 N_14_M9_d N_SET_M9_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.773
+ $Y=0.027
M10 N_11_M10_d N_4_M10_g N_14_M10_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.827 $Y=0.027
M11 N_7_M11_d N_6_M11_g N_11_M11_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.881 $Y=0.027
M12 N_7_M12_d N_SET_M12_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.989
+ $Y=0.027
M13 N_12_M13_d N_RESET_M13_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.043
+ $Y=0.027
M14 VSS N_11_M14_g N_12_M14_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.097
+ $Y=0.027
M15 N_14_M15_d N_12_M15_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=1.151
+ $Y=0.027
M16 N_QN_M16_d N_11_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.027
M17 VDD N_CLK_M17_g N_4_M17_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M18 N_6_M18_d N_4_M18_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M19 N_16_M19_d N_D_M19_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M20 N_9_M20_d N_6_M20_g N_16_M20_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M21 N_17_M21_d N_4_M21_g N_9_M21_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.449 $Y=0.216
M22 N_19_M22_d N_7_M22_g N_17_M22_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.557 $Y=0.216
M23 VDD N_RESET_M23_g N_19_M23_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.611
+ $Y=0.216
M24 N_20_M24_d N_SET_M24_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.665
+ $Y=0.189
M25 N_7_M25_d N_9_M25_g N_20_M25_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.719 $Y=0.189
M26 N_11_M26_d N_4_M26_g N_7_M26_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.827 $Y=0.216
M27 N_21_M27_d N_6_M27_g N_11_M27_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.881 $Y=0.189
M28 N_22_M28_d N_12_M28_g N_21_M28_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.935 $Y=0.189
M29 VDD N_SET_M29_g N_22_M29_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.989
+ $Y=0.189
M30 N_23_M30_d N_RESET_M30_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=1.043
+ $Y=0.189
M31 N_12_M31_d N_11_M31_g N_23_M31_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
+ $X=1.097 $Y=0.189
M32 N_QN_M32_d N_11_M32_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.162
*
* 
* .include "ASYNC_DFFHx1_ASAP7_75t_SRAM.pex.sp.ASYNC_DFFHX1_ASAP7_75T_SRAM.pxi"
* BEGIN of "./ASYNC_DFFHx1_ASAP7_75t_SRAM.pex.sp.ASYNC_DFFHX1_ASAP7_75T_SRAM.pxi"
* File: ASYNC_DFFHx1_ASAP7_75t_SRAM.pex.sp.ASYNC_DFFHX1_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:17:25 2017
* 
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_13_p N_CLK_M17_g CLK
+ N_CLK_c_6_p VSS PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%CLK
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M18_g N_4_M3_g N_4_c_37_p
+ N_4_c_46_p N_4_M21_g N_4_M10_g N_4_c_50_p N_4_M26_g N_4_M0_s N_4_c_23_n
+ N_4_M17_s N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_28_n N_4_c_29_n
+ N_4_c_30_n N_4_c_31_n N_4_c_32_n N_4_c_41_p N_4_c_38_p N_4_c_56_p N_4_c_66_p
+ N_4_c_60_p N_4_c_71_p N_4_c_34_n N_4_c_35_n N_4_c_40_p N_4_c_59_p N_4_c_61_p
+ VSS PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%4
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_108_n N_D_M19_g N_D_c_125_p D
+ N_D_c_124_p N_D_c_111_n N_D_c_112_n N_D_c_113_n N_D_c_114_n VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%D
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%6 N_6_M4_g N_6_c_136_n N_6_M20_g N_6_M11_g
+ N_6_c_139_n N_6_M27_g N_6_M1_d N_6_M18_d N_6_c_127_n N_6_c_160_n N_6_c_141_n
+ N_6_c_128_n N_6_c_161_n N_6_c_129_n N_6_c_144_n N_6_c_145_n N_6_c_185_p
+ N_6_c_178_p N_6_c_130_n N_6_c_149_n N_6_c_151_n N_6_c_155_n N_6_c_131_n
+ N_6_c_132_n N_6_c_157_n N_6_c_133_n N_6_c_190_p N_6_c_201_p VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%6
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_217_n N_7_M22_g N_7_M8_s N_7_M7_d
+ N_7_c_261_p N_7_M11_d N_7_M12_d N_7_c_262_p N_7_M25_d N_7_c_263_p N_7_M26_s
+ N_7_c_218_n N_7_c_249_p N_7_c_219_n N_7_c_220_n N_7_c_248_p N_7_c_221_n
+ N_7_c_222_n N_7_c_258_p N_7_c_305_p N_7_c_253_p N_7_c_247_p N_7_c_240_p
+ N_7_c_233_p N_7_c_216_n N_7_c_236_p N_7_c_223_n N_7_c_224_n N_7_c_293_p
+ N_7_c_280_p N_7_c_289_p N_7_c_241_p N_7_c_267_p N_7_c_225_n N_7_c_246_p
+ N_7_c_260_p N_7_c_226_n N_7_c_244_p N_7_c_228_n N_7_c_229_n N_7_c_287_p
+ N_7_c_271_p VSS PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%7
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%RESET N_RESET_M6_g N_RESET_c_323_n N_RESET_M23_g
+ N_RESET_M13_g N_RESET_c_352_p N_RESET_M30_g N_RESET_c_310_n RESET
+ N_RESET_c_329_n N_RESET_c_311_n N_RESET_c_355_p N_RESET_c_332_n
+ N_RESET_c_312_n N_RESET_c_313_n N_RESET_c_314_n N_RESET_c_320_n
+ N_RESET_c_335_n N_RESET_c_336_n N_RESET_c_339_p N_RESET_c_315_n VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%RESET
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%9 N_9_M8_g N_9_c_367_n N_9_M25_g N_9_M4_s N_9_M3_d
+ N_9_c_412_p N_9_M20_d N_9_c_380_n N_9_M21_s N_9_c_388_n N_9_c_382_n
+ N_9_c_368_n N_9_c_389_n N_9_c_398_n N_9_c_370_n N_9_c_372_n N_9_c_385_n
+ N_9_c_418_p N_9_c_373_n N_9_c_374_n N_9_c_375_n N_9_c_376_n N_9_c_377_n
+ N_9_c_378_n VSS PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%9
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%SET N_SET_M7_g N_SET_M24_g N_SET_M9_g N_SET_M12_g
+ N_SET_c_429_n N_SET_M29_g SET N_SET_c_434_n N_SET_c_461_n VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%SET
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%11 N_11_M14_g N_11_c_521_n N_11_M31_g N_11_M16_g
+ N_11_c_557_p N_11_M32_g N_11_M11_s N_11_M10_d N_11_c_502_n N_11_M27_s
+ N_11_M26_d N_11_c_503_n N_11_c_505_n N_11_c_546_p N_11_c_493_n N_11_c_495_n
+ N_11_c_492_n N_11_c_524_n N_11_c_558_p N_11_c_534_p N_11_c_526_n N_11_c_559_p
+ N_11_c_500_n N_11_c_512_n N_11_c_514_n N_11_c_516_n N_11_c_517_n N_11_c_518_n
+ N_11_c_519_n VSS PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%11
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%12 N_12_c_564_n N_12_c_582_n N_12_c_583_n
+ N_12_c_586_n N_12_c_562_n N_12_M28_g N_12_M15_g N_12_c_591_n N_12_M14_s
+ N_12_M13_d N_12_c_569_n N_12_M31_d VSS PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%12
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%13 N_13_M4_d N_13_c_599_n N_13_M6_s N_13_M5_d
+ N_13_c_602_n N_13_c_603_n N_13_c_596_n N_13_c_605_n N_13_c_607_n N_13_c_598_n
+ VSS PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%13
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%14 N_14_M10_s N_14_M9_d N_14_c_613_n N_14_M15_d
+ N_14_c_615_n N_14_c_620_n N_14_c_621_n N_14_c_608_n N_14_c_629_n VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%14
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%QN N_QN_M16_d N_QN_M32_d QN N_QN_c_637_n VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%QN
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%16 N_16_M19_d N_16_M20_s N_16_c_638_n VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%16
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%17 N_17_M21_d N_17_M22_s N_17_c_647_n VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%17
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%18 N_18_M3_s N_18_M2_d VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%18
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%19 N_19_M23_s N_19_M22_d VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%19
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%20 N_20_M25_s N_20_M24_d VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%20
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%21 N_21_M28_s N_21_M27_d VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%21
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%22 N_22_M29_s N_22_M28_d VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%22
x_PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%23 N_23_M31_s N_23_M30_d VSS
+ PM_ASYNC_DFFHX1_ASAP7_75T_SRAM%23
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_23_n 3.57152e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 CLK N_4_c_24_n 0.00135805f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.144
cc_4 CLK N_4_c_25_n 2.75361e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.07
cc_5 CLK N_4_c_26_n 0.00135805f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.107
cc_6 N_CLK_c_6_p N_4_c_27_n 0.0014229f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2
cc_7 N_CLK_c_6_p N_4_c_28_n 2.75361e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2125
cc_8 CLK N_4_c_29_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_6_p N_4_c_30_n 5.03453e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_6_p N_4_c_31_n 0.00123168f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.153
cc_11 CLK N_4_c_32_n 4.37953e-19 $X=0.082 $Y=0.119 $X2=0.175 $Y2=0.153
cc_12 N_CLK_c_6_p N_4_c_32_n 0.00154146f $X=0.081 $Y=0.135 $X2=0.175 $Y2=0.153
cc_13 N_CLK_c_13_p N_4_c_34_n 0.0011431f $X=0.081 $Y=0.135 $X2=0.151 $Y2=0.135
cc_14 CLK N_4_c_35_n 0.00190651f $X=0.082 $Y=0.119 $X2=0.151 $Y2=0.135
cc_15 CLK N_6_c_127_n 6.37157e-19 $X=0.082 $Y=0.119 $X2=0 $Y2=0
cc_16 N_CLK_c_6_p N_6_c_128_n 6.45547e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.045
cc_17 N_CLK_c_6_p N_6_c_129_n 7.79176e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.2
cc_18 N_CLK_c_6_p N_6_c_130_n 3.83659e-19 $X=0.081 $Y=0.135 $X2=0.0505 $Y2=0.234
cc_19 CLK N_6_c_131_n 7.86679e-19 $X=0.082 $Y=0.119 $X2=0.838 $Y2=0.153
cc_20 CLK N_6_c_132_n 3.35174e-19 $X=0.082 $Y=0.119 $X2=0.838 $Y2=0.153
cc_21 N_CLK_c_6_p N_6_c_133_n 3.35174e-19 $X=0.081 $Y=0.135 $X2=0.735 $Y2=0.153
cc_22 N_4_M3_g N_D_M2_g 0.00341068f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_23 N_4_c_37_p N_D_c_108_n 0.00112574f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_4_c_38_p N_D_c_108_n 3.1268e-19 $X=0.364 $Y=0.153 $X2=0.081 $Y2=0.135
cc_25 N_4_c_34_n N_D_c_108_n 2.54877e-19 $X=0.151 $Y=0.135 $X2=0.081 $Y2=0.135
cc_26 N_4_c_40_p N_D_c_111_n 4.05496e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_27 N_4_c_41_p N_D_c_112_n 4.46721e-19 $X=0.263 $Y=0.153 $X2=0 $Y2=0
cc_28 N_4_c_38_p N_D_c_113_n 4.46721e-19 $X=0.364 $Y=0.153 $X2=0 $Y2=0
cc_29 N_4_c_41_p N_D_c_114_n 9.35374e-19 $X=0.263 $Y=0.153 $X2=0 $Y2=0
cc_30 N_4_c_40_p N_D_c_114_n 2.69506e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_31 N_4_M3_g N_6_M4_g 0.00355599f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_32 N_4_c_46_p N_6_M4_g 0.00360681f $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.054
cc_33 N_4_c_37_p N_6_c_136_n 9.95945e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_34 N_4_c_46_p N_6_c_136_n 0.00103912f $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.135
cc_35 N_4_M10_g N_6_M11_g 0.00360681f $X=0.837 $Y=0.054 $X2=0 $Y2=0
cc_36 N_4_c_50_p N_6_c_139_n 0.00149895f $X=0.837 $Y=0.111 $X2=0 $Y2=0
cc_37 N_4_c_35_n N_6_c_127_n 2.97444e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_32_n N_6_c_141_n 2.38327e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_35_n N_6_c_128_n 3.21026e-19 $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_41_p N_6_c_129_n 2.46239e-19 $X=0.263 $Y=0.153 $X2=0 $Y2=0
cc_41 N_4_c_32_n N_6_c_144_n 2.31165e-19 $X=0.175 $Y=0.153 $X2=0 $Y2=0
cc_42 N_4_c_56_p N_6_c_145_n 2.46239e-19 $X=0.4115 $Y=0.153 $X2=0 $Y2=0
cc_43 N_4_c_41_p N_6_c_130_n 0.0278758f $X=0.263 $Y=0.153 $X2=0 $Y2=0
cc_44 N_4_c_40_p N_6_c_130_n 4.50946e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_45 N_4_c_59_p N_6_c_130_n 2.98641e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_60_p N_6_c_149_n 0.0278758f $X=0.632 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_61_p N_6_c_149_n 3.05992e-19 $X=0.838 $Y=0.113 $X2=0 $Y2=0
cc_48 N_4_c_56_p N_6_c_151_n 5.90855e-19 $X=0.4115 $Y=0.153 $X2=0 $Y2=0
cc_49 N_4_c_60_p N_6_c_151_n 2.40893e-19 $X=0.632 $Y=0.153 $X2=0 $Y2=0
cc_50 N_4_c_40_p N_6_c_151_n 0.00211678f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_51 N_4_c_59_p N_6_c_151_n 0.00210743f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_52 N_4_c_66_p N_6_c_155_n 2.23575e-19 $X=0.838 $Y=0.153 $X2=0 $Y2=0
cc_53 N_4_c_61_p N_6_c_155_n 0.00298694f $X=0.838 $Y=0.113 $X2=0 $Y2=0
cc_54 N_4_c_41_p N_6_c_157_n 8.79704e-19 $X=0.263 $Y=0.153 $X2=0 $Y2=0
cc_55 N_4_c_35_n N_6_c_157_n 0.00528524f $X=0.151 $Y=0.135 $X2=0 $Y2=0
cc_56 N_4_c_46_p N_7_M5_g 2.62226e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.054
cc_57 N_4_c_71_p N_7_c_216_n 0.00105927f $X=0.735 $Y=0.153 $X2=0 $Y2=0
cc_58 N_4_c_60_p N_RESET_c_310_n 0.00106702f $X=0.632 $Y=0.153 $X2=0 $Y2=0
cc_59 N_4_c_71_p N_RESET_c_311_n 2.46239e-19 $X=0.735 $Y=0.153 $X2=0 $Y2=0
cc_60 N_4_c_71_p N_RESET_c_312_n 0.00878705f $X=0.735 $Y=0.153 $X2=0 $Y2=0
cc_61 N_4_c_66_p N_RESET_c_313_n 0.00878705f $X=0.838 $Y=0.153 $X2=0 $Y2=0
cc_62 N_4_c_61_p N_RESET_c_314_n 0.00105485f $X=0.838 $Y=0.113 $X2=0 $Y2=0
cc_63 N_4_c_71_p N_RESET_c_315_n 2.16564e-19 $X=0.735 $Y=0.153 $X2=0 $Y2=0
cc_64 N_4_M10_g N_9_M8_g 2.62226e-19 $X=0.837 $Y=0.054 $X2=0.081 $Y2=0.054
cc_65 N_4_c_50_p N_9_c_367_n 7.72364e-19 $X=0.837 $Y=0.111 $X2=0.081 $Y2=0.135
cc_66 N_4_c_46_p N_9_c_368_n 3.49806e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_67 N_4_c_59_p N_9_c_368_n 3.81288e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_68 N_4_c_60_p N_9_c_370_n 0.00119816f $X=0.632 $Y=0.153 $X2=0 $Y2=0
cc_69 N_4_c_59_p N_9_c_370_n 0.0024197f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_70 N_4_c_59_p N_9_c_372_n 0.00215948f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_71 N_4_c_56_p N_9_c_373_n 3.3297e-19 $X=0.4115 $Y=0.153 $X2=0 $Y2=0
cc_72 N_4_c_60_p N_9_c_374_n 3.14696e-19 $X=0.632 $Y=0.153 $X2=0 $Y2=0
cc_73 N_4_c_71_p N_9_c_375_n 0.00324726f $X=0.735 $Y=0.153 $X2=0 $Y2=0
cc_74 N_4_c_71_p N_9_c_376_n 2.1652e-19 $X=0.735 $Y=0.153 $X2=0 $Y2=0
cc_75 N_4_c_56_p N_9_c_377_n 0.00324726f $X=0.4115 $Y=0.153 $X2=0 $Y2=0
cc_76 N_4_c_60_p N_9_c_378_n 0.00324726f $X=0.632 $Y=0.153 $X2=0 $Y2=0
cc_77 N_4_M10_g N_SET_M9_g 0.00353416f $X=0.837 $Y=0.054 $X2=0 $Y2=0
cc_78 N_4_M10_g N_SET_c_429_n 0.0026337f $X=0.837 $Y=0.054 $X2=0 $Y2=0
cc_79 N_4_c_50_p N_SET_c_429_n 0.0017762f $X=0.837 $Y=0.111 $X2=0 $Y2=0
cc_80 N_4_c_61_p N_SET_c_429_n 0.0025321f $X=0.838 $Y=0.113 $X2=0 $Y2=0
cc_81 N_4_c_50_p SET 2.54502e-19 $X=0.837 $Y=0.111 $X2=0 $Y2=0
cc_82 N_4_c_61_p SET 0.00283263f $X=0.838 $Y=0.113 $X2=0 $Y2=0
cc_83 N_4_c_66_p N_SET_c_434_n 5.90485e-19 $X=0.838 $Y=0.153 $X2=0 $Y2=0
cc_84 N_4_c_66_p N_11_c_492_n 6.36189e-19 $X=0.838 $Y=0.153 $X2=0 $Y2=0
cc_85 N_4_M10_g N_12_c_562_n 3.04066e-19 $X=0.837 $Y=0.054 $X2=0.081 $Y2=0.135
cc_86 N_4_c_46_p N_13_c_596_n 3.75215e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_87 N_4_c_59_p N_13_c_596_n 2.37912e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_88 N_4_c_66_p N_14_c_608_n 2.43239e-19 $X=0.838 $Y=0.153 $X2=0 $Y2=0
cc_89 N_4_M3_g N_16_c_638_n 0.00442838f $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_90 N_4_c_37_p N_16_c_638_n 0.00393643f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_91 N_4_c_38_p N_16_c_638_n 4.52862e-19 $X=0.364 $Y=0.153 $X2=0 $Y2=0
cc_92 N_4_c_40_p N_16_c_638_n 0.0015121f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_93 N_D_M2_g N_6_M4_g 2.92202e-19 $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_94 D N_6_c_160_n 0.00153722f $X=0.244 $Y=0.082 $X2=0 $Y2=0
cc_95 N_D_c_114_n N_6_c_161_n 0.00153722f $X=0.243 $Y=0.135 $X2=0.018 $Y2=0.225
cc_96 N_D_c_114_n N_6_c_129_n 0.00153722f $X=0.243 $Y=0.135 $X2=0.018 $Y2=0.2
cc_97 N_D_c_108_n N_6_c_130_n 2.11873e-19 $X=0.297 $Y=0.135 $X2=0.0505 $Y2=0.234
cc_98 N_D_c_114_n N_6_c_130_n 0.00134413f $X=0.243 $Y=0.135 $X2=0.0505 $Y2=0.234
cc_99 D N_6_c_131_n 0.00153722f $X=0.244 $Y=0.082 $X2=0.838 $Y2=0.153
cc_100 D N_6_c_132_n 0.00153722f $X=0.244 $Y=0.082 $X2=0.838 $Y2=0.153
cc_101 N_D_c_124_p N_6_c_157_n 0.00153722f $X=0.243 $Y=0.123 $X2=0.632 $Y2=0.153
cc_102 N_D_c_125_p N_6_c_133_n 0.00153722f $X=0.243 $Y=0.126 $X2=0.735 $Y2=0.153
cc_103 D N_9_c_377_n 2.22013e-19 $X=0.244 $Y=0.082 $X2=0.0505 $Y2=0.036
cc_104 N_6_c_130_n N_7_c_217_n 4.23437e-19 $X=0.741 $Y=0.189 $X2=0.081 $Y2=0.135
cc_105 N_6_c_149_n N_7_c_218_n 6.84883e-19 $X=0.852 $Y=0.189 $X2=0 $Y2=0
cc_106 N_6_c_130_n N_7_c_219_n 6.87626e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_107 N_6_c_130_n N_7_c_220_n 3.92349e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_108 N_6_c_130_n N_7_c_221_n 4.18502e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_109 N_6_c_130_n N_7_c_222_n 9.37967e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_110 N_6_c_130_n N_7_c_223_n 8.1356e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_111 N_6_c_130_n N_7_c_224_n 3.92349e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_112 N_6_c_149_n N_7_c_225_n 2.46239e-19 $X=0.852 $Y=0.189 $X2=0 $Y2=0
cc_113 N_6_c_178_p N_7_c_226_n 2.93332e-19 $X=0.891 $Y=0.189 $X2=0 $Y2=0
cc_114 N_6_c_149_n N_7_c_226_n 0.0140767f $X=0.852 $Y=0.189 $X2=0 $Y2=0
cc_115 N_6_c_130_n N_7_c_228_n 7.24284e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_116 N_6_c_149_n N_7_c_229_n 3.16423e-19 $X=0.852 $Y=0.189 $X2=0 $Y2=0
cc_117 N_6_c_130_n RESET 0.0012955f $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_118 N_6_c_130_n N_RESET_c_312_n 0.00100574f $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_119 N_6_c_149_n N_RESET_c_313_n 0.00100574f $X=0.852 $Y=0.189 $X2=0 $Y2=0
cc_120 N_6_c_185_p N_RESET_c_314_n 0.00100574f $X=0.891 $Y=0.189 $X2=0 $Y2=0
cc_121 N_6_c_155_n N_RESET_c_320_n 8.58654e-19 $X=0.891 $Y=0.111 $X2=0 $Y2=0
cc_122 N_6_c_130_n N_9_c_380_n 2.04929e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_123 N_6_c_151_n N_9_c_380_n 0.00115602f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_124 N_6_c_130_n N_9_c_382_n 0.00110489f $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_125 N_6_c_190_p N_9_c_370_n 4.11789e-19 $X=0.405 $Y=0.178 $X2=0 $Y2=0
cc_126 N_6_c_145_n N_9_c_372_n 4.11789e-19 $X=0.405 $Y=0.189 $X2=0 $Y2=0
cc_127 N_6_c_130_n N_9_c_385_n 0.00109006f $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_128 N_6_c_130_n N_9_c_377_n 9.78803e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_129 N_6_M11_g N_SET_M9_g 2.98134e-19 $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_130 N_6_M11_g N_SET_M12_g 2.92202e-19 $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_131 N_6_M11_g N_SET_c_429_n 0.0016486f $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_132 N_6_c_139_n N_SET_c_429_n 0.00204145f $X=0.891 $Y=0.111 $X2=0 $Y2=0
cc_133 N_6_c_130_n N_SET_c_429_n 4.15894e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_134 N_6_c_149_n N_SET_c_429_n 3.98282e-19 $X=0.852 $Y=0.189 $X2=0 $Y2=0
cc_135 N_6_c_155_n N_SET_c_429_n 0.00205489f $X=0.891 $Y=0.111 $X2=0 $Y2=0
cc_136 N_6_c_201_p N_SET_c_429_n 4.75629e-19 $X=0.891 $Y=0.173 $X2=0 $Y2=0
cc_137 N_6_M11_g N_11_c_493_n 3.09683e-19 $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_138 N_6_c_155_n N_11_c_493_n 5.25723e-19 $X=0.891 $Y=0.111 $X2=0 $Y2=0
cc_139 N_6_c_139_n N_11_c_495_n 4.82891e-19 $X=0.891 $Y=0.111 $X2=0 $Y2=0
cc_140 N_6_c_185_p N_11_c_495_n 3.64939e-19 $X=0.891 $Y=0.189 $X2=0 $Y2=0
cc_141 N_6_c_178_p N_11_c_495_n 2.60223e-19 $X=0.891 $Y=0.189 $X2=0 $Y2=0
cc_142 N_6_c_155_n N_11_c_495_n 0.00914084f $X=0.891 $Y=0.111 $X2=0 $Y2=0
cc_143 N_6_c_155_n N_11_c_492_n 2.7717e-19 $X=0.891 $Y=0.111 $X2=0 $Y2=0
cc_144 N_6_M11_g N_11_c_500_n 0.00206017f $X=0.891 $Y=0.0405 $X2=0 $Y2=0
cc_145 N_6_c_178_p N_11_c_500_n 0.00148428f $X=0.891 $Y=0.189 $X2=0 $Y2=0
cc_146 N_6_M11_g N_12_c_562_n 0.00355599f $X=0.891 $Y=0.0405 $X2=0.081 $Y2=0.135
cc_147 N_6_c_130_n N_16_c_638_n 9.26664e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_148 N_6_c_151_n N_16_c_638_n 0.00115662f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_149 N_6_c_130_n N_17_c_647_n 9.27655e-19 $X=0.741 $Y=0.189 $X2=0 $Y2=0
cc_150 N_7_M5_g N_RESET_M6_g 0.00328721f $X=0.567 $Y=0.054 $X2=0.135 $Y2=0.054
cc_151 N_7_c_222_n N_RESET_M6_g 2.50234e-19 $X=0.668 $Y=0.225 $X2=0.135
+ $Y2=0.054
cc_152 N_7_c_216_n N_RESET_c_323_n 2.70122e-19 $X=0.702 $Y=0.173 $X2=0.135
+ $Y2=0.135
cc_153 N_7_c_233_p N_RESET_c_310_n 4.04895e-19 $X=0.702 $Y=0.133 $X2=0 $Y2=0
cc_154 N_7_c_217_n RESET 3.90177e-19 $X=0.567 $Y=0.18 $X2=0 $Y2=0
cc_155 N_7_c_222_n RESET 0.00500136f $X=0.668 $Y=0.225 $X2=0 $Y2=0
cc_156 N_7_c_236_p RESET 4.04895e-19 $X=0.702 $Y=0.18 $X2=0 $Y2=0
cc_157 N_7_c_223_n RESET 0.00109903f $X=0.702 $Y=0.198 $X2=0 $Y2=0
cc_158 N_7_c_219_n N_RESET_c_329_n 0.00146693f $X=0.567 $Y=0.18 $X2=0.837
+ $Y2=0.111
cc_159 N_7_c_216_n N_RESET_c_329_n 4.04895e-19 $X=0.702 $Y=0.173 $X2=0.837
+ $Y2=0.111
cc_160 N_7_c_240_p N_RESET_c_311_n 0.00101662f $X=0.702 $Y=0.126 $X2=0 $Y2=0
cc_161 N_7_c_241_p N_RESET_c_332_n 0.00156236f $X=0.972 $Y=0.168 $X2=0.056
+ $Y2=0.216
cc_162 N_7_c_240_p N_RESET_c_312_n 5.07186e-19 $X=0.702 $Y=0.126 $X2=0 $Y2=0
cc_163 N_7_c_226_n N_RESET_c_320_n 2.31241e-19 $X=0.905 $Y=0.225 $X2=0.018
+ $Y2=0.045
cc_164 N_7_c_244_p N_RESET_c_335_n 2.31241e-19 $X=0.913 $Y=0.225 $X2=0.018
+ $Y2=0.144
cc_165 N_7_c_241_p N_RESET_c_336_n 0.00116776f $X=0.972 $Y=0.168 $X2=0.018
+ $Y2=0.07
cc_166 N_7_c_246_p N_RESET_c_336_n 2.31241e-19 $X=0.994 $Y=0.225 $X2=0.018
+ $Y2=0.07
cc_167 N_7_c_247_p N_9_c_367_n 5.43243e-19 $X=0.702 $Y=0.108 $X2=0.135 $Y2=0.135
cc_168 N_7_c_248_p N_9_c_388_n 5.07262e-19 $X=0.576 $Y=0.225 $X2=0.837
+ $Y2=0.2295
cc_169 N_7_c_249_p N_9_c_389_n 5.07262e-19 $X=0.567 $Y=0.216 $X2=0.071 $Y2=0.216
cc_170 N_7_c_219_n N_9_c_372_n 5.07262e-19 $X=0.567 $Y=0.18 $X2=0.018 $Y2=0.045
cc_171 N_7_c_217_n N_9_c_385_n 2.12288e-19 $X=0.567 $Y=0.18 $X2=0.018 $Y2=0.144
cc_172 N_7_c_220_n N_9_c_385_n 5.07262e-19 $X=0.567 $Y=0.207 $X2=0.018 $Y2=0.144
cc_173 N_7_c_253_p N_9_c_375_n 0.00108015f $X=0.702 $Y=0.072 $X2=0.054 $Y2=0.036
cc_174 N_7_c_253_p N_9_c_376_n 0.00438159f $X=0.702 $Y=0.072 $X2=0.047 $Y2=0.036
cc_175 N_7_c_240_p N_9_c_376_n 0.00193057f $X=0.702 $Y=0.126 $X2=0.047 $Y2=0.036
cc_176 N_7_c_229_n N_9_c_376_n 2.06687e-19 $X=0.747 $Y=0.225 $X2=0.047 $Y2=0.036
cc_177 N_7_M5_g N_SET_M7_g 2.20386e-19 $X=0.567 $Y=0.054 $X2=0.135 $Y2=0.054
cc_178 N_7_c_258_p N_SET_M7_g 3.55898e-19 $X=0.6805 $Y=0.225 $X2=0.135 $Y2=0.054
cc_179 N_7_c_218_n N_SET_M9_g 0.00370848f $X=0.812 $Y=0.2295 $X2=0.351
+ $Y2=0.0675
cc_180 N_7_c_260_p N_SET_M12_g 8.17918e-19 $X=0.994 $Y=0.225 $X2=0.459 $Y2=0.135
cc_181 N_7_c_261_p N_SET_c_429_n 6.2404e-19 $X=0.702 $Y=0.0405 $X2=0.459
+ $Y2=0.2295
cc_182 N_7_c_262_p N_SET_c_429_n 6.53599e-19 $X=0.974 $Y=0.0405 $X2=0.459
+ $Y2=0.2295
cc_183 N_7_c_263_p N_SET_c_429_n 2.8383e-19 $X=0.754 $Y=0.216 $X2=0.459
+ $Y2=0.2295
cc_184 N_7_c_218_n N_SET_c_429_n 0.00555074f $X=0.812 $Y=0.2295 $X2=0.459
+ $Y2=0.2295
cc_185 N_7_c_216_n N_SET_c_429_n 0.0461621f $X=0.702 $Y=0.173 $X2=0.459
+ $Y2=0.2295
cc_186 N_7_c_241_p N_SET_c_429_n 0.0020951f $X=0.972 $Y=0.168 $X2=0.459
+ $Y2=0.2295
cc_187 N_7_c_267_p N_SET_c_429_n 9.77809e-19 $X=0.972 $Y=0.192 $X2=0.459
+ $Y2=0.2295
cc_188 N_7_c_246_p N_SET_c_429_n 2.30766e-19 $X=0.994 $Y=0.225 $X2=0.459
+ $Y2=0.2295
cc_189 N_7_c_228_n N_SET_c_429_n 7.70908e-19 $X=0.729 $Y=0.225 $X2=0.459
+ $Y2=0.2295
cc_190 N_7_c_229_n N_SET_c_429_n 3.03524e-19 $X=0.747 $Y=0.225 $X2=0.459
+ $Y2=0.2295
cc_191 N_7_c_271_p N_SET_c_429_n 2.16231e-19 $X=0.9875 $Y=0.225 $X2=0.459
+ $Y2=0.2295
cc_192 N_7_c_218_n N_SET_c_434_n 5.03908e-19 $X=0.812 $Y=0.2295 $X2=0 $Y2=0
cc_193 N_7_c_233_p N_SET_c_434_n 3.35238e-19 $X=0.702 $Y=0.133 $X2=0 $Y2=0
cc_194 N_7_c_216_n N_SET_c_434_n 3.35238e-19 $X=0.702 $Y=0.173 $X2=0 $Y2=0
cc_195 N_7_c_247_p N_SET_c_461_n 3.35238e-19 $X=0.702 $Y=0.108 $X2=0.018
+ $Y2=0.07
cc_196 N_7_c_262_p N_11_c_502_n 0.00194094f $X=0.974 $Y=0.0405 $X2=0.837
+ $Y2=0.054
cc_197 N_7_c_218_n N_11_c_503_n 0.00376276f $X=0.812 $Y=0.2295 $X2=0.837
+ $Y2=0.2295
cc_198 N_7_c_226_n N_11_c_503_n 5.51168e-19 $X=0.905 $Y=0.225 $X2=0.837
+ $Y2=0.2295
cc_199 N_7_c_262_p N_11_c_505_n 0.00218053f $X=0.974 $Y=0.0405 $X2=0.837
+ $Y2=0.2295
cc_200 N_7_c_280_p N_11_c_505_n 0.00171412f $X=0.972 $Y=0.045 $X2=0.837
+ $Y2=0.2295
cc_201 N_7_c_241_p N_11_c_492_n 0.00111708f $X=0.972 $Y=0.168 $X2=0.018
+ $Y2=0.107
cc_202 N_7_c_246_p N_11_c_492_n 0.00310274f $X=0.994 $Y=0.225 $X2=0.018
+ $Y2=0.107
cc_203 N_7_c_271_p N_11_c_492_n 2.49288e-19 $X=0.9875 $Y=0.225 $X2=0.018
+ $Y2=0.107
cc_204 N_7_c_267_p N_11_c_500_n 2.73999e-19 $X=0.972 $Y=0.192 $X2=0.351
+ $Y2=0.153
cc_205 N_7_c_226_n N_11_c_500_n 3.68491e-19 $X=0.905 $Y=0.225 $X2=0.351
+ $Y2=0.153
cc_206 N_7_c_246_p N_11_c_512_n 3.11447e-19 $X=0.994 $Y=0.225 $X2=0.351
+ $Y2=0.153
cc_207 N_7_c_287_p N_11_c_512_n 0.00171412f $X=0.981 $Y=0.225 $X2=0.351
+ $Y2=0.153
cc_208 N_7_c_262_p N_11_c_514_n 3.35225e-19 $X=0.974 $Y=0.0405 $X2=0.263
+ $Y2=0.153
cc_209 N_7_c_289_p N_11_c_514_n 0.00171412f $X=0.972 $Y=0.103 $X2=0.263
+ $Y2=0.153
cc_210 N_7_c_262_p N_11_c_516_n 0.0385594f $X=0.974 $Y=0.0405 $X2=0.459
+ $Y2=0.153
cc_211 N_7_c_241_p N_11_c_517_n 0.00171412f $X=0.972 $Y=0.168 $X2=0.459
+ $Y2=0.153
cc_212 N_7_c_267_p N_11_c_518_n 0.00171412f $X=0.972 $Y=0.192 $X2=0.364
+ $Y2=0.153
cc_213 N_7_c_293_p N_11_c_519_n 0.00171412f $X=0.972 $Y=0.216 $X2=0.4115
+ $Y2=0.153
cc_214 N_7_M12_d N_12_c_564_n 2.25873e-19 $X=0.989 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_215 N_7_c_262_p N_12_c_564_n 0.00154164f $X=0.974 $Y=0.0405 $X2=0.135
+ $Y2=0.054
cc_216 N_7_c_289_p N_12_c_564_n 0.00228569f $X=0.972 $Y=0.103 $X2=0.135
+ $Y2=0.054
cc_217 N_7_c_241_p N_12_c_564_n 0.0437738f $X=0.972 $Y=0.168 $X2=0.135 $Y2=0.054
cc_218 N_7_c_262_p N_12_c_562_n 0.00268304f $X=0.974 $Y=0.0405 $X2=0.459
+ $Y2=0.135
cc_219 N_7_c_289_p N_12_c_569_n 6.51818e-19 $X=0.972 $Y=0.103 $X2=0.056
+ $Y2=0.216
cc_220 N_7_M5_g N_13_c_598_n 4.71295e-19 $X=0.567 $Y=0.054 $X2=0.837 $Y2=0.111
cc_221 N_7_c_262_p N_14_c_608_n 5.31664e-19 $X=0.974 $Y=0.0405 $X2=0.459
+ $Y2=0.2295
cc_222 N_7_c_280_p N_14_c_608_n 7.44496e-19 $X=0.972 $Y=0.045 $X2=0.459
+ $Y2=0.2295
cc_223 N_7_c_289_p N_14_c_608_n 3.13568e-19 $X=0.972 $Y=0.103 $X2=0.459
+ $Y2=0.2295
cc_224 N_7_c_221_n N_19_M23_s 3.16072e-19 $X=0.608 $Y=0.225 $X2=0.135 $Y2=0.054
cc_225 N_7_c_305_p N_20_M25_s 2.40538e-19 $X=0.702 $Y=0.216 $X2=0.135 $Y2=0.054
cc_226 N_7_c_223_n N_20_M25_s 4.55529e-19 $X=0.702 $Y=0.198 $X2=0.135 $Y2=0.054
cc_227 N_7_c_293_p N_22_M29_s 2.06543e-19 $X=0.972 $Y=0.216 $X2=0.135 $Y2=0.054
cc_228 N_7_c_267_p N_22_M29_s 2.55017e-19 $X=0.972 $Y=0.192 $X2=0.135 $Y2=0.054
cc_229 N_7_c_287_p N_22_M29_s 5.91249e-19 $X=0.981 $Y=0.225 $X2=0.135 $Y2=0.054
cc_230 N_RESET_M6_g N_9_M8_g 2.20386e-19 $X=0.621 $Y=0.054 $X2=0.135 $Y2=0.054
cc_231 N_RESET_c_339_p N_9_c_398_n 3.87136e-19 $X=0.63 $Y=0.117 $X2=0.056
+ $Y2=0.216
cc_232 N_RESET_c_310_n N_9_c_370_n 3.87136e-19 $X=0.621 $Y=0.159 $X2=0 $Y2=0
cc_233 N_RESET_c_312_n N_9_c_376_n 8.88087e-19 $X=0.752 $Y=0.117 $X2=0.047
+ $Y2=0.036
cc_234 N_RESET_c_311_n N_9_c_378_n 2.46239e-19 $X=0.646 $Y=0.117 $X2=0 $Y2=0
cc_235 N_RESET_c_312_n N_9_c_378_n 0.010102f $X=0.752 $Y=0.117 $X2=0 $Y2=0
cc_236 N_RESET_c_315_n N_9_c_378_n 2.61262e-19 $X=0.638 $Y=0.117 $X2=0 $Y2=0
cc_237 N_RESET_M6_g N_SET_M7_g 0.00268443f $X=0.621 $Y=0.054 $X2=0.135 $Y2=0.054
cc_238 N_RESET_M13_g N_SET_M12_g 0.00268443f $X=1.053 $Y=0.0405 $X2=0.459
+ $Y2=0.135
cc_239 N_RESET_c_313_n N_SET_c_429_n 3.16544e-19 $X=0.778 $Y=0.117 $X2=0.459
+ $Y2=0.2295
cc_240 N_RESET_c_320_n N_SET_c_429_n 2.74499e-19 $X=0.905 $Y=0.117 $X2=0.459
+ $Y2=0.2295
cc_241 N_RESET_c_313_n SET 2.15567e-19 $X=0.778 $Y=0.117 $X2=0.071 $Y2=0.216
cc_242 N_RESET_c_314_n SET 7.58196e-19 $X=0.852 $Y=0.117 $X2=0.071 $Y2=0.216
cc_243 N_RESET_M13_g N_11_M14_g 0.00328721f $X=1.053 $Y=0.0405 $X2=0.135
+ $Y2=0.054
cc_244 N_RESET_c_352_p N_11_c_521_n 0.00112281f $X=1.053 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_245 N_RESET_c_336_n N_11_c_495_n 0.00122107f $X=0.983 $Y=0.117 $X2=0.056
+ $Y2=0.216
cc_246 N_RESET_c_336_n N_11_c_492_n 0.00636555f $X=0.983 $Y=0.117 $X2=0.018
+ $Y2=0.107
cc_247 N_RESET_c_355_p N_11_c_524_n 0.00636555f $X=1.053 $Y=0.117 $X2=0.018
+ $Y2=0.162
cc_248 N_RESET_c_332_n N_11_c_524_n 0.00143908f $X=1.053 $Y=0.117 $X2=0.018
+ $Y2=0.162
cc_249 N_RESET_c_355_p N_11_c_526_n 3.52128e-19 $X=1.053 $Y=0.117 $X2=0.0505
+ $Y2=0.036
cc_250 N_RESET_c_332_n N_11_c_526_n 0.00325783f $X=1.053 $Y=0.117 $X2=0.0505
+ $Y2=0.036
cc_251 N_RESET_M13_g N_12_c_564_n 0.00243042f $X=1.053 $Y=0.0405 $X2=0.135
+ $Y2=0.054
cc_252 N_RESET_c_352_p N_12_c_564_n 0.00201708f $X=1.053 $Y=0.135 $X2=0.135
+ $Y2=0.054
cc_253 N_RESET_c_355_p N_12_c_564_n 5.13068e-19 $X=1.053 $Y=0.117 $X2=0.135
+ $Y2=0.054
cc_254 N_RESET_c_332_n N_12_c_564_n 0.00148371f $X=1.053 $Y=0.117 $X2=0.135
+ $Y2=0.054
cc_255 N_RESET_M13_g N_12_c_562_n 2.20386e-19 $X=1.053 $Y=0.0405 $X2=0.459
+ $Y2=0.135
cc_256 N_RESET_M13_g N_12_M15_g 2.56294e-19 $X=1.053 $Y=0.0405 $X2=0.837
+ $Y2=0.054
cc_257 N_RESET_c_314_n N_14_c_608_n 0.00935401f $X=0.852 $Y=0.117 $X2=0.459
+ $Y2=0.2295
cc_258 N_9_M8_g N_SET_M7_g 0.00328721f $X=0.729 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_259 N_9_M8_g N_SET_M9_g 0.00312021f $X=0.729 $Y=0.0405 $X2=0.351 $Y2=0.0675
cc_260 N_9_M8_g N_SET_c_429_n 0.00283288f $X=0.729 $Y=0.0405 $X2=0.459
+ $Y2=0.2295
cc_261 N_9_c_367_n N_SET_c_429_n 0.00197192f $X=0.729 $Y=0.11 $X2=0.459
+ $Y2=0.2295
cc_262 N_9_c_376_n N_SET_c_429_n 4.17919e-19 $X=0.738 $Y=0.081 $X2=0.459
+ $Y2=0.2295
cc_263 N_9_c_367_n SET 3.68575e-19 $X=0.729 $Y=0.11 $X2=0.071 $Y2=0.216
cc_264 N_9_c_375_n SET 2.90481e-19 $X=0.738 $Y=0.081 $X2=0.071 $Y2=0.216
cc_265 N_9_c_376_n SET 0.00399229f $X=0.738 $Y=0.081 $X2=0.071 $Y2=0.216
cc_266 N_9_c_412_p N_13_c_599_n 0.00266305f $X=0.378 $Y=0.0675 $X2=0.135
+ $Y2=0.135
cc_267 N_9_c_380_n N_13_c_599_n 9.24647e-19 $X=0.432 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_268 N_9_c_377_n N_13_c_599_n 3.58627e-19 $X=0.632 $Y=0.081 $X2=0.135
+ $Y2=0.135
cc_269 N_9_c_377_n N_13_c_602_n 2.88367e-19 $X=0.632 $Y=0.081 $X2=0.351
+ $Y2=0.0675
cc_270 N_9_c_412_p N_13_c_603_n 5.11172e-19 $X=0.378 $Y=0.0675 $X2=0.351
+ $Y2=0.135
cc_271 N_9_c_377_n N_13_c_603_n 0.00126867f $X=0.632 $Y=0.081 $X2=0.351
+ $Y2=0.135
cc_272 N_9_c_418_p N_13_c_605_n 0.00370107f $X=0.504 $Y=0.081 $X2=0 $Y2=0
cc_273 N_9_c_377_n N_13_c_605_n 8.13509e-19 $X=0.632 $Y=0.081 $X2=0 $Y2=0
cc_274 N_9_c_377_n N_13_c_607_n 0.00106309f $X=0.632 $Y=0.081 $X2=0.837
+ $Y2=0.111
cc_275 N_9_c_412_p N_16_c_638_n 0.00137891f $X=0.378 $Y=0.0675 $X2=0.351
+ $Y2=0.0675
cc_276 N_9_c_380_n N_16_c_638_n 0.00376466f $X=0.432 $Y=0.2025 $X2=0.351
+ $Y2=0.0675
cc_277 N_9_c_382_n N_16_c_638_n 5.4984e-19 $X=0.45 $Y=0.234 $X2=0.351 $Y2=0.0675
cc_278 N_9_c_380_n N_17_c_647_n 0.00182426f $X=0.432 $Y=0.2025 $X2=0.351
+ $Y2=0.0675
cc_279 N_9_c_388_n N_17_c_647_n 0.00241571f $X=0.486 $Y=0.234 $X2=0.351
+ $Y2=0.0675
cc_280 N_9_c_389_n N_17_c_647_n 0.0417411f $X=0.495 $Y=0.225 $X2=0.351
+ $Y2=0.0675
cc_281 N_9_c_374_n N_17_c_647_n 3.16297e-19 $X=0.521 $Y=0.081 $X2=0.351
+ $Y2=0.0675
cc_282 N_SET_M12_g N_11_M14_g 2.20386e-19 $X=0.999 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_283 N_SET_c_429_n N_11_c_502_n 7.2973e-19 $X=0.999 $Y=0.159 $X2=0.837
+ $Y2=0.054
cc_284 N_SET_c_429_n N_11_c_503_n 0.00691652f $X=0.999 $Y=0.159 $X2=0.837
+ $Y2=0.2295
cc_285 N_SET_c_429_n N_11_c_495_n 0.0142846f $X=0.999 $Y=0.159 $X2=0.056
+ $Y2=0.216
cc_286 SET N_11_c_518_n 2.76553e-19 $X=0.782 $Y=0.132 $X2=0.364 $Y2=0.153
cc_287 N_SET_M12_g N_12_c_564_n 0.00274254f $X=0.999 $Y=0.0405 $X2=0.135
+ $Y2=0.054
cc_288 N_SET_c_429_n N_12_c_564_n 0.00133164f $X=0.999 $Y=0.159 $X2=0.135
+ $Y2=0.054
cc_289 N_SET_M12_g N_12_c_562_n 0.00341068f $X=0.999 $Y=0.0405 $X2=0.459
+ $Y2=0.135
cc_290 N_SET_c_429_n N_12_c_562_n 0.00251799f $X=0.999 $Y=0.159 $X2=0.459
+ $Y2=0.135
cc_291 N_SET_c_429_n N_14_c_613_n 8.13857e-19 $X=0.999 $Y=0.159 $X2=0.135
+ $Y2=0.135
cc_292 SET N_14_c_613_n 0.0313782f $X=0.782 $Y=0.132 $X2=0.135 $Y2=0.135
cc_293 N_SET_M9_g N_14_c_615_n 5.29542e-19 $X=0.783 $Y=0.054 $X2=0.351 $Y2=0.135
cc_294 SET N_14_c_615_n 0.00374033f $X=0.782 $Y=0.132 $X2=0.351 $Y2=0.135
cc_295 SET N_14_c_608_n 2.18952e-19 $X=0.782 $Y=0.132 $X2=0.459 $Y2=0.2295
cc_296 N_SET_c_429_n N_20_M25_s 0.00109397f $X=0.999 $Y=0.159 $X2=0.135
+ $Y2=0.054
cc_297 N_SET_c_429_n N_22_M29_s 0.00113446f $X=0.999 $Y=0.159 $X2=0.135
+ $Y2=0.054
cc_298 N_11_c_524_n N_12_c_564_n 3.52391e-19 $X=1.067 $Y=0.153 $X2=0.135
+ $Y2=0.054
cc_299 N_11_c_534_p N_12_c_564_n 4.54225e-19 $X=1.198 $Y=0.153 $X2=0.135
+ $Y2=0.054
cc_300 N_11_c_495_n N_12_c_582_n 2.50343e-19 $X=0.927 $Y=0.153 $X2=0 $Y2=0
cc_301 N_11_M14_g N_12_c_583_n 0.00243042f $X=1.107 $Y=0.0405 $X2=0.135
+ $Y2=0.135
cc_302 N_11_c_521_n N_12_c_583_n 0.00201708f $X=1.107 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_303 N_11_c_526_n N_12_c_583_n 0.0015034f $X=1.107 $Y=0.135 $X2=0.135
+ $Y2=0.135
cc_304 N_11_c_534_p N_12_c_586_n 0.00106459f $X=1.198 $Y=0.153 $X2=0.351
+ $Y2=0.0675
cc_305 N_11_c_526_n N_12_c_586_n 0.00102337f $X=1.107 $Y=0.135 $X2=0.351
+ $Y2=0.0675
cc_306 N_11_c_495_n N_12_c_562_n 6.34649e-19 $X=0.927 $Y=0.153 $X2=0.459
+ $Y2=0.135
cc_307 N_11_c_500_n N_12_c_562_n 9.73967e-19 $X=0.927 $Y=0.201 $X2=0.459
+ $Y2=0.135
cc_308 N_11_M14_g N_12_M15_g 0.00312021f $X=1.107 $Y=0.0405 $X2=0.837 $Y2=0.054
cc_309 N_11_c_534_p N_12_c_591_n 3.19267e-19 $X=1.198 $Y=0.153 $X2=0.837
+ $Y2=0.111
cc_310 N_11_c_502_n N_14_c_613_n 0.00276538f $X=0.864 $Y=0.054 $X2=0.135
+ $Y2=0.135
cc_311 N_11_c_546_p N_14_c_615_n 3.34076e-19 $X=0.882 $Y=0.039 $X2=0.351
+ $Y2=0.135
cc_312 N_11_c_534_p N_14_c_620_n 0.0011481f $X=1.198 $Y=0.153 $X2=0.459
+ $Y2=0.135
cc_313 N_11_c_534_p N_14_c_621_n 2.50936e-19 $X=1.198 $Y=0.153 $X2=0 $Y2=0
cc_314 N_11_c_502_n N_14_c_608_n 2.30142e-19 $X=0.864 $Y=0.054 $X2=0.459
+ $Y2=0.2295
cc_315 N_11_c_505_n N_14_c_608_n 0.00115993f $X=0.918 $Y=0.039 $X2=0.459
+ $Y2=0.2295
cc_316 N_11_c_546_p N_14_c_608_n 9.26825e-19 $X=0.882 $Y=0.039 $X2=0.459
+ $Y2=0.2295
cc_317 N_11_c_493_n N_14_c_608_n 4.78218e-19 $X=0.9 $Y=0.039 $X2=0.459
+ $Y2=0.2295
cc_318 N_11_c_492_n N_14_c_608_n 0.0011481f $X=1.008 $Y=0.153 $X2=0.459
+ $Y2=0.2295
cc_319 N_11_c_514_n N_14_c_608_n 2.15425e-19 $X=0.927 $Y=0.054 $X2=0.459
+ $Y2=0.2295
cc_320 N_11_c_516_n N_14_c_608_n 3.22466e-19 $X=0.927 $Y=0.058 $X2=0.459
+ $Y2=0.2295
cc_321 N_11_c_524_n N_14_c_629_n 0.0011481f $X=1.067 $Y=0.153 $X2=0.459
+ $Y2=0.2295
cc_322 N_11_c_557_p QN 3.33689e-19 $X=1.323 $Y=0.135 $X2=0 $Y2=0
cc_323 N_11_c_558_p QN 2.3227e-19 $X=1.323 $Y=0.153 $X2=0 $Y2=0
cc_324 N_11_c_559_p QN 0.00322962f $X=1.323 $Y=0.135 $X2=0 $Y2=0
cc_325 N_11_c_559_p N_QN_c_637_n 5.35809e-19 $X=1.323 $Y=0.135 $X2=0.837
+ $Y2=0.054
cc_326 N_11_c_500_n N_21_M28_s 0.00134416f $X=0.927 $Y=0.201 $X2=0.135 $Y2=0.054
cc_327 N_12_M15_g N_14_c_621_n 3.68583e-19 $X=1.161 $Y=0.0405 $X2=0 $Y2=0
cc_328 N_12_c_564_n N_14_c_608_n 7.14489e-19 $X=1.068 $Y=0.096 $X2=0.459
+ $Y2=0.2295
cc_329 N_12_c_583_n N_14_c_629_n 4.31546e-19 $X=1.146 $Y=0.096 $X2=0.459
+ $Y2=0.2295
cc_330 N_12_c_569_n N_14_c_629_n 5.93699e-19 $X=1.08 $Y=0.0405 $X2=0.459
+ $Y2=0.2295

* END of "./ASYNC_DFFHx1_ASAP7_75t_SRAM.pex.sp.ASYNC_DFFHX1_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: ICGx1_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:31:37 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "ICGx1_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./ICGx1_ASAP7_75t_SRAM.pex.sp.pex"
* File: ICGx1_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:31:37 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_ICGX1_ASAP7_75T_SRAM%ENA 2 5 7 12 14 VSS
c8 14 VSS 0.00202376f $X=0.081 $Y=0.137
c9 12 VSS 0.00719777f $X=0.082 $Y=0.125
c10 5 VSS 0.002666f $X=0.081 $Y=0.135
c11 2 VSS 0.0610973f $X=0.081 $Y=0.054
r12 12 14 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.125 $X2=0.081 $Y2=0.137
r13 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.137 $X2=0.081
+ $Y2=0.137
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%SE 2 5 7 10 VSS
c11 10 VSS 0.00136133f $X=0.135 $Y=0.125
c12 5 VSS 0.00157649f $X=0.135 $Y=0.135
c13 2 VSS 0.056849f $X=0.135 $Y=0.054
r14 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.125 $X2=0.135 $Y2=0.137
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.137 $X2=0.135
+ $Y2=0.137
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%5 2 5 7 9 10 13 14 17 19 24 26 28 36 40 44 45 46 47
+ 49 VSS
c23 51 VSS 3.08662e-19 $X=0.189 $Y=0.206
c24 49 VSS 9.26001e-20 $X=0.189 $Y=0.198
c25 47 VSS 3.45068e-20 $X=0.189 $Y=0.127
c26 46 VSS 6.5293e-19 $X=0.189 $Y=0.119
c27 45 VSS 4.30607e-19 $X=0.189 $Y=0.09
c28 44 VSS 2.54814e-19 $X=0.189 $Y=0.076
c29 43 VSS 5.02744e-19 $X=0.189 $Y=0.072
c30 40 VSS 8.26035e-19 $X=0.189 $Y=0.135
c31 36 VSS 0.00146362f $X=0.144 $Y=0.036
c32 35 VSS 0.00266146f $X=0.126 $Y=0.036
c33 30 VSS 0.00201059f $X=0.108 $Y=0.036
c34 28 VSS 0.00804964f $X=0.18 $Y=0.036
c35 27 VSS 0.00324205f $X=0.162 $Y=0.233
c36 26 VSS 0.00135162f $X=0.144 $Y=0.233
c37 25 VSS 0.003458f $X=0.126 $Y=0.233
c38 24 VSS 0.00525509f $X=0.09 $Y=0.233
c39 19 VSS 0.00468477f $X=0.18 $Y=0.233
c40 17 VSS 0.00188709f $X=0.056 $Y=0.216
c41 14 VSS 4.96055e-19 $X=0.071 $Y=0.216
c42 13 VSS 0.00796456f $X=0.108 $Y=0.054
c43 9 VSS 5.3314e-19 $X=0.125 $Y=0.054
c44 5 VSS 0.00138612f $X=0.189 $Y=0.135
c45 2 VSS 0.0577976f $X=0.189 $Y=0.0675
r46 52 53 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.223 $X2=0.189 $Y2=0.2235
r47 51 52 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.206 $X2=0.189 $Y2=0.223
r48 50 51 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.199 $X2=0.189 $Y2=0.206
r49 49 50 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.198 $X2=0.189 $Y2=0.199
r50 48 49 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.184 $X2=0.189 $Y2=0.198
r51 46 47 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.119 $X2=0.189 $Y2=0.127
r52 45 46 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.09 $X2=0.189 $Y2=0.119
r53 44 45 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.076 $X2=0.189 $Y2=0.09
r54 43 44 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.072 $X2=0.189 $Y2=0.076
r55 42 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.063 $X2=0.189 $Y2=0.072
r56 40 48 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.184
r57 40 47 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.127
r58 38 53 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.224 $X2=0.189 $Y2=0.2235
r59 37 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r60 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r61 30 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r62 28 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r63 28 36 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.144 $Y2=0.036
r64 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.233 $X2=0.162 $Y2=0.233
r65 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.233 $X2=0.144 $Y2=0.233
r66 24 25 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.233 $X2=0.126 $Y2=0.233
r67 21 24 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.233 $X2=0.09 $Y2=0.233
r68 19 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.233 $X2=0.189 $Y2=0.224
r69 19 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.233 $X2=0.162 $Y2=0.233
r70 17 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.233 $X2=0.054
+ $Y2=0.233
r71 14 17 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r72 13 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r73 10 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.054 $X2=0.108 $Y2=0.054
r74 9 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.054 $X2=0.108 $Y2=0.054
r75 5 40 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r76 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r77 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%CLK 2 5 8 14 17 19 22 27 30 33 35 40 42 45 47 48 49
+ 52 65 66 69 70 71 75 80 91 92 VSS
c90 102 VSS 1.751e-20 $X=0.621 $Y=0.15
c91 92 VSS 6.23569e-19 $X=0.405 $Y=0.134
c92 91 VSS 0.00814038f $X=0.405 $Y=0.134
c93 80 VSS 2.48826e-19 $X=0.621 $Y=0.133
c94 75 VSS 9.46764e-19 $X=0.243 $Y=0.133
c95 71 VSS 6.07691e-19 $X=0.6015 $Y=0.153
c96 70 VSS 0.00403965f $X=0.582 $Y=0.153
c97 69 VSS 0.00101808f $X=0.621 $Y=0.153
c98 68 VSS 0.00158411f $X=0.621 $Y=0.153
c99 66 VSS 0.00143958f $X=0.3595 $Y=0.153
c100 65 VSS 0.00275092f $X=0.296 $Y=0.153
c101 52 VSS 0.00121984f $X=0.756 $Y=0.162
c102 49 VSS 1.21131e-19 $X=0.6935 $Y=0.187
c103 48 VSS 1.74568e-19 $X=0.688 $Y=0.187
c104 47 VSS 4.53034e-19 $X=0.684 $Y=0.187
c105 46 VSS 0.00441397f $X=0.666 $Y=0.187
c106 43 VSS 9.76836e-19 $X=0.63 $Y=0.187
c107 42 VSS 0.00277821f $X=0.747 $Y=0.187
c108 40 VSS 6.61017e-19 $X=0.3555 $Y=0.1335
c109 33 VSS 0.00699063f $X=0.783 $Y=0.162
c110 30 VSS 0.0600574f $X=0.783 $Y=0.0675
c111 22 VSS 0.0600791f $X=0.729 $Y=0.0675
c112 17 VSS 0.00236251f $X=0.621 $Y=0.135
c113 14 VSS 0.0620989f $X=0.621 $Y=0.0675
c114 8 VSS 0.0605267f $X=0.351 $Y=0.0405
c115 2 VSS 0.0605313f $X=0.243 $Y=0.1335
r116 101 102 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.147 $X2=0.621 $Y2=0.15
r117 91 92 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.405 $Y=0.134
+ $X2=0.405 $Y2=0.134
r118 80 101 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.133 $X2=0.621 $Y2=0.147
r119 70 71 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.582
+ $Y=0.153 $X2=0.6015 $Y2=0.153
r120 69 102 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.621 $Y2=0.15
r121 68 71 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.6015 $Y2=0.153
r122 68 69 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.621 $Y=0.153 $X2=0.621
+ $Y2=0.153
r123 65 66 4.31173 $w=1.8e-08 $l=6.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.296
+ $Y=0.153 $X2=0.3595 $Y2=0.153
r124 64 92 0.725694 $w=3.2e-08 $l=3.36861e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4305 $Y=0.153 $X2=0.405 $Y2=0.134
r125 63 70 10.7963 $w=1.8e-08 $l=1.59e-07 $layer=M2 $thickness=3.6e-08 $X=0.423
+ $Y=0.153 $X2=0.582 $Y2=0.153
r126 63 66 4.31173 $w=1.8e-08 $l=6.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.423
+ $Y=0.153 $X2=0.3595 $Y2=0.153
r127 63 64 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.423 $Y=0.153 $X2=0.423
+ $Y2=0.153
r128 60 75 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.133
r129 59 65 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.296 $Y2=0.153
r130 59 60 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.153 $X2=0.243
+ $Y2=0.153
r131 57 69 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.178 $X2=0.621 $Y2=0.153
r132 52 53 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.756 $Y=0.162 $X2=0.756
+ $Y2=0.162
r133 50 52 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.178 $X2=0.756 $Y2=0.162
r134 48 49 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.187 $X2=0.6935 $Y2=0.187
r135 47 48 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.187 $X2=0.688 $Y2=0.187
r136 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.187 $X2=0.684 $Y2=0.187
r137 45 49 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.699
+ $Y=0.187 $X2=0.6935 $Y2=0.187
r138 43 57 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.63 $Y=0.187 $X2=0.621 $Y2=0.178
r139 43 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.187 $X2=0.666 $Y2=0.187
r140 42 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.747 $Y=0.187 $X2=0.756 $Y2=0.178
r141 42 45 3.25926 $w=1.8e-08 $l=4.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.187 $X2=0.699 $Y2=0.187
r142 40 91 41.0143 $w=2.5e-08 $l=4.95e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.3555 $Y=0.1335 $X2=0.405 $Y2=0.1335
r143 33 53 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.783
+ $Y=0.162 $X2=0.756 $Y2=0.162
r144 33 35 202.311 $w=2e-08 $l=5.4e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.162 $X2=0.783 $Y2=0.216
r145 30 33 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.162
r146 25 53 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.162 $X2=0.756 $Y2=0.162
r147 25 27 202.311 $w=2e-08 $l=5.4e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.162 $X2=0.729 $Y2=0.216
r148 22 25 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.162
r149 17 80 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.133 $X2=0.621
+ $Y2=0.133
r150 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2025
r151 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r152 11 40 4.28571 $w=2.1e-08 $l=4.5e-09 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.1335 $X2=0.3555 $Y2=0.1335
r153 8 11 348.425 $w=2e-08 $l=9.3e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0405 $X2=0.351 $Y2=0.1335
r154 2 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.133 $X2=0.243
+ $Y2=0.133
r155 2 5 258.509 $w=2e-08 $l=6.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1335 $X2=0.243 $Y2=0.2025
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%7 2 5 7 9 12 14 17 22 32 34 35 41 43 48 51 52 64 65
+ 67 71 VSS
c61 72 VSS 2.26979e-19 $X=0.308 $Y=0.189
c62 71 VSS 4.78866e-20 $X=0.306 $Y=0.189
c63 67 VSS 4.14661e-19 $X=0.568 $Y=0.222
c64 65 VSS 8.31219e-19 $X=0.568 $Y=0.1525
c65 64 VSS 3.2551e-19 $X=0.568 $Y=0.116
c66 52 VSS 7.99983e-19 $X=0.568 $Y=0.189
c67 51 VSS 0.00784196f $X=0.568 $Y=0.189
c68 48 VSS 7.00345e-19 $X=0.31 $Y=0.189
c69 44 VSS 8.31083e-19 $X=0.5855 $Y=0.232
c70 43 VSS 0.00225204f $X=0.577 $Y=0.232
c71 41 VSS 0.00296213f $X=0.594 $Y=0.232
c72 35 VSS 1.60717e-19 $X=0.5855 $Y=0.086
c73 34 VSS 2.76555e-19 $X=0.577 $Y=0.086
c74 32 VSS 6.35967e-19 $X=0.594 $Y=0.086
c75 22 VSS 0.00293691f $X=0.297 $Y=0.133
c76 17 VSS 0.00522363f $X=0.596 $Y=0.2025
c77 14 VSS 4.06194e-19 $X=0.611 $Y=0.2025
c78 12 VSS 0.006146f $X=0.596 $Y=0.0675
c79 9 VSS 3.3425e-19 $X=0.611 $Y=0.0675
c80 5 VSS 0.00108474f $X=0.297 $Y=0.1335
c81 2 VSS 0.0591582f $X=0.297 $Y=0.0675
r82 71 72 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.189 $X2=0.308 $Y2=0.189
r83 68 71 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.306 $Y2=0.189
r84 66 67 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.196 $X2=0.568 $Y2=0.222
r85 64 65 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.116 $X2=0.568 $Y2=0.1525
r86 52 66 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.189 $X2=0.568 $Y2=0.196
r87 52 65 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.189 $X2=0.568 $Y2=0.1525
r88 51 52 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.568 $Y=0.189 $X2=0.568
+ $Y2=0.189
r89 48 72 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.31
+ $Y=0.189 $X2=0.308 $Y2=0.189
r90 47 51 17.5185 $w=1.8e-08 $l=2.58e-07 $layer=M2 $thickness=3.6e-08 $X=0.31
+ $Y=0.189 $X2=0.568 $Y2=0.189
r91 47 48 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.31 $Y=0.189 $X2=0.31
+ $Y2=0.189
r92 43 44 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.577
+ $Y=0.232 $X2=0.5855 $Y2=0.232
r93 41 44 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.232 $X2=0.5855 $Y2=0.232
r94 38 67 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.223 $X2=0.568 $Y2=0.222
r95 37 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.232 $X2=0.577 $Y2=0.232
r96 37 38 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.232 $X2=0.568 $Y2=0.223
r97 34 35 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.577
+ $Y=0.086 $X2=0.5855 $Y2=0.086
r98 32 35 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.086 $X2=0.5855 $Y2=0.086
r99 29 64 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.095 $X2=0.568 $Y2=0.116
r100 28 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.086 $X2=0.577 $Y2=0.086
r101 28 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.086 $X2=0.568 $Y2=0.095
r102 20 68 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.18 $X2=0.297 $Y2=0.189
r103 20 22 3.19136 $w=1.8e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.18 $X2=0.297 $Y2=0.133
r104 17 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.232
+ $X2=0.594 $Y2=0.232
r105 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2025 $X2=0.596 $Y2=0.2025
r106 12 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.086
+ $X2=0.594 $Y2=0.086
r107 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0675 $X2=0.596 $Y2=0.0675
r108 5 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.133 $X2=0.297
+ $Y2=0.133
r109 5 7 359.664 $w=2e-08 $l=9.6e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.1335 $X2=0.297 $Y2=0.2295
r110 2 5 247.269 $w=2e-08 $l=6.6e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.1335
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%8 2 5 7 9 12 14 17 19 21 30 31 34 35 36 37 38 39 40
+ 42 VSS
c35 48 VSS 0.00202496f $X=0.503 $Y=0.233
c36 47 VSS 0.00196262f $X=0.5125 $Y=0.233
c37 42 VSS 0.00220406f $X=0.486 $Y=0.233
c38 40 VSS 4.74628e-19 $X=0.5125 $Y=0.2115
c39 39 VSS 4.02544e-19 $X=0.5125 $Y=0.199
c40 38 VSS 0.00108412f $X=0.5125 $Y=0.181
c41 37 VSS 3.28082e-19 $X=0.5125 $Y=0.162
c42 36 VSS 7.74522e-19 $X=0.5125 $Y=0.144
c43 35 VSS 6.76213e-19 $X=0.5125 $Y=0.12
c44 34 VSS 7.4117e-19 $X=0.5125 $Y=0.224
c45 32 VSS 2.34081e-20 $X=0.4795 $Y=0.082
c46 31 VSS 3.47256e-19 $X=0.473 $Y=0.082
c47 30 VSS 5.61168e-19 $X=0.447 $Y=0.082
c48 29 VSS 1.3164e-20 $X=0.414 $Y=0.082
c49 21 VSS 3.43763e-19 $X=0.406 $Y=0.082
c50 19 VSS 6.74711e-19 $X=0.503 $Y=0.082
c51 17 VSS 0.0029927f $X=0.484 $Y=0.2295
c52 12 VSS 0.0170022f $X=0.484 $Y=0.0405
c53 5 VSS 0.00244059f $X=0.405 $Y=0.082
c54 2 VSS 0.058916f $X=0.405 $Y=0.0405
r55 48 49 0.322531 $w=1.8e-08 $l=4.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.503
+ $Y=0.233 $X2=0.50775 $Y2=0.233
r56 47 49 0.322531 $w=1.8e-08 $l=4.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.233 $X2=0.50775 $Y2=0.233
r57 42 48 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.233 $X2=0.503 $Y2=0.233
r58 39 40 0.793941 $w=1.9e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.199 $X2=0.5125 $Y2=0.2115
r59 38 39 1.14327 $w=1.9e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.181 $X2=0.5125 $Y2=0.199
r60 37 38 1.20679 $w=1.9e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.162 $X2=0.5125 $Y2=0.181
r61 36 37 1.14327 $w=1.9e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.144 $X2=0.5125 $Y2=0.162
r62 35 36 1.52437 $w=1.9e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.12 $X2=0.5125 $Y2=0.144
r63 34 47 0.0384781 $w=1.9e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.224 $X2=0.5125 $Y2=0.233
r64 34 40 0.793941 $w=1.9e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.224 $X2=0.5125 $Y2=0.2115
r65 33 35 1.84194 $w=1.9e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.091 $X2=0.5125 $Y2=0.12
r66 31 32 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.473
+ $Y=0.082 $X2=0.4795 $Y2=0.082
r67 30 31 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.082 $X2=0.473 $Y2=0.082
r68 29 30 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.082 $X2=0.447 $Y2=0.082
r69 27 32 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.082 $X2=0.4795 $Y2=0.082
r70 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.082 $X2=0.486
+ $Y2=0.082
r71 21 29 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.406
+ $Y=0.082 $X2=0.414 $Y2=0.082
r72 19 33 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.503 $Y=0.082 $X2=0.5125 $Y2=0.091
r73 19 27 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.503
+ $Y=0.082 $X2=0.486 $Y2=0.082
r74 17 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.233 $X2=0.486
+ $Y2=0.233
r75 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2295 $X2=0.484 $Y2=0.2295
r76 12 28 35.8185 $w=2.4e-08 $l=4.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0405 $X2=0.486 $Y2=0.082
r77 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0405 $X2=0.484 $Y2=0.0405
r78 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.406 $Y=0.082 $X2=0.406
+ $Y2=0.082
r79 5 7 552.609 $w=2e-08 $l=1.475e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.082 $X2=0.405 $Y2=0.2295
r80 2 5 155.48 $w=2e-08 $l=4.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0405 $X2=0.405 $Y2=0.082
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%9 2 5 7 10 13 15 18 21 23 25 30 33 37 38 41 43 49
+ 50 53 58 59 60 61 62 64 65 67 68 69 70 72 75 77 79 86 88 89 90 91 93 94 95 96
+ 97 98 101 107 110 VSS
c103 113 VSS 8.41179e-20 $X=0.837 $Y=0.125
c104 110 VSS 3.87592e-19 $X=0.837 $Y=0.133
c105 107 VSS 3.24618e-19 $X=0.837 $Y=0.108
c106 101 VSS 6.17137e-19 $X=0.675 $Y=0.133
c107 99 VSS 4.28973e-19 $X=0.675 $Y=0.108
c108 98 VSS 1.77849e-19 $X=0.358 $Y=0.19
c109 97 VSS 0.00171031f $X=0.358 $Y=0.036
c110 96 VSS 3.16771e-19 $X=0.7965 $Y=0.108
c111 95 VSS 2.5364e-19 $X=0.765 $Y=0.108
c112 94 VSS 7.79718e-20 $X=0.747 $Y=0.108
c113 93 VSS 0.00155044f $X=0.742 $Y=0.108
c114 91 VSS 6.48597e-19 $X=0.828 $Y=0.108
c115 90 VSS 8.07734e-20 $X=0.675 $Y=0.097
c116 89 VSS 4.90266e-19 $X=0.675 $Y=0.095
c117 88 VSS 1.49364e-19 $X=0.675 $Y=0.081
c118 87 VSS 1.86503e-19 $X=0.675 $Y=0.077
c119 86 VSS 5.68609e-19 $X=0.675 $Y=0.073
c120 85 VSS 8.45284e-19 $X=0.675 $Y=0.063
c121 84 VSS 6.05801e-20 $X=0.675 $Y=0.099
c122 80 VSS 5.02745e-19 $X=0.453 $Y=0.19
c123 79 VSS 0.00172533f $X=0.447 $Y=0.19
c124 78 VSS 3.27114e-19 $X=0.396 $Y=0.19
c125 77 VSS 0.00110887f $X=0.392 $Y=0.19
c126 75 VSS 8.20031e-19 $X=0.459 $Y=0.19
c127 72 VSS 0.00146505f $X=0.63 $Y=0.036
c128 71 VSS 2.9457e-19 $X=0.612 $Y=0.036
c129 70 VSS 0.00428093f $X=0.609 $Y=0.036
c130 69 VSS 0.00316044f $X=0.559 $Y=0.036
c131 68 VSS 0.0128572f $X=0.522 $Y=0.036
c132 67 VSS 0.00218374f $X=0.392 $Y=0.036
c133 65 VSS 0.00760762f $X=0.666 $Y=0.036
c134 64 VSS 7.19963e-19 $X=0.358 $Y=0.223
c135 62 VSS 3.15222e-19 $X=0.358 $Y=0.18
c136 61 VSS 3.80467e-19 $X=0.358 $Y=0.162
c137 60 VSS 5.42963e-19 $X=0.358 $Y=0.12
c138 59 VSS 2.16018e-19 $X=0.358 $Y=0.091
c139 57 VSS 5.84318e-19 $X=0.358 $Y=0.072
c140 53 VSS 0.00229455f $X=0.324 $Y=0.036
c141 50 VSS 0.00436152f $X=0.349 $Y=0.036
c142 49 VSS 0.00260946f $X=0.324 $Y=0.232
c143 48 VSS 0.00204527f $X=0.288 $Y=0.232
c144 43 VSS 0.00103077f $X=0.27 $Y=0.232
c145 41 VSS 0.00444971f $X=0.349 $Y=0.232
c146 40 VSS 6.58864e-19 $X=0.27 $Y=0.2295
c147 37 VSS 0.00129546f $X=0.27 $Y=0.2025
c148 32 VSS 5.70081e-19 $X=0.324 $Y=0.0405
c149 21 VSS 0.00222895f $X=0.837 $Y=0.135
c150 18 VSS 0.0576513f $X=0.837 $Y=0.0675
c151 13 VSS 0.00240787f $X=0.675 $Y=0.135
c152 10 VSS 0.0575264f $X=0.675 $Y=0.0675
c153 5 VSS 0.00191265f $X=0.459 $Y=0.19
c154 2 VSS 0.0630025f $X=0.459 $Y=0.0405
r155 112 113 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.117 $X2=0.837 $Y2=0.125
r156 110 113 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.133 $X2=0.837 $Y2=0.125
r157 107 112 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.108 $X2=0.837 $Y2=0.117
r158 103 104 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.116 $X2=0.675 $Y2=0.117
r159 101 104 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.133 $X2=0.675 $Y2=0.117
r160 99 103 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.108 $X2=0.675 $Y2=0.116
r161 95 96 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.765
+ $Y=0.108 $X2=0.7965 $Y2=0.108
r162 94 95 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.108 $X2=0.765 $Y2=0.108
r163 93 94 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.742
+ $Y=0.108 $X2=0.747 $Y2=0.108
r164 92 99 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.108 $X2=0.675 $Y2=0.108
r165 92 93 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.108 $X2=0.742 $Y2=0.108
r166 91 107 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.108 $X2=0.837 $Y2=0.108
r167 91 96 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.108 $X2=0.7965 $Y2=0.108
r168 89 90 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.095 $X2=0.675 $Y2=0.097
r169 88 89 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.081 $X2=0.675 $Y2=0.095
r170 87 88 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.077 $X2=0.675 $Y2=0.081
r171 86 87 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.073 $X2=0.675 $Y2=0.077
r172 85 86 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.063 $X2=0.675 $Y2=0.073
r173 84 99 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.099 $X2=0.675 $Y2=0.108
r174 84 90 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.099 $X2=0.675 $Y2=0.097
r175 83 85 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.045 $X2=0.675 $Y2=0.063
r176 79 80 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.19 $X2=0.453 $Y2=0.19
r177 78 79 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.19 $X2=0.447 $Y2=0.19
r178 77 78 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.392
+ $Y=0.19 $X2=0.396 $Y2=0.19
r179 75 80 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.19 $X2=0.453 $Y2=0.19
r180 73 98 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.19 $X2=0.358 $Y2=0.19
r181 73 77 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.19 $X2=0.392 $Y2=0.19
r182 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.63 $Y2=0.036
r183 70 71 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.609
+ $Y=0.036 $X2=0.612 $Y2=0.036
r184 69 70 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.559
+ $Y=0.036 $X2=0.609 $Y2=0.036
r185 68 69 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.559 $Y2=0.036
r186 67 68 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.392
+ $Y=0.036 $X2=0.522 $Y2=0.036
r187 66 97 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.036 $X2=0.358 $Y2=0.036
r188 66 67 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.036 $X2=0.392 $Y2=0.036
r189 65 83 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.036 $X2=0.675 $Y2=0.045
r190 65 72 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.63 $Y2=0.036
r191 63 98 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.199 $X2=0.358 $Y2=0.19
r192 63 64 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.199 $X2=0.358 $Y2=0.223
r193 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.162 $X2=0.358 $Y2=0.18
r194 60 61 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.12 $X2=0.358 $Y2=0.162
r195 59 60 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.091 $X2=0.358 $Y2=0.12
r196 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.073 $X2=0.358 $Y2=0.091
r197 57 58 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.072 $X2=0.358 $Y2=0.073
r198 56 98 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.181 $X2=0.358 $Y2=0.19
r199 56 62 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.181 $X2=0.358 $Y2=0.18
r200 55 97 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.045 $X2=0.358 $Y2=0.036
r201 55 57 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.045 $X2=0.358 $Y2=0.072
r202 52 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r203 50 97 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.349
+ $Y=0.036 $X2=0.358 $Y2=0.036
r204 50 52 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.349
+ $Y=0.036 $X2=0.324 $Y2=0.036
r205 48 49 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.232 $X2=0.324 $Y2=0.232
r206 43 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.232 $X2=0.288 $Y2=0.232
r207 41 64 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.349 $Y=0.232 $X2=0.358 $Y2=0.223
r208 41 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.349
+ $Y=0.232 $X2=0.324 $Y2=0.232
r209 38 40 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2295 $X2=0.27 $Y2=0.2295
r210 37 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.232 $X2=0.27
+ $Y2=0.232
r211 34 40 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2655 $Y=0.216 $X2=0.27 $Y2=0.2295
r212 34 37 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2655 $Y=0.216 $X2=0.2655 $Y2=0.189
r213 33 37 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.189 $X2=0.2655 $Y2=0.189
r214 30 32 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0405 $X2=0.324 $Y2=0.0405
r215 29 53 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r216 26 32 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.054 $X2=0.324 $Y2=0.0405
r217 26 29 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.054 $X2=0.3195 $Y2=0.081
r218 25 29 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.081 $X2=0.3195 $Y2=0.081
r219 21 110 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.133
+ $X2=0.837 $Y2=0.133
r220 21 23 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.216
r221 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0675 $X2=0.837 $Y2=0.135
r222 13 101 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.133
+ $X2=0.675 $Y2=0.133
r223 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.216
r224 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0675 $X2=0.675 $Y2=0.135
r225 5 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.19 $X2=0.459
+ $Y2=0.19
r226 5 7 147.987 $w=2e-08 $l=3.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.19 $X2=0.459 $Y2=0.2295
r227 2 5 560.102 $w=2e-08 $l=1.495e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0405 $X2=0.459 $Y2=0.19
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%10 2 5 7 9 10 13 14 15 18 19 20 32 33 34 39 46 49
+ 51 52 60 VSS
c33 60 VSS 0.00355073f $X=0.837 $Y=0.228
c34 59 VSS 1.56305e-19 $X=0.837 $Y=0.225
c35 58 VSS 7.65866e-19 $X=0.837 $Y=0.222
c36 56 VSS 0.00240875f $X=0.837 $Y=0.231
c37 52 VSS 4.00315e-19 $X=0.837 $Y=0.197
c38 51 VSS 5.55947e-19 $X=0.891 $Y=0.1675
c39 49 VSS 3.52663e-19 $X=0.891 $Y=0.1175
c40 46 VSS 1.57883e-19 $X=0.891 $Y=0.136
c41 44 VSS 2.26686e-19 $X=0.891 $Y=0.188
c42 41 VSS 0.00388157f $X=0.882 $Y=0.197
c43 40 VSS 0.00379396f $X=0.879 $Y=0.072
c44 39 VSS 0.00352836f $X=0.846 $Y=0.072
c45 34 VSS 6.46932e-20 $X=0.882 $Y=0.072
c46 33 VSS 0.00231927f $X=0.7875 $Y=0.231
c47 32 VSS 0.00805297f $X=0.765 $Y=0.231
c48 23 VSS 0.00658906f $X=0.81 $Y=0.216
c49 19 VSS 6.59309e-19 $X=0.827 $Y=0.216
c50 18 VSS 0.0060288f $X=0.702 $Y=0.216
c51 14 VSS 7.72153e-19 $X=0.719 $Y=0.216
c52 13 VSS 0.004367f $X=0.756 $Y=0.0675
c53 9 VSS 7.90436e-19 $X=0.773 $Y=0.0675
c54 5 VSS 0.00165529f $X=0.891 $Y=0.136
c55 2 VSS 0.061904f $X=0.891 $Y=0.0675
r56 59 60 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.228
r57 58 59 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.222 $X2=0.837 $Y2=0.225
r58 57 58 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.206 $X2=0.837 $Y2=0.222
r59 56 60 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.231 $X2=0.837 $Y2=0.228
r60 52 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.197 $X2=0.837 $Y2=0.206
r61 50 51 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.147 $X2=0.891 $Y2=0.1675
r62 48 49 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.099 $X2=0.891 $Y2=0.1175
r63 46 50 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.136 $X2=0.891 $Y2=0.147
r64 46 49 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.136 $X2=0.891 $Y2=0.1175
r65 44 51 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.188 $X2=0.891 $Y2=0.1675
r66 43 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.081 $X2=0.891 $Y2=0.099
r67 42 52 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.197 $X2=0.837 $Y2=0.197
r68 41 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.197 $X2=0.891 $Y2=0.188
r69 41 42 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.197 $X2=0.846 $Y2=0.197
r70 39 40 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.072 $X2=0.879 $Y2=0.072
r71 36 39 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.072 $X2=0.846 $Y2=0.072
r72 34 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.072 $X2=0.891 $Y2=0.081
r73 34 40 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.072 $X2=0.879 $Y2=0.072
r74 32 33 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.765
+ $Y=0.231 $X2=0.7875 $Y2=0.231
r75 30 33 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.231 $X2=0.7875 $Y2=0.231
r76 26 32 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.231 $X2=0.765 $Y2=0.231
r77 24 56 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.231 $X2=0.837 $Y2=0.231
r78 24 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.231 $X2=0.81 $Y2=0.231
r79 23 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.231 $X2=0.81
+ $Y2=0.231
r80 20 23 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.216 $X2=0.81 $Y2=0.216
r81 19 23 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.216 $X2=0.81 $Y2=0.216
r82 18 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.231 $X2=0.702
+ $Y2=0.231
r83 15 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.216 $X2=0.702 $Y2=0.216
r84 14 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.216 $X2=0.702 $Y2=0.216
r85 13 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.072 $X2=0.756
+ $Y2=0.072
r86 10 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.756 $Y2=0.0675
r87 9 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.756 $Y2=0.0675
r88 5 46 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.136 $X2=0.891
+ $Y2=0.136
r89 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.136 $X2=0.891 $Y2=0.2025
r90 2 5 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.0675 $X2=0.891 $Y2=0.136
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%GCLK 1 6 9 11 14 17 25 27 VSS
c7 29 VSS 4.30151e-19 $X=0.945 $Y=0.2155
c8 27 VSS 0.00211336f $X=0.945 $Y=0.1145
c9 26 VSS 8.85605e-19 $X=0.945 $Y=0.063
c10 25 VSS 0.00385168f $X=0.945 $Y=0.166
c11 23 VSS 4.55454e-19 $X=0.945 $Y=0.225
c12 17 VSS 0.00196563f $X=0.918 $Y=0.234
c13 15 VSS 0.00604756f $X=0.936 $Y=0.234
c14 14 VSS 0.00623927f $X=0.918 $Y=0.036
c15 11 VSS 0.0100986f $X=0.936 $Y=0.036
c16 9 VSS 0.00664317f $X=0.916 $Y=0.2025
c17 4 VSS 2.69461e-19 $X=0.916 $Y=0.0675
r18 28 29 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.206 $X2=0.945 $Y2=0.2155
r19 26 27 3.49691 $w=1.8e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.063 $X2=0.945 $Y2=0.1145
r20 25 28 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.166 $X2=0.945 $Y2=0.206
r21 25 27 3.49691 $w=1.8e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.166 $X2=0.945 $Y2=0.1145
r22 23 29 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.2155
r23 22 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.063
r24 15 23 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r25 15 17 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.918 $Y2=0.234
r26 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.036 $X2=0.918
+ $Y2=0.036
r27 11 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r28 11 13 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.918 $Y2=0.036
r29 9 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.234 $X2=0.918
+ $Y2=0.234
r30 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.901
+ $Y=0.2025 $X2=0.916 $Y2=0.2025
r31 4 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.918
+ $Y=0.0675 $X2=0.918 $Y2=0.036
r32 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.901
+ $Y=0.0675 $X2=0.916 $Y2=0.0675
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%12 1 6 9 VSS
c9 9 VSS 0.0194635f $X=0.272 $Y=0.0675
c10 6 VSS 3.61939e-19 $X=0.287 $Y=0.0675
c11 4 VSS 3.25039e-19 $X=0.214 $Y=0.0675
r12 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.272 $Y2=0.0675
r13 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.214
+ $Y=0.0675 $X2=0.272 $Y2=0.0675
r14 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.214 $Y2=0.0675
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%13 1 2 5 VSS
c5 5 VSS 0.00582405f $X=0.216 $Y=0.2025
c6 1 VSS 6.50078e-19 $X=0.233 $Y=0.2025
r7 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.2025 $X2=0.216 $Y2=0.2025
r8 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.216 $Y2=0.2025
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%14 1 6 9 VSS
c10 9 VSS 0.0186419f $X=0.38 $Y=0.2295
c11 6 VSS 3.72954e-19 $X=0.395 $Y=0.2295
c12 4 VSS 3.77944e-19 $X=0.322 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.2295 $X2=0.38 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.2295 $X2=0.38 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2295 $X2=0.322 $Y2=0.2295
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%15 1 2 5 VSS
c4 5 VSS 0.004225f $X=0.378 $Y=0.0405
c5 1 VSS 6.8236e-19 $X=0.395 $Y=0.0405
r6 2 5 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.0405 $X2=0.378 $Y2=0.0405
r7 1 5 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0405 $X2=0.378 $Y2=0.0405
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%16 1 2 VSS
c1 1 VSS 0.00221026f $X=0.719 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0675 $X2=0.685 $Y2=0.0675
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%17 1 2 VSS
c2 1 VSS 0.00230546f $X=0.827 $Y=0.0675
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.827
+ $Y=0.0675 $X2=0.793 $Y2=0.0675
.ends

.subckt PM_ICGX1_ASAP7_75T_SRAM%18 1 2 VSS
c0 1 VSS 0.00242486f $X=0.125 $Y=0.216
r1 1 2 25.1852 $w=5.4e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.216 $X2=0.091 $Y2=0.216
.ends


* END of "./ICGx1_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt ICGx1_ASAP7_75t_SRAM  VSS VDD ENA SE CLK GCLK
* 
* GCLK	GCLK
* CLK	CLK
* SE	SE
* ENA	ENA
M0 N_5_M0_d N_ENA_M0_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 VSS N_SE_M1_g N_5_M1_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 N_12_M2_d N_5_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_9_M3_d N_7_M3_g N_12_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M4 N_15_M4_d N_CLK_M4_g N_9_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.341
+ $Y=0.027
M5 VSS N_8_M5_g N_15_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.395
+ $Y=0.027
M6 N_8_M6_d N_9_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449 $Y=0.027
M7 VSS N_CLK_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M8 VSS N_9_M8_g N_16_M8_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M9 N_16_M9_d N_CLK_M9_g N_10_M9_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M10 N_17_M10_d N_CLK_M10_g N_10_M10_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.773 $Y=0.027
M11 VSS N_9_M11_g N_17_M11_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.027
M12 N_GCLK_M12_d N_10_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.027
M13 N_18_M13_d N_ENA_M13_g N_5_M13_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.071 $Y=0.189
M14 VDD N_SE_M14_g N_18_M14_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M15 N_13_M15_d N_5_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M16 N_9_M16_d N_CLK_M16_g N_13_M16_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M17 N_14_M17_d N_7_M17_g N_9_M17_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.287 $Y=0.216
M18 VDD N_8_M18_g N_14_M18_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.395
+ $Y=0.216
M19 N_8_M19_d N_9_M19_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.216
M20 VDD N_CLK_M20_g N_7_M20_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M21 N_10_M21_d N_9_M21_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.665
+ $Y=0.189
M22 VDD N_CLK_M22_g N_10_M22_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.719
+ $Y=0.189
M23 VDD N_CLK_M23_g N_10_M23_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.773
+ $Y=0.189
M24 N_10_M24_d N_9_M24_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.827
+ $Y=0.189
M25 N_GCLK_M25_d N_10_M25_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.162
*
* 
* .include "ICGx1_ASAP7_75t_SRAM.pex.sp.ICGX1_ASAP7_75T_SRAM.pxi"
* BEGIN of "./ICGx1_ASAP7_75t_SRAM.pex.sp.ICGX1_ASAP7_75T_SRAM.pxi"
* File: ICGx1_ASAP7_75t_SRAM.pex.sp.ICGX1_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:31:37 2017
* 
x_PM_ICGX1_ASAP7_75T_SRAM%ENA N_ENA_M0_g N_ENA_c_2_p N_ENA_M13_g ENA N_ENA_c_6_p
+ VSS PM_ICGX1_ASAP7_75T_SRAM%ENA
x_PM_ICGX1_ASAP7_75T_SRAM%SE N_SE_M1_g N_SE_c_10_n N_SE_M14_g SE VSS
+ PM_ICGX1_ASAP7_75T_SRAM%SE
x_PM_ICGX1_ASAP7_75T_SRAM%5 N_5_M2_g N_5_c_26_n N_5_M15_g N_5_M1_s N_5_M0_d
+ N_5_c_21_n N_5_M13_s N_5_c_22_n N_5_c_40_p N_5_c_23_n N_5_c_27_n N_5_c_41_p
+ N_5_c_29_n N_5_c_34_p N_5_c_37_p N_5_c_31_n N_5_c_38_p N_5_c_35_p N_5_c_39_p
+ VSS PM_ICGX1_ASAP7_75T_SRAM%5
x_PM_ICGX1_ASAP7_75T_SRAM%CLK N_CLK_c_43_n N_CLK_M16_g N_CLK_M4_g N_CLK_M7_g
+ N_CLK_c_85_p N_CLK_M20_g N_CLK_M9_g N_CLK_M22_g N_CLK_M10_g N_CLK_c_108_p
+ N_CLK_M23_g N_CLK_c_51_p N_CLK_c_118_p CLK N_CLK_c_84_p N_CLK_c_109_p
+ N_CLK_c_110_p N_CLK_c_111_p N_CLK_c_46_n N_CLK_c_56_p N_CLK_c_53_p
+ N_CLK_c_59_p N_CLK_c_52_p N_CLK_c_47_n N_CLK_c_66_p N_CLK_c_69_p N_CLK_c_62_p
+ VSS PM_ICGX1_ASAP7_75T_SRAM%CLK
x_PM_ICGX1_ASAP7_75T_SRAM%7 N_7_M3_g N_7_c_139_n N_7_M17_g N_7_M7_s N_7_c_141_n
+ N_7_M20_s N_7_c_142_n N_7_c_134_n N_7_c_147_n N_7_c_161_p N_7_c_148_n
+ N_7_c_191_p N_7_c_162_p N_7_c_149_n N_7_c_150_n N_7_c_152_n N_7_c_163_p
+ N_7_c_154_n N_7_c_156_n N_7_c_136_n VSS PM_ICGX1_ASAP7_75T_SRAM%7
x_PM_ICGX1_ASAP7_75T_SRAM%8 N_8_M5_g N_8_c_219_p N_8_M18_g N_8_M6_d N_8_c_197_n
+ N_8_M19_d N_8_c_207_n N_8_c_209_n N_8_c_198_n N_8_c_199_n N_8_c_201_n
+ N_8_c_210_n N_8_c_211_n N_8_c_202_n N_8_c_203_n N_8_c_213_n N_8_c_214_n
+ N_8_c_215_n N_8_c_216_n VSS PM_ICGX1_ASAP7_75T_SRAM%8
x_PM_ICGX1_ASAP7_75T_SRAM%9 N_9_M6_g N_9_c_231_n N_9_M19_g N_9_M8_g N_9_c_236_n
+ N_9_M21_g N_9_M11_g N_9_c_302_p N_9_M24_g N_9_M3_d N_9_M4_s N_9_M16_d
+ N_9_c_239_n N_9_M17_s N_9_c_269_n N_9_c_229_n N_9_c_270_n N_9_c_242_n
+ N_9_c_243_n N_9_c_275_n N_9_c_276_n N_9_c_244_n N_9_c_245_n N_9_c_250_n
+ N_9_c_325_p N_9_c_303_p N_9_c_328_p N_9_c_295_n N_9_c_251_n N_9_c_279_n
+ N_9_c_252_n N_9_c_282_n N_9_c_254_n N_9_c_256_n N_9_c_310_p N_9_c_285_n
+ N_9_c_304_p N_9_c_286_n N_9_c_331_p N_9_c_258_n N_9_c_261_n N_9_c_262_n
+ N_9_c_263_n N_9_c_329_p N_9_c_287_n N_9_c_265_n N_9_c_313_p N_9_c_312_p VSS
+ PM_ICGX1_ASAP7_75T_SRAM%9
x_PM_ICGX1_ASAP7_75T_SRAM%10 N_10_M12_g N_10_c_343_n N_10_M25_g N_10_M10_s
+ N_10_M9_s N_10_c_333_n N_10_M22_s N_10_M21_d N_10_c_334_n N_10_M24_d
+ N_10_M23_s N_10_c_336_n N_10_c_338_n N_10_c_359_p N_10_c_340_n N_10_c_353_n
+ N_10_c_354_n N_10_c_357_p N_10_c_355_n N_10_c_356_n VSS
+ PM_ICGX1_ASAP7_75T_SRAM%10
x_PM_ICGX1_ASAP7_75T_SRAM%GCLK N_GCLK_M12_d N_GCLK_M25_d N_GCLK_c_365_n
+ N_GCLK_c_366_n N_GCLK_c_368_n N_GCLK_c_369_n GCLK N_GCLK_c_371_n VSS
+ PM_ICGX1_ASAP7_75T_SRAM%GCLK
x_PM_ICGX1_ASAP7_75T_SRAM%12 N_12_M2_d N_12_M3_s N_12_c_372_n VSS
+ PM_ICGX1_ASAP7_75T_SRAM%12
x_PM_ICGX1_ASAP7_75T_SRAM%13 N_13_M16_s N_13_M15_d N_13_c_381_n VSS
+ PM_ICGX1_ASAP7_75T_SRAM%13
x_PM_ICGX1_ASAP7_75T_SRAM%14 N_14_M17_d N_14_M18_s N_14_c_386_n VSS
+ PM_ICGX1_ASAP7_75T_SRAM%14
x_PM_ICGX1_ASAP7_75T_SRAM%15 N_15_M5_s N_15_M4_d N_15_c_396_n VSS
+ PM_ICGX1_ASAP7_75T_SRAM%15
x_PM_ICGX1_ASAP7_75T_SRAM%16 N_16_M9_d N_16_M8_s VSS PM_ICGX1_ASAP7_75T_SRAM%16
x_PM_ICGX1_ASAP7_75T_SRAM%17 N_17_M11_s N_17_M10_d VSS PM_ICGX1_ASAP7_75T_SRAM%17
x_PM_ICGX1_ASAP7_75T_SRAM%18 N_18_M14_s N_18_M13_d VSS PM_ICGX1_ASAP7_75T_SRAM%18
cc_1 N_ENA_M0_g N_SE_M1_g 0.00328721f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_ENA_c_2_p N_SE_c_10_n 9.35826e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 ENA SE 0.00588002f $X=0.082 $Y=0.125 $X2=0.135 $Y2=0.125
cc_4 N_ENA_M0_g N_5_M2_g 2.13359e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 ENA N_5_c_21_n 6.06976e-19 $X=0.082 $Y=0.125 $X2=0.135 $Y2=0.137
cc_6 N_ENA_c_6_p N_5_c_22_n 0.00176249f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_7 N_ENA_M0_g N_5_c_23_n 2.28086e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_8 N_ENA_c_6_p N_5_c_23_n 0.00499899f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_9 N_SE_M1_g N_5_M2_g 0.00268443f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_10 N_SE_c_10_n N_5_c_26_n 9.11034e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_11 N_SE_M1_g N_5_c_27_n 2.59938e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_12 SE N_5_c_27_n 0.00123553f $X=0.135 $Y=0.125 $X2=0 $Y2=0
cc_13 N_SE_M1_g N_5_c_29_n 2.84283e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_14 SE N_5_c_29_n 0.001038f $X=0.135 $Y=0.125 $X2=0 $Y2=0
cc_15 SE N_5_c_31_n 0.00457266f $X=0.135 $Y=0.125 $X2=0 $Y2=0
cc_16 N_SE_M1_g N_CLK_c_43_n 2.13359e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_17 N_5_M2_g N_CLK_c_43_n 0.00341068f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_18 N_5_c_26_n N_CLK_c_43_n 8.10277e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.054
cc_19 N_5_c_34_p N_CLK_c_46_n 3.51913e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_20 N_5_c_35_p N_CLK_c_47_n 0.00253596f $X=0.189 $Y=0.127 $X2=0 $Y2=0
cc_21 N_5_M2_g N_7_M3_g 2.82885e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_22 N_5_c_37_p N_7_c_134_n 3.23824e-19 $X=0.189 $Y=0.076 $X2=0 $Y2=0
cc_23 N_5_c_38_p N_7_c_134_n 2.18117e-19 $X=0.189 $Y=0.119 $X2=0 $Y2=0
cc_24 N_5_c_39_p N_7_c_136_n 2.18117e-19 $X=0.189 $Y=0.198 $X2=0 $Y2=0
cc_25 N_5_c_40_p N_9_c_229_n 4.49022e-19 $X=0.18 $Y=0.233 $X2=0 $Y2=0
cc_26 N_5_c_41_p N_12_c_372_n 0.00246673f $X=0.18 $Y=0.036 $X2=0 $Y2=0
cc_27 N_5_c_34_p N_13_c_381_n 0.00181721f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_28 N_CLK_c_43_n N_7_M3_g 0.00355599f $X=0.243 $Y=0.1335 $X2=0.135 $Y2=0.054
cc_29 N_CLK_M4_g N_7_M3_g 0.00355599f $X=0.351 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_30 N_CLK_c_43_n N_7_c_139_n 8.50652e-19 $X=0.243 $Y=0.1335 $X2=0.135
+ $Y2=0.135
cc_31 N_CLK_c_51_p N_7_c_139_n 9.47532e-19 $X=0.3555 $Y=0.1335 $X2=0.135
+ $Y2=0.135
cc_32 N_CLK_c_52_p N_7_c_141_n 2.51466e-19 $X=0.6015 $Y=0.153 $X2=0.135
+ $Y2=0.137
cc_33 N_CLK_c_53_p N_7_c_142_n 6.13009e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_34 N_CLK_c_52_p N_7_c_142_n 2.98103e-19 $X=0.6015 $Y=0.153 $X2=0 $Y2=0
cc_35 N_CLK_c_46_n N_7_c_134_n 0.0010183f $X=0.296 $Y=0.153 $X2=0 $Y2=0
cc_36 N_CLK_c_56_p N_7_c_134_n 5.3655e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_37 N_CLK_c_47_n N_7_c_134_n 0.00252905f $X=0.243 $Y=0.133 $X2=0 $Y2=0
cc_38 N_CLK_c_52_p N_7_c_147_n 2.62247e-19 $X=0.6015 $Y=0.153 $X2=0 $Y2=0
cc_39 N_CLK_c_59_p N_7_c_148_n 2.62247e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_40 N_CLK_c_56_p N_7_c_149_n 2.46239e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_41 N_CLK_c_56_p N_7_c_150_n 0.0242262f $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_42 N_CLK_c_62_p N_7_c_150_n 4.84045e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_43 N_CLK_c_53_p N_7_c_152_n 0.0017697f $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_44 N_CLK_c_59_p N_7_c_152_n 4.75571e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_45 N_CLK_c_59_p N_7_c_154_n 4.04804e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_46 N_CLK_c_66_p N_7_c_154_n 0.00167205f $X=0.621 $Y=0.133 $X2=0 $Y2=0
cc_47 N_CLK_c_59_p N_7_c_156_n 2.46239e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_48 N_CLK_M4_g N_8_M5_g 0.00341068f $X=0.351 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_49 N_CLK_c_69_p N_8_M5_g 0.00207156f $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.054
cc_50 N_CLK_c_62_p N_8_M5_g 2.24185e-19 $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.054
cc_51 N_CLK_c_59_p N_8_c_197_n 2.35254e-19 $X=0.582 $Y=0.153 $X2=0.135 $Y2=0.137
cc_52 N_CLK_c_62_p N_8_c_198_n 8.28523e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_53 N_CLK_c_59_p N_8_c_199_n 3.19268e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_54 N_CLK_c_62_p N_8_c_199_n 0.00100806f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_55 N_CLK_c_59_p N_8_c_201_n 9.01736e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_56 N_CLK_c_62_p N_8_c_202_n 3.57731e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_57 N_CLK_c_59_p N_8_c_203_n 6.50246e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_58 N_CLK_c_62_p N_8_c_203_n 4.93535e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_59 N_CLK_M4_g N_9_M6_g 2.13359e-19 $X=0.351 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_60 N_CLK_c_59_p N_9_c_231_n 2.15534e-19 $X=0.582 $Y=0.153 $X2=0.135 $Y2=0.135
cc_61 N_CLK_M7_g N_9_M8_g 0.00268443f $X=0.621 $Y=0.0675 $X2=0.135 $Y2=0.125
cc_62 N_CLK_M9_g N_9_M8_g 0.00328721f $X=0.729 $Y=0.0675 $X2=0.135 $Y2=0.125
cc_63 N_CLK_M10_g N_9_M8_g 2.48122e-19 $X=0.783 $Y=0.0675 $X2=0.135 $Y2=0.125
cc_64 N_CLK_c_84_p N_9_M8_g 3.92861e-19 $X=0.684 $Y=0.187 $X2=0.135 $Y2=0.125
cc_65 N_CLK_c_85_p N_9_c_236_n 0.0010353f $X=0.621 $Y=0.135 $X2=0.135 $Y2=0.137
cc_66 N_CLK_M9_g N_9_M11_g 2.48122e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_67 N_CLK_M10_g N_9_M11_g 0.00328721f $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_68 N_CLK_c_46_n N_9_c_239_n 3.0124e-19 $X=0.296 $Y=0.153 $X2=0 $Y2=0
cc_69 N_CLK_c_47_n N_9_c_239_n 5.62774e-19 $X=0.243 $Y=0.133 $X2=0 $Y2=0
cc_70 N_CLK_c_46_n N_9_c_229_n 3.44788e-19 $X=0.296 $Y=0.153 $X2=0 $Y2=0
cc_71 N_CLK_c_56_p N_9_c_242_n 4.44284e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_72 N_CLK_c_56_p N_9_c_243_n 2.54113e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_73 N_CLK_M4_g N_9_c_244_n 2.69763e-19 $X=0.351 $Y=0.0405 $X2=0 $Y2=0
cc_74 N_CLK_c_51_p N_9_c_245_n 5.33107e-19 $X=0.3555 $Y=0.1335 $X2=0 $Y2=0
cc_75 N_CLK_c_56_p N_9_c_245_n 4.41663e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_76 N_CLK_c_59_p N_9_c_245_n 3.17785e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_77 N_CLK_c_69_p N_9_c_245_n 0.00207315f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_78 N_CLK_c_62_p N_9_c_245_n 0.00252282f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_79 N_CLK_M4_g N_9_c_250_n 2.92102e-19 $X=0.351 $Y=0.0405 $X2=0 $Y2=0
cc_80 N_CLK_c_59_p N_9_c_251_n 6.2848e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_81 N_CLK_M7_g N_9_c_252_n 3.73075e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_82 N_CLK_c_66_p N_9_c_252_n 4.18576e-19 $X=0.621 $Y=0.133 $X2=0 $Y2=0
cc_83 N_CLK_c_59_p N_9_c_254_n 2.73788e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_84 N_CLK_c_69_p N_9_c_254_n 3.82241e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_85 N_CLK_c_59_p N_9_c_256_n 3.8223e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_86 N_CLK_c_62_p N_9_c_256_n 0.00487387f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_87 N_CLK_M9_g N_9_c_258_n 5.5355e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_88 N_CLK_c_108_p N_9_c_258_n 7.26266e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_89 N_CLK_c_109_p N_9_c_258_n 8.01493e-19 $X=0.688 $Y=0.187 $X2=0 $Y2=0
cc_90 N_CLK_c_110_p N_9_c_261_n 8.01493e-19 $X=0.6935 $Y=0.187 $X2=0 $Y2=0
cc_91 N_CLK_c_111_p N_9_c_262_n 0.00118098f $X=0.756 $Y=0.162 $X2=0 $Y2=0
cc_92 N_CLK_M10_g N_9_c_263_n 3.81593e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_93 N_CLK_c_108_p N_9_c_263_n 8.51921e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_94 N_CLK_c_84_p N_9_c_265_n 9.869e-19 $X=0.684 $Y=0.187 $X2=0 $Y2=0
cc_95 N_CLK_c_66_p N_9_c_265_n 0.00110905f $X=0.621 $Y=0.133 $X2=0 $Y2=0
cc_96 N_CLK_M10_g N_10_M12_g 2.13359e-19 $X=0.783 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_97 N_CLK_c_108_p N_10_c_333_n 7.52823e-19 $X=0.783 $Y=0.162 $X2=0.135
+ $Y2=0.137
cc_98 N_CLK_c_118_p N_10_c_334_n 0.049634f $X=0.747 $Y=0.187 $X2=0 $Y2=0
cc_99 N_CLK_c_110_p N_10_c_334_n 0.0086729f $X=0.6935 $Y=0.187 $X2=0 $Y2=0
cc_100 N_CLK_M9_g N_10_c_336_n 2.89162e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_101 N_CLK_c_110_p N_10_c_336_n 0.00454542f $X=0.6935 $Y=0.187 $X2=0 $Y2=0
cc_102 N_CLK_M10_g N_10_c_338_n 2.82957e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_103 N_CLK_c_108_p N_10_c_338_n 3.8451e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_104 N_CLK_M10_g N_10_c_340_n 3.96202e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_105 N_CLK_c_43_n N_12_c_372_n 0.00569573f $X=0.243 $Y=0.1335 $X2=0.135
+ $Y2=0.125
cc_106 N_CLK_c_46_n N_12_c_372_n 3.78132e-19 $X=0.296 $Y=0.153 $X2=0.135
+ $Y2=0.125
cc_107 N_CLK_c_47_n N_12_c_372_n 3.48512e-19 $X=0.243 $Y=0.133 $X2=0.135
+ $Y2=0.125
cc_108 N_CLK_c_47_n N_13_c_381_n 5.62774e-19 $X=0.243 $Y=0.133 $X2=0.135
+ $Y2=0.135
cc_109 N_CLK_M4_g N_14_c_386_n 0.00280362f $X=0.351 $Y=0.0405 $X2=0.135
+ $Y2=0.125
cc_110 N_CLK_c_51_p N_14_c_386_n 2.06383e-19 $X=0.3555 $Y=0.1335 $X2=0.135
+ $Y2=0.125
cc_111 N_CLK_c_69_p N_14_c_386_n 9.52591e-19 $X=0.405 $Y=0.134 $X2=0.135
+ $Y2=0.125
cc_112 N_CLK_c_69_p N_15_c_396_n 8.7631e-19 $X=0.405 $Y=0.134 $X2=0.135
+ $Y2=0.135
cc_113 N_7_M3_g N_8_M5_g 2.82885e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_114 N_7_c_141_n N_8_c_197_n 0.00121003f $X=0.596 $Y=0.0675 $X2=0 $Y2=0
cc_115 N_7_c_142_n N_8_c_207_n 4.7624e-19 $X=0.596 $Y=0.2025 $X2=0.056 $Y2=0.216
cc_116 N_7_c_150_n N_8_c_207_n 2.60284e-19 $X=0.568 $Y=0.189 $X2=0.056 $Y2=0.216
cc_117 N_7_c_161_p N_8_c_209_n 0.00134983f $X=0.577 $Y=0.086 $X2=0.18 $Y2=0.233
cc_118 N_7_c_162_p N_8_c_210_n 0.00134983f $X=0.577 $Y=0.232 $X2=0 $Y2=0
cc_119 N_7_c_163_p N_8_c_211_n 0.00134983f $X=0.568 $Y=0.116 $X2=0.126 $Y2=0.036
cc_120 N_7_c_154_n N_8_c_203_n 0.00134983f $X=0.568 $Y=0.1525 $X2=0.189
+ $Y2=0.045
cc_121 N_7_c_152_n N_8_c_213_n 0.00134983f $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.224
cc_122 N_7_c_150_n N_8_c_214_n 6.67324e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.135
cc_123 N_7_c_156_n N_8_c_215_n 0.00134983f $X=0.568 $Y=0.222 $X2=0.189 $Y2=0.135
cc_124 N_7_c_150_n N_8_c_216_n 5.91796e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.063
cc_125 N_7_c_142_n N_9_c_231_n 2.39572e-19 $X=0.596 $Y=0.2025 $X2=0.189
+ $Y2=0.135
cc_126 N_7_c_134_n N_9_c_239_n 0.00130909f $X=0.297 $Y=0.133 $X2=0.189 $Y2=0.045
cc_127 N_7_c_150_n N_9_c_269_n 5.00653e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.135
cc_128 N_7_M3_g N_9_c_270_n 2.70372e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.198
cc_129 N_7_c_149_n N_9_c_270_n 4.88088e-19 $X=0.31 $Y=0.189 $X2=0.189 $Y2=0.198
cc_130 N_7_c_150_n N_9_c_270_n 3.79017e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.198
cc_131 N_7_c_136_n N_9_c_270_n 0.00265354f $X=0.306 $Y=0.189 $X2=0.189 $Y2=0.198
cc_132 N_7_c_134_n N_9_c_243_n 0.0011395f $X=0.297 $Y=0.133 $X2=0.189 $Y2=0.2235
cc_133 N_7_c_134_n N_9_c_275_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_134 N_7_c_134_n N_9_c_276_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_135 N_7_c_134_n N_9_c_244_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_136 N_7_c_134_n N_9_c_245_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_137 N_7_M7_s N_9_c_279_n 3.12749e-19 $X=0.611 $Y=0.0675 $X2=0 $Y2=0
cc_138 N_7_c_141_n N_9_c_279_n 0.00290811f $X=0.596 $Y=0.0675 $X2=0 $Y2=0
cc_139 N_7_c_161_p N_9_c_279_n 0.0027674f $X=0.577 $Y=0.086 $X2=0 $Y2=0
cc_140 N_7_c_150_n N_9_c_282_n 2.35423e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_141 N_7_c_150_n N_9_c_254_n 3.37429e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_142 N_7_c_150_n N_9_c_256_n 6.95518e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_143 N_7_c_147_n N_9_c_285_n 3.43042e-19 $X=0.594 $Y=0.086 $X2=0 $Y2=0
cc_144 N_7_c_163_p N_9_c_286_n 2.63767e-19 $X=0.568 $Y=0.116 $X2=0 $Y2=0
cc_145 N_7_c_149_n N_9_c_287_n 0.00126174f $X=0.31 $Y=0.189 $X2=0 $Y2=0
cc_146 N_7_c_150_n N_9_c_287_n 4.35645e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_147 N_7_c_191_p N_10_c_336_n 2.63066e-19 $X=0.594 $Y=0.232 $X2=0 $Y2=0
cc_148 N_7_c_134_n N_12_c_372_n 0.00330923f $X=0.297 $Y=0.133 $X2=0.125
+ $Y2=0.054
cc_149 N_7_c_150_n N_14_c_386_n 3.19426e-19 $X=0.568 $Y=0.189 $X2=0.125
+ $Y2=0.054
cc_150 N_8_M5_g N_9_M6_g 0.00268443f $X=0.405 $Y=0.0405 $X2=0.243 $Y2=0.1335
cc_151 N_8_c_201_n N_9_M6_g 5.07993e-19 $X=0.473 $Y=0.082 $X2=0.243 $Y2=0.1335
cc_152 N_8_c_219_p N_9_c_243_n 5.2508e-19 $X=0.405 $Y=0.082 $X2=0.756 $Y2=0.162
cc_153 N_8_c_198_n N_9_c_276_n 0.00112828f $X=0.406 $Y=0.082 $X2=0.243 $Y2=0.153
cc_154 N_8_c_211_n N_9_c_244_n 2.05549e-19 $X=0.5125 $Y=0.12 $X2=0.243 $Y2=0.153
cc_155 N_8_c_213_n N_9_c_245_n 2.05549e-19 $X=0.5125 $Y=0.181 $X2=0 $Y2=0
cc_156 N_8_M5_g N_9_c_295_n 2.1403e-19 $X=0.405 $Y=0.0405 $X2=0.621 $Y2=0.153
cc_157 N_8_c_197_n N_9_c_295_n 0.00315628f $X=0.484 $Y=0.0405 $X2=0.621
+ $Y2=0.153
cc_158 N_8_c_198_n N_9_c_295_n 0.00735896f $X=0.406 $Y=0.082 $X2=0.621 $Y2=0.153
cc_159 N_8_c_214_n N_9_c_282_n 9.42345e-19 $X=0.5125 $Y=0.199 $X2=0.243
+ $Y2=0.133
cc_160 N_8_c_216_n N_9_c_282_n 2.89066e-19 $X=0.486 $Y=0.233 $X2=0.243 $Y2=0.133
cc_161 N_8_M5_g N_9_c_256_n 5.18398e-19 $X=0.405 $Y=0.0405 $X2=0.621 $Y2=0.133
cc_162 N_9_M11_g N_10_M12_g 0.00268443f $X=0.837 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_163 N_9_c_302_p N_10_c_343_n 9.58586e-19 $X=0.837 $Y=0.135 $X2=0.189
+ $Y2=0.135
cc_164 N_9_c_303_p N_10_c_333_n 6.30417e-19 $X=0.666 $Y=0.036 $X2=0.108
+ $Y2=0.054
cc_165 N_9_c_304_p N_10_c_333_n 2.62833e-19 $X=0.675 $Y=0.095 $X2=0.108
+ $Y2=0.054
cc_166 N_9_c_261_n N_10_c_333_n 5.00181e-19 $X=0.747 $Y=0.108 $X2=0.108
+ $Y2=0.054
cc_167 N_9_c_262_n N_10_c_333_n 0.00105563f $X=0.765 $Y=0.108 $X2=0.108
+ $Y2=0.054
cc_168 N_9_c_263_n N_10_c_333_n 5.00181e-19 $X=0.7965 $Y=0.108 $X2=0.108
+ $Y2=0.054
cc_169 N_9_c_258_n N_10_c_338_n 4.7867e-19 $X=0.742 $Y=0.108 $X2=0 $Y2=0
cc_170 N_9_M11_g N_10_c_340_n 3.37536e-19 $X=0.837 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_171 N_9_c_310_p N_10_c_340_n 5.50762e-19 $X=0.675 $Y=0.073 $X2=0.189
+ $Y2=0.135
cc_172 N_9_c_261_n N_10_c_340_n 0.00883267f $X=0.747 $Y=0.108 $X2=0.189
+ $Y2=0.135
cc_173 N_9_c_312_p N_10_c_353_n 0.00104908f $X=0.837 $Y=0.133 $X2=0.189
+ $Y2=0.119
cc_174 N_9_c_313_p N_10_c_354_n 0.00104908f $X=0.837 $Y=0.108 $X2=0.189
+ $Y2=0.198
cc_175 N_9_c_312_p N_10_c_355_n 8.04994e-19 $X=0.837 $Y=0.133 $X2=0.189
+ $Y2=0.223
cc_176 N_9_c_262_n N_10_c_356_n 4.7867e-19 $X=0.765 $Y=0.108 $X2=0 $Y2=0
cc_177 N_9_c_239_n N_12_c_372_n 0.00144308f $X=0.27 $Y=0.2025 $X2=0.125
+ $Y2=0.054
cc_178 N_9_c_242_n N_12_c_372_n 5.41912e-19 $X=0.349 $Y=0.036 $X2=0.125
+ $Y2=0.054
cc_179 N_9_c_243_n N_12_c_372_n 0.00307808f $X=0.324 $Y=0.036 $X2=0.125
+ $Y2=0.054
cc_180 N_9_c_239_n N_13_c_381_n 0.00390769f $X=0.27 $Y=0.2025 $X2=0.189
+ $Y2=0.135
cc_181 N_9_c_229_n N_13_c_381_n 3.931e-19 $X=0.27 $Y=0.232 $X2=0.189 $Y2=0.135
cc_182 N_9_c_239_n N_14_c_386_n 0.00165821f $X=0.27 $Y=0.2025 $X2=0.125
+ $Y2=0.054
cc_183 N_9_c_269_n N_14_c_386_n 0.00263901f $X=0.349 $Y=0.232 $X2=0.125
+ $Y2=0.054
cc_184 N_9_c_270_n N_14_c_386_n 0.00105007f $X=0.324 $Y=0.232 $X2=0.125
+ $Y2=0.054
cc_185 N_9_c_243_n N_14_c_386_n 5.71406e-19 $X=0.324 $Y=0.036 $X2=0.125
+ $Y2=0.054
cc_186 N_9_c_325_p N_14_c_386_n 0.0127725f $X=0.358 $Y=0.223 $X2=0.125 $Y2=0.054
cc_187 N_9_c_254_n N_14_c_386_n 2.57332e-19 $X=0.392 $Y=0.19 $X2=0.125 $Y2=0.054
cc_188 N_9_c_243_n N_15_c_396_n 0.00179714f $X=0.324 $Y=0.036 $X2=0.189
+ $Y2=0.135
cc_189 N_9_c_328_p N_15_c_396_n 0.00159984f $X=0.392 $Y=0.036 $X2=0.189
+ $Y2=0.135
cc_190 N_9_c_329_p N_15_c_396_n 4.19603e-19 $X=0.358 $Y=0.036 $X2=0.189
+ $Y2=0.135
cc_191 N_9_c_258_n N_16_M9_d 5.62141e-19 $X=0.742 $Y=0.108 $X2=0.189 $Y2=0.0675
cc_192 N_9_c_331_p N_17_M11_s 4.38445e-19 $X=0.828 $Y=0.108 $X2=0.189 $Y2=0.0675
cc_193 N_10_c_357_p N_GCLK_c_365_n 0.00134945f $X=0.891 $Y=0.1675 $X2=0 $Y2=0
cc_194 N_10_M12_g N_GCLK_c_366_n 2.25273e-19 $X=0.891 $Y=0.0675 $X2=0.351
+ $Y2=0.1335
cc_195 N_10_c_359_p N_GCLK_c_366_n 0.0022432f $X=0.882 $Y=0.072 $X2=0.351
+ $Y2=0.1335
cc_196 N_10_c_359_p N_GCLK_c_368_n 0.00137679f $X=0.882 $Y=0.072 $X2=0.621
+ $Y2=0.0675
cc_197 N_10_c_356_n N_GCLK_c_369_n 3.33464e-19 $X=0.837 $Y=0.228 $X2=0.621
+ $Y2=0.135
cc_198 N_10_c_353_n GCLK 0.00272952f $X=0.891 $Y=0.136 $X2=0.729 $Y2=0.162
cc_199 N_10_c_359_p N_GCLK_c_371_n 0.00272952f $X=0.882 $Y=0.072 $X2=0.729
+ $Y2=0.216
cc_200 N_10_c_340_n N_17_M11_s 4.99504e-19 $X=0.846 $Y=0.072 $X2=0.243
+ $Y2=0.1335
cc_201 N_12_c_372_n N_13_c_381_n 9.62374e-19 $X=0.272 $Y=0.0675 $X2=0.189
+ $Y2=0.135

* END of "./ICGx1_ASAP7_75t_SRAM.pex.sp.ICGX1_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: ICGx2_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:32:00 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "ICGx2_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./ICGx2_ASAP7_75t_SRAM.pex.sp.pex"
* File: ICGx2_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:32:00 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_ICGX2_ASAP7_75T_SRAM%ENA 2 5 7 12 14 VSS
c8 14 VSS 0.00202376f $X=0.081 $Y=0.137
c9 12 VSS 0.00719777f $X=0.082 $Y=0.125
c10 5 VSS 0.002666f $X=0.081 $Y=0.135
c11 2 VSS 0.0610973f $X=0.081 $Y=0.054
r12 12 14 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.125 $X2=0.081 $Y2=0.137
r13 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.137 $X2=0.081
+ $Y2=0.137
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%SE 2 5 7 10 VSS
c11 10 VSS 0.00136133f $X=0.135 $Y=0.125
c12 5 VSS 0.00157649f $X=0.135 $Y=0.135
c13 2 VSS 0.056849f $X=0.135 $Y=0.054
r14 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.125 $X2=0.135 $Y2=0.137
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.137 $X2=0.135
+ $Y2=0.137
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%5 2 5 7 9 10 13 14 17 19 24 26 28 36 40 44 45 46 47
+ 49 VSS
c23 51 VSS 3.08662e-19 $X=0.189 $Y=0.206
c24 49 VSS 9.26001e-20 $X=0.189 $Y=0.198
c25 47 VSS 3.45068e-20 $X=0.189 $Y=0.127
c26 46 VSS 6.5293e-19 $X=0.189 $Y=0.119
c27 45 VSS 4.30607e-19 $X=0.189 $Y=0.09
c28 44 VSS 2.54814e-19 $X=0.189 $Y=0.076
c29 43 VSS 5.02744e-19 $X=0.189 $Y=0.072
c30 40 VSS 8.26035e-19 $X=0.189 $Y=0.135
c31 36 VSS 0.00146362f $X=0.144 $Y=0.036
c32 35 VSS 0.00266146f $X=0.126 $Y=0.036
c33 30 VSS 0.00201059f $X=0.108 $Y=0.036
c34 28 VSS 0.00804964f $X=0.18 $Y=0.036
c35 27 VSS 0.00324205f $X=0.162 $Y=0.233
c36 26 VSS 0.00135162f $X=0.144 $Y=0.233
c37 25 VSS 0.003458f $X=0.126 $Y=0.233
c38 24 VSS 0.00525509f $X=0.09 $Y=0.233
c39 19 VSS 0.00468477f $X=0.18 $Y=0.233
c40 17 VSS 0.00188709f $X=0.056 $Y=0.216
c41 14 VSS 4.96055e-19 $X=0.071 $Y=0.216
c42 13 VSS 0.00796456f $X=0.108 $Y=0.054
c43 9 VSS 5.3314e-19 $X=0.125 $Y=0.054
c44 5 VSS 0.00138612f $X=0.189 $Y=0.135
c45 2 VSS 0.0577976f $X=0.189 $Y=0.0675
r46 52 53 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.223 $X2=0.189 $Y2=0.2235
r47 51 52 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.206 $X2=0.189 $Y2=0.223
r48 50 51 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.199 $X2=0.189 $Y2=0.206
r49 49 50 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.198 $X2=0.189 $Y2=0.199
r50 48 49 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.184 $X2=0.189 $Y2=0.198
r51 46 47 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.119 $X2=0.189 $Y2=0.127
r52 45 46 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.09 $X2=0.189 $Y2=0.119
r53 44 45 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.076 $X2=0.189 $Y2=0.09
r54 43 44 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.072 $X2=0.189 $Y2=0.076
r55 42 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.063 $X2=0.189 $Y2=0.072
r56 40 48 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.184
r57 40 47 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.127
r58 38 53 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.224 $X2=0.189 $Y2=0.2235
r59 37 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r60 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r61 30 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r62 28 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r63 28 36 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.144 $Y2=0.036
r64 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.233 $X2=0.162 $Y2=0.233
r65 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.233 $X2=0.144 $Y2=0.233
r66 24 25 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.233 $X2=0.126 $Y2=0.233
r67 21 24 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.233 $X2=0.09 $Y2=0.233
r68 19 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.233 $X2=0.189 $Y2=0.224
r69 19 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.233 $X2=0.162 $Y2=0.233
r70 17 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.233 $X2=0.054
+ $Y2=0.233
r71 14 17 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r72 13 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r73 10 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.054 $X2=0.108 $Y2=0.054
r74 9 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.054 $X2=0.108 $Y2=0.054
r75 5 40 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r76 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r77 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%CLK 2 5 8 14 17 19 22 27 30 33 35 40 42 45 47 48 49
+ 52 65 66 69 70 71 75 80 91 92 VSS
c90 102 VSS 1.751e-20 $X=0.621 $Y=0.15
c91 92 VSS 6.23569e-19 $X=0.405 $Y=0.134
c92 91 VSS 0.00814038f $X=0.405 $Y=0.134
c93 80 VSS 2.48826e-19 $X=0.621 $Y=0.133
c94 75 VSS 9.46764e-19 $X=0.243 $Y=0.133
c95 71 VSS 6.07691e-19 $X=0.6015 $Y=0.153
c96 70 VSS 0.00403965f $X=0.582 $Y=0.153
c97 69 VSS 0.00101808f $X=0.621 $Y=0.153
c98 68 VSS 0.00158411f $X=0.621 $Y=0.153
c99 66 VSS 0.00143958f $X=0.3595 $Y=0.153
c100 65 VSS 0.00275092f $X=0.296 $Y=0.153
c101 52 VSS 0.00127303f $X=0.756 $Y=0.162
c102 49 VSS 1.21131e-19 $X=0.6935 $Y=0.187
c103 48 VSS 1.74568e-19 $X=0.688 $Y=0.187
c104 47 VSS 4.53034e-19 $X=0.684 $Y=0.187
c105 46 VSS 0.00441397f $X=0.666 $Y=0.187
c106 43 VSS 9.76836e-19 $X=0.63 $Y=0.187
c107 42 VSS 0.00283826f $X=0.747 $Y=0.187
c108 40 VSS 6.61017e-19 $X=0.3555 $Y=0.1335
c109 33 VSS 0.00699063f $X=0.783 $Y=0.162
c110 30 VSS 0.0600574f $X=0.783 $Y=0.0675
c111 22 VSS 0.0600791f $X=0.729 $Y=0.0675
c112 17 VSS 0.00236251f $X=0.621 $Y=0.135
c113 14 VSS 0.0620989f $X=0.621 $Y=0.0675
c114 8 VSS 0.0605267f $X=0.351 $Y=0.0405
c115 2 VSS 0.0605313f $X=0.243 $Y=0.1335
r116 101 102 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.147 $X2=0.621 $Y2=0.15
r117 91 92 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.405 $Y=0.134
+ $X2=0.405 $Y2=0.134
r118 80 101 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.133 $X2=0.621 $Y2=0.147
r119 70 71 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.582
+ $Y=0.153 $X2=0.6015 $Y2=0.153
r120 69 102 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.621 $Y2=0.15
r121 68 71 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.6015 $Y2=0.153
r122 68 69 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.621 $Y=0.153 $X2=0.621
+ $Y2=0.153
r123 65 66 4.31173 $w=1.8e-08 $l=6.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.296
+ $Y=0.153 $X2=0.3595 $Y2=0.153
r124 64 92 0.725694 $w=3.2e-08 $l=3.36861e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4305 $Y=0.153 $X2=0.405 $Y2=0.134
r125 63 70 10.7963 $w=1.8e-08 $l=1.59e-07 $layer=M2 $thickness=3.6e-08 $X=0.423
+ $Y=0.153 $X2=0.582 $Y2=0.153
r126 63 66 4.31173 $w=1.8e-08 $l=6.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.423
+ $Y=0.153 $X2=0.3595 $Y2=0.153
r127 63 64 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.423 $Y=0.153 $X2=0.423
+ $Y2=0.153
r128 60 75 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.133
r129 59 65 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.296 $Y2=0.153
r130 59 60 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.153 $X2=0.243
+ $Y2=0.153
r131 57 69 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.178 $X2=0.621 $Y2=0.153
r132 52 53 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.756 $Y=0.162 $X2=0.756
+ $Y2=0.162
r133 50 52 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.178 $X2=0.756 $Y2=0.162
r134 48 49 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.187 $X2=0.6935 $Y2=0.187
r135 47 48 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.187 $X2=0.688 $Y2=0.187
r136 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.187 $X2=0.684 $Y2=0.187
r137 45 49 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.699
+ $Y=0.187 $X2=0.6935 $Y2=0.187
r138 43 57 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.63 $Y=0.187 $X2=0.621 $Y2=0.178
r139 43 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.187 $X2=0.666 $Y2=0.187
r140 42 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.747 $Y=0.187 $X2=0.756 $Y2=0.178
r141 42 45 3.25926 $w=1.8e-08 $l=4.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.187 $X2=0.699 $Y2=0.187
r142 40 91 41.0143 $w=2.5e-08 $l=4.95e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.3555 $Y=0.1335 $X2=0.405 $Y2=0.1335
r143 33 53 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.783
+ $Y=0.162 $X2=0.756 $Y2=0.162
r144 33 35 202.311 $w=2e-08 $l=5.4e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.162 $X2=0.783 $Y2=0.216
r145 30 33 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.162
r146 25 53 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.162 $X2=0.756 $Y2=0.162
r147 25 27 202.311 $w=2e-08 $l=5.4e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.162 $X2=0.729 $Y2=0.216
r148 22 25 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.162
r149 17 80 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.133 $X2=0.621
+ $Y2=0.133
r150 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2025
r151 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r152 11 40 4.28571 $w=2.1e-08 $l=4.5e-09 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.1335 $X2=0.3555 $Y2=0.1335
r153 8 11 348.425 $w=2e-08 $l=9.3e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0405 $X2=0.351 $Y2=0.1335
r154 2 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.133 $X2=0.243
+ $Y2=0.133
r155 2 5 258.509 $w=2e-08 $l=6.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1335 $X2=0.243 $Y2=0.2025
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%7 2 5 7 9 12 14 17 22 32 34 35 41 43 48 51 52 64 65
+ 67 71 VSS
c61 72 VSS 2.26979e-19 $X=0.308 $Y=0.189
c62 71 VSS 4.78866e-20 $X=0.306 $Y=0.189
c63 67 VSS 4.14661e-19 $X=0.568 $Y=0.222
c64 65 VSS 8.31219e-19 $X=0.568 $Y=0.1525
c65 64 VSS 3.2551e-19 $X=0.568 $Y=0.116
c66 52 VSS 7.99983e-19 $X=0.568 $Y=0.189
c67 51 VSS 0.00784196f $X=0.568 $Y=0.189
c68 48 VSS 7.00345e-19 $X=0.31 $Y=0.189
c69 44 VSS 8.31083e-19 $X=0.5855 $Y=0.232
c70 43 VSS 0.00225204f $X=0.577 $Y=0.232
c71 41 VSS 0.00296213f $X=0.594 $Y=0.232
c72 35 VSS 1.60717e-19 $X=0.5855 $Y=0.086
c73 34 VSS 2.76555e-19 $X=0.577 $Y=0.086
c74 32 VSS 6.35967e-19 $X=0.594 $Y=0.086
c75 22 VSS 0.00293691f $X=0.297 $Y=0.133
c76 17 VSS 0.00522363f $X=0.596 $Y=0.2025
c77 14 VSS 4.06194e-19 $X=0.611 $Y=0.2025
c78 12 VSS 0.006146f $X=0.596 $Y=0.0675
c79 9 VSS 3.3425e-19 $X=0.611 $Y=0.0675
c80 5 VSS 0.00108474f $X=0.297 $Y=0.1335
c81 2 VSS 0.0591582f $X=0.297 $Y=0.0675
r82 71 72 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.189 $X2=0.308 $Y2=0.189
r83 68 71 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.306 $Y2=0.189
r84 66 67 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.196 $X2=0.568 $Y2=0.222
r85 64 65 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.116 $X2=0.568 $Y2=0.1525
r86 52 66 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.189 $X2=0.568 $Y2=0.196
r87 52 65 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.189 $X2=0.568 $Y2=0.1525
r88 51 52 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.568 $Y=0.189 $X2=0.568
+ $Y2=0.189
r89 48 72 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.31
+ $Y=0.189 $X2=0.308 $Y2=0.189
r90 47 51 17.5185 $w=1.8e-08 $l=2.58e-07 $layer=M2 $thickness=3.6e-08 $X=0.31
+ $Y=0.189 $X2=0.568 $Y2=0.189
r91 47 48 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.31 $Y=0.189 $X2=0.31
+ $Y2=0.189
r92 43 44 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.577
+ $Y=0.232 $X2=0.5855 $Y2=0.232
r93 41 44 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.232 $X2=0.5855 $Y2=0.232
r94 38 67 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.223 $X2=0.568 $Y2=0.222
r95 37 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.232 $X2=0.577 $Y2=0.232
r96 37 38 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.232 $X2=0.568 $Y2=0.223
r97 34 35 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.577
+ $Y=0.086 $X2=0.5855 $Y2=0.086
r98 32 35 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.086 $X2=0.5855 $Y2=0.086
r99 29 64 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.095 $X2=0.568 $Y2=0.116
r100 28 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.086 $X2=0.577 $Y2=0.086
r101 28 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.086 $X2=0.568 $Y2=0.095
r102 20 68 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.18 $X2=0.297 $Y2=0.189
r103 20 22 3.19136 $w=1.8e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.18 $X2=0.297 $Y2=0.133
r104 17 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.232
+ $X2=0.594 $Y2=0.232
r105 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2025 $X2=0.596 $Y2=0.2025
r106 12 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.086
+ $X2=0.594 $Y2=0.086
r107 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0675 $X2=0.596 $Y2=0.0675
r108 5 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.133 $X2=0.297
+ $Y2=0.133
r109 5 7 359.664 $w=2e-08 $l=9.6e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.1335 $X2=0.297 $Y2=0.2295
r110 2 5 247.269 $w=2e-08 $l=6.6e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.1335
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%8 2 5 7 9 12 14 17 19 21 30 31 34 35 36 37 38 39 40
+ 42 VSS
c35 48 VSS 0.00202496f $X=0.503 $Y=0.233
c36 47 VSS 0.00196262f $X=0.5125 $Y=0.233
c37 42 VSS 0.00220406f $X=0.486 $Y=0.233
c38 40 VSS 4.74628e-19 $X=0.5125 $Y=0.2115
c39 39 VSS 4.02544e-19 $X=0.5125 $Y=0.199
c40 38 VSS 0.00108412f $X=0.5125 $Y=0.181
c41 37 VSS 3.28082e-19 $X=0.5125 $Y=0.162
c42 36 VSS 7.74522e-19 $X=0.5125 $Y=0.144
c43 35 VSS 6.76213e-19 $X=0.5125 $Y=0.12
c44 34 VSS 7.4117e-19 $X=0.5125 $Y=0.224
c45 32 VSS 2.34081e-20 $X=0.4795 $Y=0.082
c46 31 VSS 3.47256e-19 $X=0.473 $Y=0.082
c47 30 VSS 5.61168e-19 $X=0.447 $Y=0.082
c48 29 VSS 1.3164e-20 $X=0.414 $Y=0.082
c49 21 VSS 3.43763e-19 $X=0.406 $Y=0.082
c50 19 VSS 6.74711e-19 $X=0.503 $Y=0.082
c51 17 VSS 0.0029927f $X=0.484 $Y=0.2295
c52 12 VSS 0.0170022f $X=0.484 $Y=0.0405
c53 5 VSS 0.00244059f $X=0.405 $Y=0.082
c54 2 VSS 0.058916f $X=0.405 $Y=0.0405
r55 48 49 0.322531 $w=1.8e-08 $l=4.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.503
+ $Y=0.233 $X2=0.50775 $Y2=0.233
r56 47 49 0.322531 $w=1.8e-08 $l=4.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.233 $X2=0.50775 $Y2=0.233
r57 42 48 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.233 $X2=0.503 $Y2=0.233
r58 39 40 0.793941 $w=1.9e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.199 $X2=0.5125 $Y2=0.2115
r59 38 39 1.14327 $w=1.9e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.181 $X2=0.5125 $Y2=0.199
r60 37 38 1.20679 $w=1.9e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.162 $X2=0.5125 $Y2=0.181
r61 36 37 1.14327 $w=1.9e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.144 $X2=0.5125 $Y2=0.162
r62 35 36 1.52437 $w=1.9e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.12 $X2=0.5125 $Y2=0.144
r63 34 47 0.0384781 $w=1.9e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.224 $X2=0.5125 $Y2=0.233
r64 34 40 0.793941 $w=1.9e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.224 $X2=0.5125 $Y2=0.2115
r65 33 35 1.84194 $w=1.9e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.091 $X2=0.5125 $Y2=0.12
r66 31 32 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.473
+ $Y=0.082 $X2=0.4795 $Y2=0.082
r67 30 31 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.082 $X2=0.473 $Y2=0.082
r68 29 30 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.082 $X2=0.447 $Y2=0.082
r69 27 32 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.082 $X2=0.4795 $Y2=0.082
r70 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.082 $X2=0.486
+ $Y2=0.082
r71 21 29 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.406
+ $Y=0.082 $X2=0.414 $Y2=0.082
r72 19 33 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.503 $Y=0.082 $X2=0.5125 $Y2=0.091
r73 19 27 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.503
+ $Y=0.082 $X2=0.486 $Y2=0.082
r74 17 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.233 $X2=0.486
+ $Y2=0.233
r75 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2295 $X2=0.484 $Y2=0.2295
r76 12 28 35.8185 $w=2.4e-08 $l=4.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0405 $X2=0.486 $Y2=0.082
r77 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0405 $X2=0.484 $Y2=0.0405
r78 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.406 $Y=0.082 $X2=0.406
+ $Y2=0.082
r79 5 7 552.609 $w=2e-08 $l=1.475e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.082 $X2=0.405 $Y2=0.2295
r80 2 5 155.48 $w=2e-08 $l=4.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0405 $X2=0.405 $Y2=0.082
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%9 2 5 7 10 13 15 18 21 23 25 30 33 37 38 41 43 49
+ 50 53 58 59 60 61 62 64 65 67 68 69 70 72 75 77 79 86 88 89 90 91 93 94 95 96
+ 97 98 101 107 110 VSS
c104 113 VSS 8.63727e-20 $X=0.837 $Y=0.125
c105 110 VSS 3.89134e-19 $X=0.837 $Y=0.133
c106 107 VSS 3.25689e-19 $X=0.837 $Y=0.108
c107 101 VSS 6.17137e-19 $X=0.675 $Y=0.133
c108 99 VSS 4.28973e-19 $X=0.675 $Y=0.108
c109 98 VSS 1.77849e-19 $X=0.358 $Y=0.19
c110 97 VSS 0.00171031f $X=0.358 $Y=0.036
c111 96 VSS 3.16771e-19 $X=0.7965 $Y=0.108
c112 95 VSS 2.5364e-19 $X=0.765 $Y=0.108
c113 94 VSS 7.79718e-20 $X=0.747 $Y=0.108
c114 93 VSS 0.00155044f $X=0.742 $Y=0.108
c115 91 VSS 6.48597e-19 $X=0.828 $Y=0.108
c116 90 VSS 8.07734e-20 $X=0.675 $Y=0.097
c117 89 VSS 4.90266e-19 $X=0.675 $Y=0.095
c118 88 VSS 1.49364e-19 $X=0.675 $Y=0.081
c119 87 VSS 1.86503e-19 $X=0.675 $Y=0.077
c120 86 VSS 5.68609e-19 $X=0.675 $Y=0.073
c121 85 VSS 8.45284e-19 $X=0.675 $Y=0.063
c122 84 VSS 6.05801e-20 $X=0.675 $Y=0.099
c123 80 VSS 5.02745e-19 $X=0.453 $Y=0.19
c124 79 VSS 0.00172533f $X=0.447 $Y=0.19
c125 78 VSS 3.27114e-19 $X=0.396 $Y=0.19
c126 77 VSS 0.00110887f $X=0.392 $Y=0.19
c127 75 VSS 8.20031e-19 $X=0.459 $Y=0.19
c128 72 VSS 0.00146505f $X=0.63 $Y=0.036
c129 71 VSS 2.9457e-19 $X=0.612 $Y=0.036
c130 70 VSS 0.00428093f $X=0.609 $Y=0.036
c131 69 VSS 0.00316044f $X=0.559 $Y=0.036
c132 68 VSS 0.0128572f $X=0.522 $Y=0.036
c133 67 VSS 0.00218374f $X=0.392 $Y=0.036
c134 65 VSS 0.0076085f $X=0.666 $Y=0.036
c135 64 VSS 7.19963e-19 $X=0.358 $Y=0.223
c136 62 VSS 3.15222e-19 $X=0.358 $Y=0.18
c137 61 VSS 3.80467e-19 $X=0.358 $Y=0.162
c138 60 VSS 5.42963e-19 $X=0.358 $Y=0.12
c139 59 VSS 2.16018e-19 $X=0.358 $Y=0.091
c140 57 VSS 5.84318e-19 $X=0.358 $Y=0.072
c141 53 VSS 0.00229455f $X=0.324 $Y=0.036
c142 50 VSS 0.00436152f $X=0.349 $Y=0.036
c143 49 VSS 0.00260946f $X=0.324 $Y=0.232
c144 48 VSS 0.00204527f $X=0.288 $Y=0.232
c145 43 VSS 0.00103077f $X=0.27 $Y=0.232
c146 41 VSS 0.00444971f $X=0.349 $Y=0.232
c147 40 VSS 6.58864e-19 $X=0.27 $Y=0.2295
c148 37 VSS 0.00129546f $X=0.27 $Y=0.2025
c149 32 VSS 5.70081e-19 $X=0.324 $Y=0.0405
c150 21 VSS 0.00210626f $X=0.837 $Y=0.135
c151 18 VSS 0.0569001f $X=0.837 $Y=0.0675
c152 13 VSS 0.00240787f $X=0.675 $Y=0.135
c153 10 VSS 0.0575264f $X=0.675 $Y=0.0675
c154 5 VSS 0.00191265f $X=0.459 $Y=0.19
c155 2 VSS 0.0630025f $X=0.459 $Y=0.0405
r156 112 113 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.117 $X2=0.837 $Y2=0.125
r157 110 113 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.133 $X2=0.837 $Y2=0.125
r158 107 112 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.108 $X2=0.837 $Y2=0.117
r159 103 104 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.116 $X2=0.675 $Y2=0.117
r160 101 104 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.133 $X2=0.675 $Y2=0.117
r161 99 103 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.108 $X2=0.675 $Y2=0.116
r162 95 96 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.765
+ $Y=0.108 $X2=0.7965 $Y2=0.108
r163 94 95 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.108 $X2=0.765 $Y2=0.108
r164 93 94 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.742
+ $Y=0.108 $X2=0.747 $Y2=0.108
r165 92 99 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.108 $X2=0.675 $Y2=0.108
r166 92 93 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.108 $X2=0.742 $Y2=0.108
r167 91 107 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.108 $X2=0.837 $Y2=0.108
r168 91 96 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.108 $X2=0.7965 $Y2=0.108
r169 89 90 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.095 $X2=0.675 $Y2=0.097
r170 88 89 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.081 $X2=0.675 $Y2=0.095
r171 87 88 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.077 $X2=0.675 $Y2=0.081
r172 86 87 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.073 $X2=0.675 $Y2=0.077
r173 85 86 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.063 $X2=0.675 $Y2=0.073
r174 84 99 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.099 $X2=0.675 $Y2=0.108
r175 84 90 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.099 $X2=0.675 $Y2=0.097
r176 83 85 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.045 $X2=0.675 $Y2=0.063
r177 79 80 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.19 $X2=0.453 $Y2=0.19
r178 78 79 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.19 $X2=0.447 $Y2=0.19
r179 77 78 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.392
+ $Y=0.19 $X2=0.396 $Y2=0.19
r180 75 80 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.19 $X2=0.453 $Y2=0.19
r181 73 98 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.19 $X2=0.358 $Y2=0.19
r182 73 77 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.19 $X2=0.392 $Y2=0.19
r183 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.63 $Y2=0.036
r184 70 71 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.609
+ $Y=0.036 $X2=0.612 $Y2=0.036
r185 69 70 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.559
+ $Y=0.036 $X2=0.609 $Y2=0.036
r186 68 69 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.559 $Y2=0.036
r187 67 68 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.392
+ $Y=0.036 $X2=0.522 $Y2=0.036
r188 66 97 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.036 $X2=0.358 $Y2=0.036
r189 66 67 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.036 $X2=0.392 $Y2=0.036
r190 65 83 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.036 $X2=0.675 $Y2=0.045
r191 65 72 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.63 $Y2=0.036
r192 63 98 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.199 $X2=0.358 $Y2=0.19
r193 63 64 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.199 $X2=0.358 $Y2=0.223
r194 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.162 $X2=0.358 $Y2=0.18
r195 60 61 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.12 $X2=0.358 $Y2=0.162
r196 59 60 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.091 $X2=0.358 $Y2=0.12
r197 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.073 $X2=0.358 $Y2=0.091
r198 57 58 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.072 $X2=0.358 $Y2=0.073
r199 56 98 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.181 $X2=0.358 $Y2=0.19
r200 56 62 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.181 $X2=0.358 $Y2=0.18
r201 55 97 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.045 $X2=0.358 $Y2=0.036
r202 55 57 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.045 $X2=0.358 $Y2=0.072
r203 52 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r204 50 97 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.349
+ $Y=0.036 $X2=0.358 $Y2=0.036
r205 50 52 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.349
+ $Y=0.036 $X2=0.324 $Y2=0.036
r206 48 49 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.232 $X2=0.324 $Y2=0.232
r207 43 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.232 $X2=0.288 $Y2=0.232
r208 41 64 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.349 $Y=0.232 $X2=0.358 $Y2=0.223
r209 41 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.349
+ $Y=0.232 $X2=0.324 $Y2=0.232
r210 38 40 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2295 $X2=0.27 $Y2=0.2295
r211 37 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.232 $X2=0.27
+ $Y2=0.232
r212 34 40 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2655 $Y=0.216 $X2=0.27 $Y2=0.2295
r213 34 37 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2655 $Y=0.216 $X2=0.2655 $Y2=0.189
r214 33 37 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.189 $X2=0.2655 $Y2=0.189
r215 30 32 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0405 $X2=0.324 $Y2=0.0405
r216 29 53 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r217 26 32 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.054 $X2=0.324 $Y2=0.0405
r218 26 29 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.054 $X2=0.3195 $Y2=0.081
r219 25 29 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.081 $X2=0.3195 $Y2=0.081
r220 21 110 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.133
+ $X2=0.837 $Y2=0.133
r221 21 23 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.216
r222 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0675 $X2=0.837 $Y2=0.135
r223 13 101 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.133
+ $X2=0.675 $Y2=0.133
r224 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.216
r225 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0675 $X2=0.675 $Y2=0.135
r226 5 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.19 $X2=0.459
+ $Y2=0.19
r227 5 7 147.987 $w=2e-08 $l=3.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.19 $X2=0.459 $Y2=0.2295
r228 2 5 560.102 $w=2e-08 $l=1.495e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0405 $X2=0.459 $Y2=0.19
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%10 2 7 10 13 15 17 18 21 22 23 26 27 28 40 41 42 47
+ 54 57 59 60 68 VSS
c43 68 VSS 0.00355073f $X=0.837 $Y=0.228
c44 67 VSS 1.56305e-19 $X=0.837 $Y=0.225
c45 66 VSS 7.65866e-19 $X=0.837 $Y=0.222
c46 64 VSS 0.00240875f $X=0.837 $Y=0.231
c47 60 VSS 4.03714e-19 $X=0.837 $Y=0.197
c48 59 VSS 5.64067e-19 $X=0.891 $Y=0.1675
c49 57 VSS 3.61137e-19 $X=0.891 $Y=0.1175
c50 54 VSS 2.06442e-19 $X=0.891 $Y=0.136
c51 52 VSS 2.2993e-19 $X=0.891 $Y=0.188
c52 49 VSS 0.00388157f $X=0.882 $Y=0.197
c53 48 VSS 0.00379396f $X=0.879 $Y=0.072
c54 47 VSS 0.00352836f $X=0.846 $Y=0.072
c55 42 VSS 6.46932e-20 $X=0.882 $Y=0.072
c56 41 VSS 0.00231927f $X=0.7875 $Y=0.231
c57 40 VSS 0.00805297f $X=0.765 $Y=0.231
c58 31 VSS 0.00656665f $X=0.81 $Y=0.216
c59 27 VSS 6.59309e-19 $X=0.827 $Y=0.216
c60 26 VSS 0.0060288f $X=0.702 $Y=0.216
c61 22 VSS 7.72153e-19 $X=0.719 $Y=0.216
c62 21 VSS 0.004367f $X=0.756 $Y=0.0675
c63 17 VSS 7.90436e-19 $X=0.773 $Y=0.0675
c64 13 VSS 0.00379511f $X=0.945 $Y=0.136
c65 10 VSS 0.0615048f $X=0.945 $Y=0.0675
c66 2 VSS 0.0580673f $X=0.891 $Y=0.0675
r67 67 68 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.228
r68 66 67 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.222 $X2=0.837 $Y2=0.225
r69 65 66 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.206 $X2=0.837 $Y2=0.222
r70 64 68 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.231 $X2=0.837 $Y2=0.228
r71 60 65 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.197 $X2=0.837 $Y2=0.206
r72 58 59 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.147 $X2=0.891 $Y2=0.1675
r73 56 57 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.099 $X2=0.891 $Y2=0.1175
r74 54 58 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.136 $X2=0.891 $Y2=0.147
r75 54 57 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.136 $X2=0.891 $Y2=0.1175
r76 52 59 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.188 $X2=0.891 $Y2=0.1675
r77 51 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.081 $X2=0.891 $Y2=0.099
r78 50 60 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.197 $X2=0.837 $Y2=0.197
r79 49 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.197 $X2=0.891 $Y2=0.188
r80 49 50 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.197 $X2=0.846 $Y2=0.197
r81 47 48 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.072 $X2=0.879 $Y2=0.072
r82 44 47 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.072 $X2=0.846 $Y2=0.072
r83 42 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.072 $X2=0.891 $Y2=0.081
r84 42 48 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.072 $X2=0.879 $Y2=0.072
r85 40 41 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.765
+ $Y=0.231 $X2=0.7875 $Y2=0.231
r86 38 41 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.231 $X2=0.7875 $Y2=0.231
r87 34 40 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.231 $X2=0.765 $Y2=0.231
r88 32 64 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.231 $X2=0.837 $Y2=0.231
r89 32 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.231 $X2=0.81 $Y2=0.231
r90 31 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.231 $X2=0.81
+ $Y2=0.231
r91 28 31 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.216 $X2=0.81 $Y2=0.216
r92 27 31 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.216 $X2=0.81 $Y2=0.216
r93 26 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.231 $X2=0.702
+ $Y2=0.231
r94 23 26 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.216 $X2=0.702 $Y2=0.216
r95 22 26 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.216 $X2=0.702 $Y2=0.216
r96 21 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.072 $X2=0.756
+ $Y2=0.072
r97 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.756 $Y2=0.0675
r98 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.756 $Y2=0.0675
r99 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.945
+ $Y=0.136 $X2=0.945 $Y2=0.2025
r100 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.0675 $X2=0.945 $Y2=0.136
r101 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.891
+ $Y=0.136 $X2=0.945 $Y2=0.136
r102 5 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.136 $X2=0.891
+ $Y2=0.136
r103 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.136 $X2=0.891 $Y2=0.2025
r104 2 5 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.0675 $X2=0.891 $Y2=0.136
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%GCLK 1 2 6 7 10 11 13 14 18 20 28 30 VSS
c16 32 VSS 4.59291e-19 $X=0.999 $Y=0.2155
c17 30 VSS 0.00281393f $X=0.999 $Y=0.1145
c18 29 VSS 8.85605e-19 $X=0.999 $Y=0.063
c19 28 VSS 0.00474646f $X=1 $Y=0.166
c20 26 VSS 4.55454e-19 $X=0.999 $Y=0.225
c21 20 VSS 0.00191539f $X=0.918 $Y=0.234
c22 18 VSS 0.0131673f $X=0.99 $Y=0.234
c23 14 VSS 0.0103019f $X=0.918 $Y=0.036
c24 13 VSS 0.00398627f $X=0.918 $Y=0.036
c25 11 VSS 0.0131334f $X=0.99 $Y=0.036
c26 10 VSS 0.0103762f $X=0.918 $Y=0.2025
c27 6 VSS 5.38922e-19 $X=0.935 $Y=0.2025
c28 1 VSS 5.38922e-19 $X=0.935 $Y=0.0675
r29 31 32 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.206 $X2=0.999 $Y2=0.2155
r30 29 30 3.49691 $w=1.8e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.063 $X2=0.999 $Y2=0.1145
r31 28 31 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.166 $X2=0.999 $Y2=0.206
r32 28 30 3.49691 $w=1.8e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.166 $X2=0.999 $Y2=0.1145
r33 26 32 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.225 $X2=0.999 $Y2=0.2155
r34 25 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.045 $X2=0.999 $Y2=0.063
r35 18 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.99 $Y=0.234 $X2=0.999 $Y2=0.225
r36 18 20 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.99
+ $Y=0.234 $X2=0.918 $Y2=0.234
r37 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.036 $X2=0.918
+ $Y2=0.036
r38 11 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.99 $Y=0.036 $X2=0.999 $Y2=0.045
r39 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.99
+ $Y=0.036 $X2=0.918 $Y2=0.036
r40 10 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.234 $X2=0.918
+ $Y2=0.234
r41 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.2025 $X2=0.918 $Y2=0.2025
r42 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.935 $Y=0.2025 $X2=0.918 $Y2=0.2025
r43 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.918
+ $Y=0.0675 $X2=0.918 $Y2=0.036
r44 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.901
+ $Y=0.0675 $X2=0.918 $Y2=0.0675
r45 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.935
+ $Y=0.0675 $X2=0.918 $Y2=0.0675
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%12 1 6 9 VSS
c9 9 VSS 0.0194635f $X=0.272 $Y=0.0675
c10 6 VSS 3.61939e-19 $X=0.287 $Y=0.0675
c11 4 VSS 3.25039e-19 $X=0.214 $Y=0.0675
r12 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.272 $Y2=0.0675
r13 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.214
+ $Y=0.0675 $X2=0.272 $Y2=0.0675
r14 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.214 $Y2=0.0675
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%13 1 2 5 VSS
c5 5 VSS 0.00582405f $X=0.216 $Y=0.2025
c6 1 VSS 6.50078e-19 $X=0.233 $Y=0.2025
r7 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.2025 $X2=0.216 $Y2=0.2025
r8 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.216 $Y2=0.2025
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%14 1 6 9 VSS
c10 9 VSS 0.0186419f $X=0.38 $Y=0.2295
c11 6 VSS 3.72954e-19 $X=0.395 $Y=0.2295
c12 4 VSS 3.77944e-19 $X=0.322 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.2295 $X2=0.38 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.2295 $X2=0.38 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2295 $X2=0.322 $Y2=0.2295
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%15 1 2 5 VSS
c4 5 VSS 0.004225f $X=0.378 $Y=0.0405
c5 1 VSS 6.8236e-19 $X=0.395 $Y=0.0405
r6 2 5 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.0405 $X2=0.378 $Y2=0.0405
r7 1 5 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0405 $X2=0.378 $Y2=0.0405
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%16 1 2 VSS
c1 1 VSS 0.00221026f $X=0.719 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0675 $X2=0.685 $Y2=0.0675
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%17 1 2 VSS
c2 1 VSS 0.00230546f $X=0.827 $Y=0.0675
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.827
+ $Y=0.0675 $X2=0.793 $Y2=0.0675
.ends

.subckt PM_ICGX2_ASAP7_75T_SRAM%18 1 2 VSS
c0 1 VSS 0.00242486f $X=0.125 $Y=0.216
r1 1 2 25.1852 $w=5.4e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.216 $X2=0.091 $Y2=0.216
.ends


* END of "./ICGx2_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt ICGx2_ASAP7_75t_SRAM  VSS VDD ENA SE CLK GCLK
* 
* GCLK	GCLK
* CLK	CLK
* SE	SE
* ENA	ENA
M0 N_5_M0_d N_ENA_M0_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 VSS N_SE_M1_g N_5_M1_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 N_12_M2_d N_5_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_9_M3_d N_7_M3_g N_12_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M4 N_15_M4_d N_CLK_M4_g N_9_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.341
+ $Y=0.027
M5 VSS N_8_M5_g N_15_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.395
+ $Y=0.027
M6 N_8_M6_d N_9_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449 $Y=0.027
M7 VSS N_CLK_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M8 VSS N_9_M8_g N_16_M8_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M9 N_16_M9_d N_CLK_M9_g N_10_M9_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M10 N_17_M10_d N_CLK_M10_g N_10_M10_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.773 $Y=0.027
M11 VSS N_9_M11_g N_17_M11_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.027
M12 N_GCLK_M12_d N_10_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.027
M13 N_GCLK_M13_d N_10_M13_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.027
M14 N_18_M14_d N_ENA_M14_g N_5_M14_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.071 $Y=0.189
M15 VDD N_SE_M15_g N_18_M15_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M16 N_13_M16_d N_5_M16_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M17 N_9_M17_d N_CLK_M17_g N_13_M17_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M18 N_14_M18_d N_7_M18_g N_9_M18_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.287 $Y=0.216
M19 VDD N_8_M19_g N_14_M19_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.395
+ $Y=0.216
M20 N_8_M20_d N_9_M20_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.216
M21 VDD N_CLK_M21_g N_7_M21_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M22 N_10_M22_d N_9_M22_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.665
+ $Y=0.189
M23 VDD N_CLK_M23_g N_10_M23_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.719
+ $Y=0.189
M24 VDD N_CLK_M24_g N_10_M24_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.773
+ $Y=0.189
M25 N_10_M25_d N_9_M25_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.827
+ $Y=0.189
M26 N_GCLK_M26_d N_10_M26_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.162
M27 N_GCLK_M27_d N_10_M27_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.162
*
* 
* .include "ICGx2_ASAP7_75t_SRAM.pex.sp.ICGX2_ASAP7_75T_SRAM.pxi"
* BEGIN of "./ICGx2_ASAP7_75t_SRAM.pex.sp.ICGX2_ASAP7_75T_SRAM.pxi"
* File: ICGx2_ASAP7_75t_SRAM.pex.sp.ICGX2_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:32:00 2017
* 
x_PM_ICGX2_ASAP7_75T_SRAM%ENA N_ENA_M0_g N_ENA_c_2_p N_ENA_M14_g ENA N_ENA_c_6_p
+ VSS PM_ICGX2_ASAP7_75T_SRAM%ENA
x_PM_ICGX2_ASAP7_75T_SRAM%SE N_SE_M1_g N_SE_c_10_n N_SE_M15_g SE VSS
+ PM_ICGX2_ASAP7_75T_SRAM%SE
x_PM_ICGX2_ASAP7_75T_SRAM%5 N_5_M2_g N_5_c_26_n N_5_M16_g N_5_M1_s N_5_M0_d
+ N_5_c_21_n N_5_M14_s N_5_c_22_n N_5_c_40_p N_5_c_23_n N_5_c_27_n N_5_c_41_p
+ N_5_c_29_n N_5_c_34_p N_5_c_37_p N_5_c_31_n N_5_c_38_p N_5_c_35_p N_5_c_39_p
+ VSS PM_ICGX2_ASAP7_75T_SRAM%5
x_PM_ICGX2_ASAP7_75T_SRAM%CLK N_CLK_c_43_n N_CLK_M17_g N_CLK_M4_g N_CLK_M7_g
+ N_CLK_c_85_p N_CLK_M21_g N_CLK_M9_g N_CLK_M23_g N_CLK_M10_g N_CLK_c_108_p
+ N_CLK_M24_g N_CLK_c_51_p N_CLK_c_118_p CLK N_CLK_c_84_p N_CLK_c_109_p
+ N_CLK_c_110_p N_CLK_c_111_p N_CLK_c_46_n N_CLK_c_56_p N_CLK_c_53_p
+ N_CLK_c_59_p N_CLK_c_52_p N_CLK_c_47_n N_CLK_c_66_p N_CLK_c_69_p N_CLK_c_62_p
+ VSS PM_ICGX2_ASAP7_75T_SRAM%CLK
x_PM_ICGX2_ASAP7_75T_SRAM%7 N_7_M3_g N_7_c_139_n N_7_M18_g N_7_M7_s N_7_c_141_n
+ N_7_M21_s N_7_c_142_n N_7_c_134_n N_7_c_147_n N_7_c_161_p N_7_c_148_n
+ N_7_c_191_p N_7_c_162_p N_7_c_149_n N_7_c_150_n N_7_c_152_n N_7_c_163_p
+ N_7_c_154_n N_7_c_156_n N_7_c_136_n VSS PM_ICGX2_ASAP7_75T_SRAM%7
x_PM_ICGX2_ASAP7_75T_SRAM%8 N_8_M5_g N_8_c_219_p N_8_M19_g N_8_M6_d N_8_c_197_n
+ N_8_M20_d N_8_c_207_n N_8_c_209_n N_8_c_198_n N_8_c_199_n N_8_c_201_n
+ N_8_c_210_n N_8_c_211_n N_8_c_202_n N_8_c_203_n N_8_c_213_n N_8_c_214_n
+ N_8_c_215_n N_8_c_216_n VSS PM_ICGX2_ASAP7_75T_SRAM%8
x_PM_ICGX2_ASAP7_75T_SRAM%9 N_9_M6_g N_9_c_231_n N_9_M20_g N_9_M8_g N_9_c_236_n
+ N_9_M22_g N_9_M11_g N_9_c_303_p N_9_M25_g N_9_M3_d N_9_M4_s N_9_M17_d
+ N_9_c_239_n N_9_M18_s N_9_c_269_n N_9_c_229_n N_9_c_270_n N_9_c_242_n
+ N_9_c_243_n N_9_c_275_n N_9_c_276_n N_9_c_244_n N_9_c_245_n N_9_c_250_n
+ N_9_c_326_p N_9_c_304_p N_9_c_329_p N_9_c_295_n N_9_c_251_n N_9_c_279_n
+ N_9_c_252_n N_9_c_282_n N_9_c_254_n N_9_c_256_n N_9_c_311_p N_9_c_285_n
+ N_9_c_305_p N_9_c_286_n N_9_c_332_p N_9_c_258_n N_9_c_261_n N_9_c_262_n
+ N_9_c_263_n N_9_c_330_p N_9_c_287_n N_9_c_265_n N_9_c_314_p N_9_c_313_p VSS
+ PM_ICGX2_ASAP7_75T_SRAM%9
x_PM_ICGX2_ASAP7_75T_SRAM%10 N_10_M12_g N_10_M26_g N_10_M13_g N_10_c_345_n
+ N_10_M27_g N_10_M10_s N_10_M9_s N_10_c_334_n N_10_M23_s N_10_M22_d
+ N_10_c_335_n N_10_M25_d N_10_M24_s N_10_c_337_n N_10_c_339_n N_10_c_366_p
+ N_10_c_341_n N_10_c_355_n N_10_c_356_n N_10_c_362_p N_10_c_357_n N_10_c_358_n
+ VSS PM_ICGX2_ASAP7_75T_SRAM%10
x_PM_ICGX2_ASAP7_75T_SRAM%GCLK N_GCLK_M13_d N_GCLK_M12_d N_GCLK_M27_d N_GCLK_M26_d
+ N_GCLK_c_378_n N_GCLK_c_380_n N_GCLK_c_381_n N_GCLK_c_384_n N_GCLK_c_386_n
+ N_GCLK_c_387_n GCLK N_GCLK_c_391_n VSS PM_ICGX2_ASAP7_75T_SRAM%GCLK
x_PM_ICGX2_ASAP7_75T_SRAM%12 N_12_M2_d N_12_M3_s N_12_c_392_n VSS
+ PM_ICGX2_ASAP7_75T_SRAM%12
x_PM_ICGX2_ASAP7_75T_SRAM%13 N_13_M17_s N_13_M16_d N_13_c_401_n VSS
+ PM_ICGX2_ASAP7_75T_SRAM%13
x_PM_ICGX2_ASAP7_75T_SRAM%14 N_14_M18_d N_14_M19_s N_14_c_406_n VSS
+ PM_ICGX2_ASAP7_75T_SRAM%14
x_PM_ICGX2_ASAP7_75T_SRAM%15 N_15_M5_s N_15_M4_d N_15_c_416_n VSS
+ PM_ICGX2_ASAP7_75T_SRAM%15
x_PM_ICGX2_ASAP7_75T_SRAM%16 N_16_M9_d N_16_M8_s VSS PM_ICGX2_ASAP7_75T_SRAM%16
x_PM_ICGX2_ASAP7_75T_SRAM%17 N_17_M11_s N_17_M10_d VSS PM_ICGX2_ASAP7_75T_SRAM%17
x_PM_ICGX2_ASAP7_75T_SRAM%18 N_18_M15_s N_18_M14_d VSS PM_ICGX2_ASAP7_75T_SRAM%18
cc_1 N_ENA_M0_g N_SE_M1_g 0.00328721f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_ENA_c_2_p N_SE_c_10_n 9.35826e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 ENA SE 0.00588002f $X=0.082 $Y=0.125 $X2=0.135 $Y2=0.125
cc_4 N_ENA_M0_g N_5_M2_g 2.13359e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 ENA N_5_c_21_n 6.06976e-19 $X=0.082 $Y=0.125 $X2=0.135 $Y2=0.137
cc_6 N_ENA_c_6_p N_5_c_22_n 0.00176249f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_7 N_ENA_M0_g N_5_c_23_n 2.28086e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_8 N_ENA_c_6_p N_5_c_23_n 0.00499899f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_9 N_SE_M1_g N_5_M2_g 0.00268443f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_10 N_SE_c_10_n N_5_c_26_n 9.11034e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_11 N_SE_M1_g N_5_c_27_n 2.59938e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_12 SE N_5_c_27_n 0.00123553f $X=0.135 $Y=0.125 $X2=0 $Y2=0
cc_13 N_SE_M1_g N_5_c_29_n 2.84283e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_14 SE N_5_c_29_n 0.001038f $X=0.135 $Y=0.125 $X2=0 $Y2=0
cc_15 SE N_5_c_31_n 0.00457266f $X=0.135 $Y=0.125 $X2=0 $Y2=0
cc_16 N_SE_M1_g N_CLK_c_43_n 2.13359e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_17 N_5_M2_g N_CLK_c_43_n 0.00341068f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_18 N_5_c_26_n N_CLK_c_43_n 8.10277e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.054
cc_19 N_5_c_34_p N_CLK_c_46_n 3.51913e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_20 N_5_c_35_p N_CLK_c_47_n 0.00253596f $X=0.189 $Y=0.127 $X2=0 $Y2=0
cc_21 N_5_M2_g N_7_M3_g 2.82885e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_22 N_5_c_37_p N_7_c_134_n 3.23824e-19 $X=0.189 $Y=0.076 $X2=0 $Y2=0
cc_23 N_5_c_38_p N_7_c_134_n 2.18117e-19 $X=0.189 $Y=0.119 $X2=0 $Y2=0
cc_24 N_5_c_39_p N_7_c_136_n 2.18117e-19 $X=0.189 $Y=0.198 $X2=0 $Y2=0
cc_25 N_5_c_40_p N_9_c_229_n 4.49022e-19 $X=0.18 $Y=0.233 $X2=0 $Y2=0
cc_26 N_5_c_41_p N_12_c_392_n 0.00246673f $X=0.18 $Y=0.036 $X2=0 $Y2=0
cc_27 N_5_c_34_p N_13_c_401_n 0.00181721f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_28 N_CLK_c_43_n N_7_M3_g 0.00355599f $X=0.243 $Y=0.1335 $X2=0.135 $Y2=0.054
cc_29 N_CLK_M4_g N_7_M3_g 0.00355599f $X=0.351 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_30 N_CLK_c_43_n N_7_c_139_n 8.50652e-19 $X=0.243 $Y=0.1335 $X2=0.135
+ $Y2=0.135
cc_31 N_CLK_c_51_p N_7_c_139_n 9.47532e-19 $X=0.3555 $Y=0.1335 $X2=0.135
+ $Y2=0.135
cc_32 N_CLK_c_52_p N_7_c_141_n 2.51466e-19 $X=0.6015 $Y=0.153 $X2=0.135
+ $Y2=0.137
cc_33 N_CLK_c_53_p N_7_c_142_n 6.13009e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_34 N_CLK_c_52_p N_7_c_142_n 2.98103e-19 $X=0.6015 $Y=0.153 $X2=0 $Y2=0
cc_35 N_CLK_c_46_n N_7_c_134_n 0.0010183f $X=0.296 $Y=0.153 $X2=0 $Y2=0
cc_36 N_CLK_c_56_p N_7_c_134_n 5.3655e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_37 N_CLK_c_47_n N_7_c_134_n 0.00252905f $X=0.243 $Y=0.133 $X2=0 $Y2=0
cc_38 N_CLK_c_52_p N_7_c_147_n 2.62247e-19 $X=0.6015 $Y=0.153 $X2=0 $Y2=0
cc_39 N_CLK_c_59_p N_7_c_148_n 2.62247e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_40 N_CLK_c_56_p N_7_c_149_n 2.46239e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_41 N_CLK_c_56_p N_7_c_150_n 0.0242262f $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_42 N_CLK_c_62_p N_7_c_150_n 4.84045e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_43 N_CLK_c_53_p N_7_c_152_n 0.0017697f $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_44 N_CLK_c_59_p N_7_c_152_n 4.75571e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_45 N_CLK_c_59_p N_7_c_154_n 4.04804e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_46 N_CLK_c_66_p N_7_c_154_n 0.00167205f $X=0.621 $Y=0.133 $X2=0 $Y2=0
cc_47 N_CLK_c_59_p N_7_c_156_n 2.46239e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_48 N_CLK_M4_g N_8_M5_g 0.00341068f $X=0.351 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_49 N_CLK_c_69_p N_8_M5_g 0.00207156f $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.054
cc_50 N_CLK_c_62_p N_8_M5_g 2.24185e-19 $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.054
cc_51 N_CLK_c_59_p N_8_c_197_n 2.35254e-19 $X=0.582 $Y=0.153 $X2=0.135 $Y2=0.137
cc_52 N_CLK_c_62_p N_8_c_198_n 8.28523e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_53 N_CLK_c_59_p N_8_c_199_n 3.19268e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_54 N_CLK_c_62_p N_8_c_199_n 0.00100806f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_55 N_CLK_c_59_p N_8_c_201_n 9.01736e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_56 N_CLK_c_62_p N_8_c_202_n 3.57731e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_57 N_CLK_c_59_p N_8_c_203_n 6.50246e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_58 N_CLK_c_62_p N_8_c_203_n 4.93535e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_59 N_CLK_M4_g N_9_M6_g 2.13359e-19 $X=0.351 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_60 N_CLK_c_59_p N_9_c_231_n 2.15534e-19 $X=0.582 $Y=0.153 $X2=0.135 $Y2=0.135
cc_61 N_CLK_M7_g N_9_M8_g 0.00268443f $X=0.621 $Y=0.0675 $X2=0.135 $Y2=0.125
cc_62 N_CLK_M9_g N_9_M8_g 0.00328721f $X=0.729 $Y=0.0675 $X2=0.135 $Y2=0.125
cc_63 N_CLK_M10_g N_9_M8_g 2.48122e-19 $X=0.783 $Y=0.0675 $X2=0.135 $Y2=0.125
cc_64 N_CLK_c_84_p N_9_M8_g 3.92861e-19 $X=0.684 $Y=0.187 $X2=0.135 $Y2=0.125
cc_65 N_CLK_c_85_p N_9_c_236_n 0.0010353f $X=0.621 $Y=0.135 $X2=0.135 $Y2=0.137
cc_66 N_CLK_M9_g N_9_M11_g 2.48122e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_67 N_CLK_M10_g N_9_M11_g 0.00328721f $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_68 N_CLK_c_46_n N_9_c_239_n 3.0124e-19 $X=0.296 $Y=0.153 $X2=0 $Y2=0
cc_69 N_CLK_c_47_n N_9_c_239_n 5.62774e-19 $X=0.243 $Y=0.133 $X2=0 $Y2=0
cc_70 N_CLK_c_46_n N_9_c_229_n 3.44788e-19 $X=0.296 $Y=0.153 $X2=0 $Y2=0
cc_71 N_CLK_c_56_p N_9_c_242_n 4.44284e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_72 N_CLK_c_56_p N_9_c_243_n 2.54113e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_73 N_CLK_M4_g N_9_c_244_n 2.69763e-19 $X=0.351 $Y=0.0405 $X2=0 $Y2=0
cc_74 N_CLK_c_51_p N_9_c_245_n 5.33107e-19 $X=0.3555 $Y=0.1335 $X2=0 $Y2=0
cc_75 N_CLK_c_56_p N_9_c_245_n 4.41663e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_76 N_CLK_c_59_p N_9_c_245_n 3.17785e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_77 N_CLK_c_69_p N_9_c_245_n 0.00207315f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_78 N_CLK_c_62_p N_9_c_245_n 0.00252282f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_79 N_CLK_M4_g N_9_c_250_n 2.92102e-19 $X=0.351 $Y=0.0405 $X2=0 $Y2=0
cc_80 N_CLK_c_59_p N_9_c_251_n 6.2848e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_81 N_CLK_M7_g N_9_c_252_n 3.73075e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_82 N_CLK_c_66_p N_9_c_252_n 4.18576e-19 $X=0.621 $Y=0.133 $X2=0 $Y2=0
cc_83 N_CLK_c_59_p N_9_c_254_n 2.73788e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_84 N_CLK_c_69_p N_9_c_254_n 3.82241e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_85 N_CLK_c_59_p N_9_c_256_n 3.8223e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_86 N_CLK_c_62_p N_9_c_256_n 0.00487387f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_87 N_CLK_M9_g N_9_c_258_n 5.5355e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_88 N_CLK_c_108_p N_9_c_258_n 7.26266e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_89 N_CLK_c_109_p N_9_c_258_n 8.01493e-19 $X=0.688 $Y=0.187 $X2=0 $Y2=0
cc_90 N_CLK_c_110_p N_9_c_261_n 8.01493e-19 $X=0.6935 $Y=0.187 $X2=0 $Y2=0
cc_91 N_CLK_c_111_p N_9_c_262_n 0.00118098f $X=0.756 $Y=0.162 $X2=0 $Y2=0
cc_92 N_CLK_M10_g N_9_c_263_n 3.81593e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_93 N_CLK_c_108_p N_9_c_263_n 8.51921e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_94 N_CLK_c_84_p N_9_c_265_n 9.869e-19 $X=0.684 $Y=0.187 $X2=0 $Y2=0
cc_95 N_CLK_c_66_p N_9_c_265_n 0.00110905f $X=0.621 $Y=0.133 $X2=0 $Y2=0
cc_96 N_CLK_M10_g N_10_M12_g 2.13359e-19 $X=0.783 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_97 N_CLK_c_108_p N_10_c_334_n 7.52823e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_98 N_CLK_c_118_p N_10_c_335_n 0.049634f $X=0.747 $Y=0.187 $X2=0 $Y2=0
cc_99 N_CLK_c_110_p N_10_c_335_n 0.0086729f $X=0.6935 $Y=0.187 $X2=0 $Y2=0
cc_100 N_CLK_M9_g N_10_c_337_n 2.89162e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_101 N_CLK_c_110_p N_10_c_337_n 0.00454542f $X=0.6935 $Y=0.187 $X2=0 $Y2=0
cc_102 N_CLK_M10_g N_10_c_339_n 2.82957e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_103 N_CLK_c_108_p N_10_c_339_n 3.8451e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_104 N_CLK_M10_g N_10_c_341_n 3.96202e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_105 N_CLK_c_43_n N_12_c_392_n 0.00569573f $X=0.243 $Y=0.1335 $X2=0.135
+ $Y2=0.125
cc_106 N_CLK_c_46_n N_12_c_392_n 3.78132e-19 $X=0.296 $Y=0.153 $X2=0.135
+ $Y2=0.125
cc_107 N_CLK_c_47_n N_12_c_392_n 3.48512e-19 $X=0.243 $Y=0.133 $X2=0.135
+ $Y2=0.125
cc_108 N_CLK_c_47_n N_13_c_401_n 5.62774e-19 $X=0.243 $Y=0.133 $X2=0.135
+ $Y2=0.135
cc_109 N_CLK_M4_g N_14_c_406_n 0.00280362f $X=0.351 $Y=0.0405 $X2=0.135
+ $Y2=0.125
cc_110 N_CLK_c_51_p N_14_c_406_n 2.06383e-19 $X=0.3555 $Y=0.1335 $X2=0.135
+ $Y2=0.125
cc_111 N_CLK_c_69_p N_14_c_406_n 9.52591e-19 $X=0.405 $Y=0.134 $X2=0.135
+ $Y2=0.125
cc_112 N_CLK_c_69_p N_15_c_416_n 8.7631e-19 $X=0.405 $Y=0.134 $X2=0.135
+ $Y2=0.135
cc_113 N_7_M3_g N_8_M5_g 2.82885e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_114 N_7_c_141_n N_8_c_197_n 0.00121003f $X=0.596 $Y=0.0675 $X2=0 $Y2=0
cc_115 N_7_c_142_n N_8_c_207_n 4.7624e-19 $X=0.596 $Y=0.2025 $X2=0.056 $Y2=0.216
cc_116 N_7_c_150_n N_8_c_207_n 2.60284e-19 $X=0.568 $Y=0.189 $X2=0.056 $Y2=0.216
cc_117 N_7_c_161_p N_8_c_209_n 0.00134983f $X=0.577 $Y=0.086 $X2=0.18 $Y2=0.233
cc_118 N_7_c_162_p N_8_c_210_n 0.00134983f $X=0.577 $Y=0.232 $X2=0 $Y2=0
cc_119 N_7_c_163_p N_8_c_211_n 0.00134983f $X=0.568 $Y=0.116 $X2=0.126 $Y2=0.036
cc_120 N_7_c_154_n N_8_c_203_n 0.00134983f $X=0.568 $Y=0.1525 $X2=0.189
+ $Y2=0.045
cc_121 N_7_c_152_n N_8_c_213_n 0.00134983f $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.224
cc_122 N_7_c_150_n N_8_c_214_n 6.67324e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.135
cc_123 N_7_c_156_n N_8_c_215_n 0.00134983f $X=0.568 $Y=0.222 $X2=0.189 $Y2=0.135
cc_124 N_7_c_150_n N_8_c_216_n 5.91796e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.063
cc_125 N_7_c_142_n N_9_c_231_n 2.39572e-19 $X=0.596 $Y=0.2025 $X2=0.189
+ $Y2=0.135
cc_126 N_7_c_134_n N_9_c_239_n 0.00130909f $X=0.297 $Y=0.133 $X2=0.189 $Y2=0.045
cc_127 N_7_c_150_n N_9_c_269_n 5.00653e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.135
cc_128 N_7_M3_g N_9_c_270_n 2.70372e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.198
cc_129 N_7_c_149_n N_9_c_270_n 4.88088e-19 $X=0.31 $Y=0.189 $X2=0.189 $Y2=0.198
cc_130 N_7_c_150_n N_9_c_270_n 3.79017e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.198
cc_131 N_7_c_136_n N_9_c_270_n 0.00265354f $X=0.306 $Y=0.189 $X2=0.189 $Y2=0.198
cc_132 N_7_c_134_n N_9_c_243_n 0.0011395f $X=0.297 $Y=0.133 $X2=0.189 $Y2=0.2235
cc_133 N_7_c_134_n N_9_c_275_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_134 N_7_c_134_n N_9_c_276_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_135 N_7_c_134_n N_9_c_244_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_136 N_7_c_134_n N_9_c_245_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_137 N_7_M7_s N_9_c_279_n 3.12749e-19 $X=0.611 $Y=0.0675 $X2=0 $Y2=0
cc_138 N_7_c_141_n N_9_c_279_n 0.00290811f $X=0.596 $Y=0.0675 $X2=0 $Y2=0
cc_139 N_7_c_161_p N_9_c_279_n 0.0027674f $X=0.577 $Y=0.086 $X2=0 $Y2=0
cc_140 N_7_c_150_n N_9_c_282_n 2.35423e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_141 N_7_c_150_n N_9_c_254_n 3.37429e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_142 N_7_c_150_n N_9_c_256_n 6.95518e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_143 N_7_c_147_n N_9_c_285_n 3.43042e-19 $X=0.594 $Y=0.086 $X2=0 $Y2=0
cc_144 N_7_c_163_p N_9_c_286_n 2.63767e-19 $X=0.568 $Y=0.116 $X2=0 $Y2=0
cc_145 N_7_c_149_n N_9_c_287_n 0.00126174f $X=0.31 $Y=0.189 $X2=0 $Y2=0
cc_146 N_7_c_150_n N_9_c_287_n 4.35645e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_147 N_7_c_191_p N_10_c_337_n 2.63066e-19 $X=0.594 $Y=0.232 $X2=0.189
+ $Y2=0.135
cc_148 N_7_c_134_n N_12_c_392_n 0.00330923f $X=0.297 $Y=0.133 $X2=0.125
+ $Y2=0.054
cc_149 N_7_c_150_n N_14_c_406_n 3.19426e-19 $X=0.568 $Y=0.189 $X2=0.125
+ $Y2=0.054
cc_150 N_8_M5_g N_9_M6_g 0.00268443f $X=0.405 $Y=0.0405 $X2=0.243 $Y2=0.1335
cc_151 N_8_c_201_n N_9_M6_g 5.07993e-19 $X=0.473 $Y=0.082 $X2=0.243 $Y2=0.1335
cc_152 N_8_c_219_p N_9_c_243_n 5.2508e-19 $X=0.405 $Y=0.082 $X2=0.756 $Y2=0.162
cc_153 N_8_c_198_n N_9_c_276_n 0.00112828f $X=0.406 $Y=0.082 $X2=0.243 $Y2=0.153
cc_154 N_8_c_211_n N_9_c_244_n 2.05549e-19 $X=0.5125 $Y=0.12 $X2=0.243 $Y2=0.153
cc_155 N_8_c_213_n N_9_c_245_n 2.05549e-19 $X=0.5125 $Y=0.181 $X2=0 $Y2=0
cc_156 N_8_M5_g N_9_c_295_n 2.1403e-19 $X=0.405 $Y=0.0405 $X2=0.621 $Y2=0.153
cc_157 N_8_c_197_n N_9_c_295_n 0.00315628f $X=0.484 $Y=0.0405 $X2=0.621
+ $Y2=0.153
cc_158 N_8_c_198_n N_9_c_295_n 0.00735896f $X=0.406 $Y=0.082 $X2=0.621 $Y2=0.153
cc_159 N_8_c_214_n N_9_c_282_n 9.42345e-19 $X=0.5125 $Y=0.199 $X2=0.243
+ $Y2=0.133
cc_160 N_8_c_216_n N_9_c_282_n 2.89066e-19 $X=0.486 $Y=0.233 $X2=0.243 $Y2=0.133
cc_161 N_8_M5_g N_9_c_256_n 5.18398e-19 $X=0.405 $Y=0.0405 $X2=0.621 $Y2=0.133
cc_162 N_9_M11_g N_10_M12_g 0.00268443f $X=0.837 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_163 N_9_M11_g N_10_M13_g 2.13359e-19 $X=0.837 $Y=0.0675 $X2=0.091 $Y2=0.054
cc_164 N_9_c_303_p N_10_c_345_n 9.85984e-19 $X=0.837 $Y=0.135 $X2=0.108
+ $Y2=0.054
cc_165 N_9_c_304_p N_10_c_334_n 6.30417e-19 $X=0.666 $Y=0.036 $X2=0.054
+ $Y2=0.233
cc_166 N_9_c_305_p N_10_c_334_n 2.62833e-19 $X=0.675 $Y=0.095 $X2=0.054
+ $Y2=0.233
cc_167 N_9_c_261_n N_10_c_334_n 5.00181e-19 $X=0.747 $Y=0.108 $X2=0.054
+ $Y2=0.233
cc_168 N_9_c_262_n N_10_c_334_n 0.00105563f $X=0.765 $Y=0.108 $X2=0.054
+ $Y2=0.233
cc_169 N_9_c_263_n N_10_c_334_n 5.00181e-19 $X=0.7965 $Y=0.108 $X2=0.054
+ $Y2=0.233
cc_170 N_9_c_258_n N_10_c_339_n 4.7867e-19 $X=0.742 $Y=0.108 $X2=0.189 $Y2=0.135
cc_171 N_9_M11_g N_10_c_341_n 3.37536e-19 $X=0.837 $Y=0.0675 $X2=0.189 $Y2=0.127
cc_172 N_9_c_311_p N_10_c_341_n 5.50762e-19 $X=0.675 $Y=0.073 $X2=0.189
+ $Y2=0.127
cc_173 N_9_c_261_n N_10_c_341_n 0.00883267f $X=0.747 $Y=0.108 $X2=0.189
+ $Y2=0.127
cc_174 N_9_c_313_p N_10_c_355_n 0.00104987f $X=0.837 $Y=0.133 $X2=0 $Y2=0
cc_175 N_9_c_314_p N_10_c_356_n 0.00104987f $X=0.837 $Y=0.108 $X2=0 $Y2=0
cc_176 N_9_c_313_p N_10_c_357_n 8.04994e-19 $X=0.837 $Y=0.133 $X2=0 $Y2=0
cc_177 N_9_c_262_n N_10_c_358_n 4.7867e-19 $X=0.765 $Y=0.108 $X2=0 $Y2=0
cc_178 N_9_c_239_n N_12_c_392_n 0.00144308f $X=0.27 $Y=0.2025 $X2=0.125
+ $Y2=0.054
cc_179 N_9_c_242_n N_12_c_392_n 5.41912e-19 $X=0.349 $Y=0.036 $X2=0.125
+ $Y2=0.054
cc_180 N_9_c_243_n N_12_c_392_n 0.00307808f $X=0.324 $Y=0.036 $X2=0.125
+ $Y2=0.054
cc_181 N_9_c_239_n N_13_c_401_n 0.00390769f $X=0.27 $Y=0.2025 $X2=0.189
+ $Y2=0.135
cc_182 N_9_c_229_n N_13_c_401_n 3.931e-19 $X=0.27 $Y=0.232 $X2=0.189 $Y2=0.135
cc_183 N_9_c_239_n N_14_c_406_n 0.00165821f $X=0.27 $Y=0.2025 $X2=0.125
+ $Y2=0.054
cc_184 N_9_c_269_n N_14_c_406_n 0.00263901f $X=0.349 $Y=0.232 $X2=0.125
+ $Y2=0.054
cc_185 N_9_c_270_n N_14_c_406_n 0.00105007f $X=0.324 $Y=0.232 $X2=0.125
+ $Y2=0.054
cc_186 N_9_c_243_n N_14_c_406_n 5.71406e-19 $X=0.324 $Y=0.036 $X2=0.125
+ $Y2=0.054
cc_187 N_9_c_326_p N_14_c_406_n 0.0127725f $X=0.358 $Y=0.223 $X2=0.125 $Y2=0.054
cc_188 N_9_c_254_n N_14_c_406_n 2.57332e-19 $X=0.392 $Y=0.19 $X2=0.125 $Y2=0.054
cc_189 N_9_c_243_n N_15_c_416_n 0.00179714f $X=0.324 $Y=0.036 $X2=0.189
+ $Y2=0.135
cc_190 N_9_c_329_p N_15_c_416_n 0.00159984f $X=0.392 $Y=0.036 $X2=0.189
+ $Y2=0.135
cc_191 N_9_c_330_p N_15_c_416_n 4.19603e-19 $X=0.358 $Y=0.036 $X2=0.189
+ $Y2=0.135
cc_192 N_9_c_258_n N_16_M9_d 5.62141e-19 $X=0.742 $Y=0.108 $X2=0.189 $Y2=0.0675
cc_193 N_9_c_332_p N_17_M11_s 4.38445e-19 $X=0.828 $Y=0.108 $X2=0.189 $Y2=0.0675
cc_194 N_10_c_345_n N_GCLK_M13_d 3.7444e-19 $X=0.945 $Y=0.136 $X2=0.243
+ $Y2=0.1335
cc_195 N_10_c_345_n N_GCLK_M27_d 3.87022e-19 $X=0.945 $Y=0.136 $X2=0 $Y2=0
cc_196 N_10_c_345_n N_GCLK_c_378_n 8.43851e-19 $X=0.945 $Y=0.136 $X2=0.351
+ $Y2=0.1335
cc_197 N_10_c_362_p N_GCLK_c_378_n 0.00157438f $X=0.891 $Y=0.1675 $X2=0.351
+ $Y2=0.1335
cc_198 N_10_M13_g N_GCLK_c_380_n 4.61823e-19 $X=0.945 $Y=0.0675 $X2=0.351
+ $Y2=0.1335
cc_199 N_10_M12_g N_GCLK_c_381_n 2.25273e-19 $X=0.891 $Y=0.0675 $X2=0.621
+ $Y2=0.0675
cc_200 N_10_c_345_n N_GCLK_c_381_n 5.85939e-19 $X=0.945 $Y=0.136 $X2=0.621
+ $Y2=0.0675
cc_201 N_10_c_366_p N_GCLK_c_381_n 0.0022316f $X=0.882 $Y=0.072 $X2=0.621
+ $Y2=0.0675
cc_202 N_10_c_345_n N_GCLK_c_384_n 7.60428e-19 $X=0.945 $Y=0.136 $X2=0.621
+ $Y2=0.0675
cc_203 N_10_c_366_p N_GCLK_c_384_n 0.00160813f $X=0.882 $Y=0.072 $X2=0.621
+ $Y2=0.0675
cc_204 N_10_M13_g N_GCLK_c_386_n 4.56718e-19 $X=0.945 $Y=0.0675 $X2=0.621
+ $Y2=0.2025
cc_205 N_10_c_345_n N_GCLK_c_387_n 5.97402e-19 $X=0.945 $Y=0.136 $X2=0 $Y2=0
cc_206 N_10_c_358_n N_GCLK_c_387_n 3.48358e-19 $X=0.837 $Y=0.228 $X2=0 $Y2=0
cc_207 N_10_c_345_n GCLK 4.01182e-19 $X=0.945 $Y=0.136 $X2=0 $Y2=0
cc_208 N_10_c_355_n GCLK 7.87781e-19 $X=0.891 $Y=0.136 $X2=0 $Y2=0
cc_209 N_10_c_366_p N_GCLK_c_391_n 7.87781e-19 $X=0.882 $Y=0.072 $X2=0.783
+ $Y2=0.0675
cc_210 N_10_c_341_n N_17_M11_s 4.99504e-19 $X=0.846 $Y=0.072 $X2=0.243
+ $Y2=0.1335
cc_211 N_12_c_392_n N_13_c_401_n 9.62374e-19 $X=0.272 $Y=0.0675 $X2=0.189
+ $Y2=0.135

* END of "./ICGx2_ASAP7_75t_SRAM.pex.sp.ICGX2_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: ICGx3_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:32:22 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "ICGx3_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./ICGx3_ASAP7_75t_SRAM.pex.sp.pex"
* File: ICGx3_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:32:22 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_ICGX3_ASAP7_75T_SRAM%ENA 2 5 7 12 14 VSS
c8 14 VSS 0.00198326f $X=0.081 $Y=0.137
c9 12 VSS 0.00715247f $X=0.082 $Y=0.125
c10 5 VSS 0.00267764f $X=0.081 $Y=0.135
c11 2 VSS 0.0610973f $X=0.081 $Y=0.054
r12 12 14 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.125 $X2=0.081 $Y2=0.137
r13 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.137 $X2=0.081
+ $Y2=0.137
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%SE 2 5 7 10 VSS
c11 10 VSS 0.0013575f $X=0.135 $Y=0.125
c12 5 VSS 0.00158698f $X=0.135 $Y=0.135
c13 2 VSS 0.056849f $X=0.135 $Y=0.054
r14 10 13 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.125 $X2=0.135 $Y2=0.137
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.137 $X2=0.135
+ $Y2=0.137
r16 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%5 2 5 7 9 10 13 14 17 19 24 26 28 36 40 44 45 46 47
+ 49 VSS
c23 51 VSS 3.08662e-19 $X=0.189 $Y=0.206
c24 49 VSS 9.26001e-20 $X=0.189 $Y=0.198
c25 47 VSS 2.30045e-20 $X=0.189 $Y=0.127
c26 46 VSS 6.5293e-19 $X=0.189 $Y=0.119
c27 45 VSS 4.30607e-19 $X=0.189 $Y=0.09
c28 44 VSS 2.54814e-19 $X=0.189 $Y=0.076
c29 43 VSS 5.02744e-19 $X=0.189 $Y=0.072
c30 40 VSS 8.26035e-19 $X=0.189 $Y=0.135
c31 36 VSS 0.00146362f $X=0.144 $Y=0.036
c32 35 VSS 0.00266146f $X=0.126 $Y=0.036
c33 30 VSS 0.00201059f $X=0.108 $Y=0.036
c34 28 VSS 0.00804964f $X=0.18 $Y=0.036
c35 27 VSS 0.00324205f $X=0.162 $Y=0.233
c36 26 VSS 0.00135162f $X=0.144 $Y=0.233
c37 25 VSS 0.00344819f $X=0.126 $Y=0.233
c38 24 VSS 0.00525503f $X=0.09 $Y=0.233
c39 19 VSS 0.00468477f $X=0.18 $Y=0.233
c40 17 VSS 0.00199178f $X=0.056 $Y=0.216
c41 14 VSS 4.96055e-19 $X=0.071 $Y=0.216
c42 13 VSS 0.0085383f $X=0.108 $Y=0.054
c43 9 VSS 5.3314e-19 $X=0.125 $Y=0.054
c44 5 VSS 0.00138247f $X=0.189 $Y=0.135
c45 2 VSS 0.0577976f $X=0.189 $Y=0.0675
r46 52 53 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.223 $X2=0.189 $Y2=0.2235
r47 51 52 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.206 $X2=0.189 $Y2=0.223
r48 50 51 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.199 $X2=0.189 $Y2=0.206
r49 49 50 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.198 $X2=0.189 $Y2=0.199
r50 48 49 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.184 $X2=0.189 $Y2=0.198
r51 46 47 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.119 $X2=0.189 $Y2=0.127
r52 45 46 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.09 $X2=0.189 $Y2=0.119
r53 44 45 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.076 $X2=0.189 $Y2=0.09
r54 43 44 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.072 $X2=0.189 $Y2=0.076
r55 42 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.063 $X2=0.189 $Y2=0.072
r56 40 48 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.184
r57 40 47 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.127
r58 38 53 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.224 $X2=0.189 $Y2=0.2235
r59 37 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r60 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r61 30 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r62 28 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r63 28 36 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.144 $Y2=0.036
r64 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.233 $X2=0.162 $Y2=0.233
r65 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.233 $X2=0.144 $Y2=0.233
r66 24 25 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.233 $X2=0.126 $Y2=0.233
r67 21 24 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.233 $X2=0.09 $Y2=0.233
r68 19 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.233 $X2=0.189 $Y2=0.224
r69 19 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.233 $X2=0.162 $Y2=0.233
r70 17 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.233 $X2=0.054
+ $Y2=0.233
r71 14 17 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r72 13 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r73 10 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.054 $X2=0.108 $Y2=0.054
r74 9 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.054 $X2=0.108 $Y2=0.054
r75 5 40 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r76 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r77 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%CLK 2 5 8 14 17 19 22 27 30 33 35 40 42 45 47 48 49
+ 52 65 66 69 70 71 75 80 91 92 VSS
c89 102 VSS 1.751e-20 $X=0.621 $Y=0.15
c90 92 VSS 6.23569e-19 $X=0.405 $Y=0.134
c91 91 VSS 0.00812781f $X=0.405 $Y=0.134
c92 80 VSS 2.48826e-19 $X=0.621 $Y=0.133
c93 75 VSS 9.46764e-19 $X=0.243 $Y=0.133
c94 71 VSS 6.07691e-19 $X=0.6015 $Y=0.153
c95 70 VSS 0.004187f $X=0.582 $Y=0.153
c96 69 VSS 0.00101808f $X=0.621 $Y=0.153
c97 68 VSS 0.00158411f $X=0.621 $Y=0.153
c98 66 VSS 0.00142963f $X=0.3595 $Y=0.153
c99 65 VSS 0.00275092f $X=0.296 $Y=0.153
c100 52 VSS 0.00127138f $X=0.756 $Y=0.162
c101 49 VSS 1.14519e-19 $X=0.6935 $Y=0.187
c102 48 VSS 1.68783e-19 $X=0.688 $Y=0.187
c103 47 VSS 4.53034e-19 $X=0.684 $Y=0.187
c104 46 VSS 0.00437089f $X=0.666 $Y=0.187
c105 43 VSS 9.76836e-19 $X=0.63 $Y=0.187
c106 42 VSS 0.00282432f $X=0.747 $Y=0.187
c107 40 VSS 6.59173e-19 $X=0.3555 $Y=0.1335
c108 33 VSS 0.00745385f $X=0.783 $Y=0.162
c109 30 VSS 0.0599108f $X=0.783 $Y=0.0675
c110 22 VSS 0.0599326f $X=0.729 $Y=0.0675
c111 17 VSS 0.00243599f $X=0.621 $Y=0.135
c112 14 VSS 0.0620989f $X=0.621 $Y=0.0675
c113 8 VSS 0.0605267f $X=0.351 $Y=0.0405
c114 2 VSS 0.0605352f $X=0.243 $Y=0.1335
r115 101 102 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.147 $X2=0.621 $Y2=0.15
r116 91 92 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.405 $Y=0.134
+ $X2=0.405 $Y2=0.134
r117 80 101 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.133 $X2=0.621 $Y2=0.147
r118 70 71 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.582
+ $Y=0.153 $X2=0.6015 $Y2=0.153
r119 69 102 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.621 $Y2=0.15
r120 68 71 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M2 $thickness=3.6e-08 $X=0.621
+ $Y=0.153 $X2=0.6015 $Y2=0.153
r121 68 69 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.621 $Y=0.153 $X2=0.621
+ $Y2=0.153
r122 65 66 4.31173 $w=1.8e-08 $l=6.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.296
+ $Y=0.153 $X2=0.3595 $Y2=0.153
r123 64 92 0.725694 $w=3.2e-08 $l=3.36861e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.4305 $Y=0.153 $X2=0.405 $Y2=0.134
r124 63 70 10.7963 $w=1.8e-08 $l=1.59e-07 $layer=M2 $thickness=3.6e-08 $X=0.423
+ $Y=0.153 $X2=0.582 $Y2=0.153
r125 63 66 4.31173 $w=1.8e-08 $l=6.35e-08 $layer=M2 $thickness=3.6e-08 $X=0.423
+ $Y=0.153 $X2=0.3595 $Y2=0.153
r126 63 64 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.423 $Y=0.153 $X2=0.423
+ $Y2=0.153
r127 60 75 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.133
r128 59 65 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.296 $Y2=0.153
r129 59 60 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.153 $X2=0.243
+ $Y2=0.153
r130 57 69 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.178 $X2=0.621 $Y2=0.153
r131 52 53 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.756 $Y=0.162 $X2=0.756
+ $Y2=0.162
r132 50 52 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.178 $X2=0.756 $Y2=0.162
r133 48 49 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.688
+ $Y=0.187 $X2=0.6935 $Y2=0.187
r134 47 48 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.187 $X2=0.688 $Y2=0.187
r135 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.187 $X2=0.684 $Y2=0.187
r136 45 49 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.699
+ $Y=0.187 $X2=0.6935 $Y2=0.187
r137 43 57 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.63 $Y=0.187 $X2=0.621 $Y2=0.178
r138 43 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.187 $X2=0.666 $Y2=0.187
r139 42 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.747 $Y=0.187 $X2=0.756 $Y2=0.178
r140 42 45 3.25926 $w=1.8e-08 $l=4.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.187 $X2=0.699 $Y2=0.187
r141 40 91 41.0143 $w=2.5e-08 $l=4.95e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.3555 $Y=0.1335 $X2=0.405 $Y2=0.1335
r142 33 53 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.783
+ $Y=0.162 $X2=0.756 $Y2=0.162
r143 33 35 202.311 $w=2e-08 $l=5.4e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.162 $X2=0.783 $Y2=0.216
r144 30 33 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.162
r145 25 53 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.162 $X2=0.756 $Y2=0.162
r146 25 27 202.311 $w=2e-08 $l=5.4e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.162 $X2=0.729 $Y2=0.216
r147 22 25 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.162
r148 17 80 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.133 $X2=0.621
+ $Y2=0.133
r149 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2025
r150 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r151 11 40 4.28571 $w=2.1e-08 $l=4.5e-09 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.1335 $X2=0.3555 $Y2=0.1335
r152 8 11 348.425 $w=2e-08 $l=9.3e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0405 $X2=0.351 $Y2=0.1335
r153 2 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.133 $X2=0.243
+ $Y2=0.133
r154 2 5 258.509 $w=2e-08 $l=6.9e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1335 $X2=0.243 $Y2=0.2025
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%7 2 5 7 9 12 14 17 22 32 34 35 41 43 48 51 52 64 65
+ 67 71 VSS
c61 72 VSS 2.26979e-19 $X=0.308 $Y=0.189
c62 71 VSS 4.78866e-20 $X=0.306 $Y=0.189
c63 67 VSS 4.14661e-19 $X=0.568 $Y=0.222
c64 65 VSS 8.24918e-19 $X=0.568 $Y=0.1525
c65 64 VSS 3.2551e-19 $X=0.568 $Y=0.116
c66 52 VSS 7.99983e-19 $X=0.568 $Y=0.189
c67 51 VSS 0.00784196f $X=0.568 $Y=0.189
c68 48 VSS 6.70853e-19 $X=0.31 $Y=0.189
c69 44 VSS 8.31083e-19 $X=0.5855 $Y=0.232
c70 43 VSS 0.00225204f $X=0.577 $Y=0.232
c71 41 VSS 0.00296213f $X=0.594 $Y=0.232
c72 35 VSS 1.50276e-19 $X=0.5855 $Y=0.086
c73 34 VSS 2.75727e-19 $X=0.577 $Y=0.086
c74 32 VSS 6.35967e-19 $X=0.594 $Y=0.086
c75 22 VSS 0.00287748f $X=0.297 $Y=0.133
c76 17 VSS 0.00554583f $X=0.596 $Y=0.2025
c77 14 VSS 4.06194e-19 $X=0.611 $Y=0.2025
c78 12 VSS 0.00700617f $X=0.596 $Y=0.0675
c79 9 VSS 3.3425e-19 $X=0.611 $Y=0.0675
c80 5 VSS 0.00109246f $X=0.297 $Y=0.1335
c81 2 VSS 0.0591582f $X=0.297 $Y=0.0675
r82 71 72 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.189 $X2=0.308 $Y2=0.189
r83 68 71 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.306 $Y2=0.189
r84 66 67 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.196 $X2=0.568 $Y2=0.222
r85 64 65 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.116 $X2=0.568 $Y2=0.1525
r86 52 66 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.189 $X2=0.568 $Y2=0.196
r87 52 65 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.189 $X2=0.568 $Y2=0.1525
r88 51 52 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.568 $Y=0.189 $X2=0.568
+ $Y2=0.189
r89 48 72 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.31
+ $Y=0.189 $X2=0.308 $Y2=0.189
r90 47 51 17.5185 $w=1.8e-08 $l=2.58e-07 $layer=M2 $thickness=3.6e-08 $X=0.31
+ $Y=0.189 $X2=0.568 $Y2=0.189
r91 47 48 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.31 $Y=0.189 $X2=0.31
+ $Y2=0.189
r92 43 44 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.577
+ $Y=0.232 $X2=0.5855 $Y2=0.232
r93 41 44 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.232 $X2=0.5855 $Y2=0.232
r94 38 67 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.223 $X2=0.568 $Y2=0.222
r95 37 43 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.232 $X2=0.577 $Y2=0.232
r96 37 38 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.232 $X2=0.568 $Y2=0.223
r97 34 35 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.577
+ $Y=0.086 $X2=0.5855 $Y2=0.086
r98 32 35 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.086 $X2=0.5855 $Y2=0.086
r99 29 64 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.095 $X2=0.568 $Y2=0.116
r100 28 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.086 $X2=0.577 $Y2=0.086
r101 28 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.568
+ $Y=0.086 $X2=0.568 $Y2=0.095
r102 20 68 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.18 $X2=0.297 $Y2=0.189
r103 20 22 3.19136 $w=1.8e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.18 $X2=0.297 $Y2=0.133
r104 17 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.232
+ $X2=0.594 $Y2=0.232
r105 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2025 $X2=0.596 $Y2=0.2025
r106 12 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.086
+ $X2=0.594 $Y2=0.086
r107 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0675 $X2=0.596 $Y2=0.0675
r108 5 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.133 $X2=0.297
+ $Y2=0.133
r109 5 7 359.664 $w=2e-08 $l=9.6e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.1335 $X2=0.297 $Y2=0.2295
r110 2 5 247.269 $w=2e-08 $l=6.6e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.1335
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%8 2 5 7 9 12 14 17 19 21 30 31 34 35 36 37 38 39 40
+ 42 VSS
c34 48 VSS 0.00202496f $X=0.503 $Y=0.233
c35 47 VSS 0.00196174f $X=0.5125 $Y=0.233
c36 42 VSS 0.00220406f $X=0.486 $Y=0.233
c37 40 VSS 4.74628e-19 $X=0.5125 $Y=0.2115
c38 39 VSS 4.02544e-19 $X=0.5125 $Y=0.199
c39 38 VSS 0.00128405f $X=0.5125 $Y=0.181
c40 37 VSS 3.27036e-19 $X=0.5125 $Y=0.162
c41 36 VSS 7.69748e-19 $X=0.5125 $Y=0.144
c42 35 VSS 8.43604e-19 $X=0.5125 $Y=0.12
c43 34 VSS 7.4117e-19 $X=0.5125 $Y=0.224
c44 32 VSS 2.34012e-20 $X=0.4795 $Y=0.082
c45 31 VSS 3.09176e-19 $X=0.473 $Y=0.082
c46 30 VSS 5.46116e-19 $X=0.447 $Y=0.082
c47 29 VSS 1.3164e-20 $X=0.414 $Y=0.082
c48 21 VSS 3.42062e-19 $X=0.406 $Y=0.082
c49 19 VSS 6.62699e-19 $X=0.503 $Y=0.082
c50 17 VSS 0.00305014f $X=0.484 $Y=0.2295
c51 12 VSS 0.00680979f $X=0.484 $Y=0.0405
c52 5 VSS 0.00260336f $X=0.405 $Y=0.082
c53 2 VSS 0.0587788f $X=0.405 $Y=0.0405
r54 48 49 0.322531 $w=1.8e-08 $l=4.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.503
+ $Y=0.233 $X2=0.50775 $Y2=0.233
r55 47 49 0.322531 $w=1.8e-08 $l=4.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.233 $X2=0.50775 $Y2=0.233
r56 42 48 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.233 $X2=0.503 $Y2=0.233
r57 39 40 0.793941 $w=1.9e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.199 $X2=0.5125 $Y2=0.2115
r58 38 39 1.14327 $w=1.9e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.181 $X2=0.5125 $Y2=0.199
r59 37 38 1.20679 $w=1.9e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.162 $X2=0.5125 $Y2=0.181
r60 36 37 1.14327 $w=1.9e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.144 $X2=0.5125 $Y2=0.162
r61 35 36 1.52437 $w=1.9e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.12 $X2=0.5125 $Y2=0.144
r62 34 47 0.0384781 $w=1.9e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.224 $X2=0.5125 $Y2=0.233
r63 34 40 0.793941 $w=1.9e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.224 $X2=0.5125 $Y2=0.2115
r64 33 35 1.84194 $w=1.9e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5125
+ $Y=0.091 $X2=0.5125 $Y2=0.12
r65 31 32 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.473
+ $Y=0.082 $X2=0.4795 $Y2=0.082
r66 30 31 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.082 $X2=0.473 $Y2=0.082
r67 29 30 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.082 $X2=0.447 $Y2=0.082
r68 27 32 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.082 $X2=0.4795 $Y2=0.082
r69 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.082 $X2=0.486
+ $Y2=0.082
r70 21 29 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.406
+ $Y=0.082 $X2=0.414 $Y2=0.082
r71 19 33 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.503 $Y=0.082 $X2=0.5125 $Y2=0.091
r72 19 27 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.503
+ $Y=0.082 $X2=0.486 $Y2=0.082
r73 17 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.233 $X2=0.486
+ $Y2=0.233
r74 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2295 $X2=0.484 $Y2=0.2295
r75 12 28 35.8185 $w=2.4e-08 $l=4.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0405 $X2=0.486 $Y2=0.082
r76 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0405 $X2=0.484 $Y2=0.0405
r77 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.406 $Y=0.082 $X2=0.406
+ $Y2=0.082
r78 5 7 552.609 $w=2e-08 $l=1.475e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.082 $X2=0.405 $Y2=0.2295
r79 2 5 155.48 $w=2e-08 $l=4.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0405 $X2=0.405 $Y2=0.082
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%9 2 5 7 10 13 15 18 21 23 25 30 33 37 38 41 43 49
+ 50 53 58 59 60 61 62 64 65 67 68 69 70 72 75 77 79 86 88 89 90 91 93 94 95 96
+ 97 98 101 107 110 VSS
c102 113 VSS 8.63727e-20 $X=0.837 $Y=0.125
c103 110 VSS 3.88312e-19 $X=0.837 $Y=0.133
c104 107 VSS 3.25689e-19 $X=0.837 $Y=0.108
c105 101 VSS 6.07255e-19 $X=0.675 $Y=0.133
c106 99 VSS 4.28973e-19 $X=0.675 $Y=0.108
c107 98 VSS 1.77849e-19 $X=0.358 $Y=0.19
c108 97 VSS 0.00171031f $X=0.358 $Y=0.036
c109 96 VSS 3.03415e-19 $X=0.7965 $Y=0.108
c110 95 VSS 2.5364e-19 $X=0.765 $Y=0.108
c111 94 VSS 7.79718e-20 $X=0.747 $Y=0.108
c112 93 VSS 0.00151883f $X=0.742 $Y=0.108
c113 91 VSS 6.2055e-19 $X=0.828 $Y=0.108
c114 90 VSS 8.07734e-20 $X=0.675 $Y=0.097
c115 89 VSS 4.90266e-19 $X=0.675 $Y=0.095
c116 88 VSS 1.49364e-19 $X=0.675 $Y=0.081
c117 87 VSS 1.86503e-19 $X=0.675 $Y=0.077
c118 86 VSS 5.68609e-19 $X=0.675 $Y=0.073
c119 85 VSS 8.45284e-19 $X=0.675 $Y=0.063
c120 84 VSS 6.05801e-20 $X=0.675 $Y=0.099
c121 80 VSS 5.01043e-19 $X=0.453 $Y=0.19
c122 79 VSS 0.00167287f $X=0.447 $Y=0.19
c123 78 VSS 3.25412e-19 $X=0.396 $Y=0.19
c124 77 VSS 0.00110887f $X=0.392 $Y=0.19
c125 75 VSS 8.00008e-19 $X=0.459 $Y=0.19
c126 72 VSS 0.00146505f $X=0.63 $Y=0.036
c127 71 VSS 2.9457e-19 $X=0.612 $Y=0.036
c128 70 VSS 0.00428093f $X=0.609 $Y=0.036
c129 69 VSS 0.00316044f $X=0.559 $Y=0.036
c130 68 VSS 0.0128446f $X=0.522 $Y=0.036
c131 67 VSS 0.00218374f $X=0.392 $Y=0.036
c132 65 VSS 0.00760784f $X=0.666 $Y=0.036
c133 64 VSS 7.19963e-19 $X=0.358 $Y=0.223
c134 62 VSS 3.15222e-19 $X=0.358 $Y=0.18
c135 61 VSS 5.76653e-19 $X=0.358 $Y=0.162
c136 60 VSS 7.37599e-19 $X=0.358 $Y=0.12
c137 59 VSS 2.16018e-19 $X=0.358 $Y=0.091
c138 57 VSS 5.27349e-19 $X=0.358 $Y=0.072
c139 53 VSS 0.00330518f $X=0.324 $Y=0.036
c140 50 VSS 0.0043866f $X=0.349 $Y=0.036
c141 49 VSS 0.00260946f $X=0.324 $Y=0.232
c142 48 VSS 0.00204527f $X=0.288 $Y=0.232
c143 43 VSS 0.00102923f $X=0.27 $Y=0.232
c144 41 VSS 0.00444971f $X=0.349 $Y=0.232
c145 40 VSS 6.58864e-19 $X=0.27 $Y=0.2295
c146 37 VSS 0.00138123f $X=0.27 $Y=0.2025
c147 32 VSS 5.70081e-19 $X=0.324 $Y=0.0405
c148 21 VSS 0.00193767f $X=0.837 $Y=0.135
c149 18 VSS 0.0569005f $X=0.837 $Y=0.0675
c150 13 VSS 0.00220177f $X=0.675 $Y=0.135
c151 10 VSS 0.0575264f $X=0.675 $Y=0.0675
c152 5 VSS 0.00218509f $X=0.459 $Y=0.19
c153 2 VSS 0.062866f $X=0.459 $Y=0.0405
r154 112 113 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.117 $X2=0.837 $Y2=0.125
r155 110 113 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.133 $X2=0.837 $Y2=0.125
r156 107 112 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.108 $X2=0.837 $Y2=0.117
r157 103 104 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.116 $X2=0.675 $Y2=0.117
r158 101 104 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.133 $X2=0.675 $Y2=0.117
r159 99 103 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.108 $X2=0.675 $Y2=0.116
r160 95 96 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.765
+ $Y=0.108 $X2=0.7965 $Y2=0.108
r161 94 95 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.747
+ $Y=0.108 $X2=0.765 $Y2=0.108
r162 93 94 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.742
+ $Y=0.108 $X2=0.747 $Y2=0.108
r163 92 99 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.108 $X2=0.675 $Y2=0.108
r164 92 93 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.108 $X2=0.742 $Y2=0.108
r165 91 107 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.108 $X2=0.837 $Y2=0.108
r166 91 96 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.108 $X2=0.7965 $Y2=0.108
r167 89 90 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.095 $X2=0.675 $Y2=0.097
r168 88 89 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.081 $X2=0.675 $Y2=0.095
r169 87 88 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.077 $X2=0.675 $Y2=0.081
r170 86 87 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.073 $X2=0.675 $Y2=0.077
r171 85 86 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.063 $X2=0.675 $Y2=0.073
r172 84 99 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.099 $X2=0.675 $Y2=0.108
r173 84 90 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.099 $X2=0.675 $Y2=0.097
r174 83 85 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.045 $X2=0.675 $Y2=0.063
r175 79 80 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.447
+ $Y=0.19 $X2=0.453 $Y2=0.19
r176 78 79 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.19 $X2=0.447 $Y2=0.19
r177 77 78 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.392
+ $Y=0.19 $X2=0.396 $Y2=0.19
r178 75 80 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.19 $X2=0.453 $Y2=0.19
r179 73 98 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.19 $X2=0.358 $Y2=0.19
r180 73 77 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.19 $X2=0.392 $Y2=0.19
r181 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.63 $Y2=0.036
r182 70 71 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.609
+ $Y=0.036 $X2=0.612 $Y2=0.036
r183 69 70 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.559
+ $Y=0.036 $X2=0.609 $Y2=0.036
r184 68 69 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.559 $Y2=0.036
r185 67 68 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.392
+ $Y=0.036 $X2=0.522 $Y2=0.036
r186 66 97 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.036 $X2=0.358 $Y2=0.036
r187 66 67 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.036 $X2=0.392 $Y2=0.036
r188 65 83 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.036 $X2=0.675 $Y2=0.045
r189 65 72 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.63 $Y2=0.036
r190 63 98 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.199 $X2=0.358 $Y2=0.19
r191 63 64 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.199 $X2=0.358 $Y2=0.223
r192 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.162 $X2=0.358 $Y2=0.18
r193 60 61 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.12 $X2=0.358 $Y2=0.162
r194 59 60 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.091 $X2=0.358 $Y2=0.12
r195 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.073 $X2=0.358 $Y2=0.091
r196 57 58 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.072 $X2=0.358 $Y2=0.073
r197 56 98 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.181 $X2=0.358 $Y2=0.19
r198 56 62 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.181 $X2=0.358 $Y2=0.18
r199 55 97 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.045 $X2=0.358 $Y2=0.036
r200 55 57 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.358
+ $Y=0.045 $X2=0.358 $Y2=0.072
r201 52 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r202 50 97 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.349
+ $Y=0.036 $X2=0.358 $Y2=0.036
r203 50 52 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.349
+ $Y=0.036 $X2=0.324 $Y2=0.036
r204 48 49 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.232 $X2=0.324 $Y2=0.232
r205 43 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.232 $X2=0.288 $Y2=0.232
r206 41 64 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.349 $Y=0.232 $X2=0.358 $Y2=0.223
r207 41 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.349
+ $Y=0.232 $X2=0.324 $Y2=0.232
r208 38 40 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2295 $X2=0.27 $Y2=0.2295
r209 37 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.232 $X2=0.27
+ $Y2=0.232
r210 34 40 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2655 $Y=0.216 $X2=0.27 $Y2=0.2295
r211 34 37 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.2655 $Y=0.216 $X2=0.2655 $Y2=0.189
r212 33 37 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.189 $X2=0.2655 $Y2=0.189
r213 30 32 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0405 $X2=0.324 $Y2=0.0405
r214 29 53 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r215 26 32 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.054 $X2=0.324 $Y2=0.0405
r216 26 29 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.3195 $Y=0.054 $X2=0.3195 $Y2=0.081
r217 25 29 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.081 $X2=0.3195 $Y2=0.081
r218 21 110 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.133
+ $X2=0.837 $Y2=0.133
r219 21 23 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.837
+ $Y=0.135 $X2=0.837 $Y2=0.216
r220 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0675 $X2=0.837 $Y2=0.135
r221 13 101 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.133
+ $X2=0.675 $Y2=0.133
r222 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.216
r223 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0675 $X2=0.675 $Y2=0.135
r224 5 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.19 $X2=0.459
+ $Y2=0.19
r225 5 7 147.987 $w=2e-08 $l=3.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.19 $X2=0.459 $Y2=0.2295
r226 2 5 560.102 $w=2e-08 $l=1.495e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0405 $X2=0.459 $Y2=0.19
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%10 2 7 10 15 18 21 23 25 26 29 30 31 34 35 36 48 49
+ 50 55 62 65 67 68 76 VSS
c45 76 VSS 0.00355073f $X=0.837 $Y=0.228
c46 75 VSS 1.56305e-19 $X=0.837 $Y=0.225
c47 74 VSS 7.66292e-19 $X=0.837 $Y=0.222
c48 72 VSS 0.00240875f $X=0.837 $Y=0.231
c49 68 VSS 4.0488e-19 $X=0.837 $Y=0.197
c50 67 VSS 6.32944e-19 $X=0.891 $Y=0.1675
c51 65 VSS 3.96463e-19 $X=0.891 $Y=0.1175
c52 62 VSS 2.31452e-19 $X=0.891 $Y=0.136
c53 60 VSS 2.2993e-19 $X=0.891 $Y=0.188
c54 57 VSS 0.00387746f $X=0.882 $Y=0.197
c55 56 VSS 0.00379396f $X=0.879 $Y=0.072
c56 55 VSS 0.00352836f $X=0.846 $Y=0.072
c57 50 VSS 6.46876e-20 $X=0.882 $Y=0.072
c58 49 VSS 0.00229769f $X=0.7875 $Y=0.231
c59 48 VSS 0.00805297f $X=0.765 $Y=0.231
c60 39 VSS 0.00656914f $X=0.81 $Y=0.216
c61 35 VSS 6.59309e-19 $X=0.827 $Y=0.216
c62 34 VSS 0.00617068f $X=0.702 $Y=0.216
c63 30 VSS 7.72153e-19 $X=0.719 $Y=0.216
c64 29 VSS 0.00468946f $X=0.756 $Y=0.0675
c65 25 VSS 7.90436e-19 $X=0.773 $Y=0.0675
c66 21 VSS 0.0120908f $X=0.999 $Y=0.136
c67 18 VSS 0.0647964f $X=0.999 $Y=0.0675
c68 10 VSS 0.0615177f $X=0.945 $Y=0.0675
c69 2 VSS 0.057881f $X=0.891 $Y=0.0675
r70 75 76 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.228
r71 74 75 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.222 $X2=0.837 $Y2=0.225
r72 73 74 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.206 $X2=0.837 $Y2=0.222
r73 72 76 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.231 $X2=0.837 $Y2=0.228
r74 68 73 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.197 $X2=0.837 $Y2=0.206
r75 66 67 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.147 $X2=0.891 $Y2=0.1675
r76 64 65 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.099 $X2=0.891 $Y2=0.1175
r77 62 66 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.136 $X2=0.891 $Y2=0.147
r78 62 65 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.136 $X2=0.891 $Y2=0.1175
r79 60 67 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.188 $X2=0.891 $Y2=0.1675
r80 59 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.081 $X2=0.891 $Y2=0.099
r81 58 68 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.197 $X2=0.837 $Y2=0.197
r82 57 60 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.197 $X2=0.891 $Y2=0.188
r83 57 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.197 $X2=0.846 $Y2=0.197
r84 55 56 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.846
+ $Y=0.072 $X2=0.879 $Y2=0.072
r85 52 55 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.072 $X2=0.846 $Y2=0.072
r86 50 59 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.072 $X2=0.891 $Y2=0.081
r87 50 56 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.072 $X2=0.879 $Y2=0.072
r88 48 49 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.765
+ $Y=0.231 $X2=0.7875 $Y2=0.231
r89 46 49 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.231 $X2=0.7875 $Y2=0.231
r90 42 48 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.231 $X2=0.765 $Y2=0.231
r91 40 72 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.231 $X2=0.837 $Y2=0.231
r92 40 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.231 $X2=0.81 $Y2=0.231
r93 39 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.231 $X2=0.81
+ $Y2=0.231
r94 36 39 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.216 $X2=0.81 $Y2=0.216
r95 35 39 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.216 $X2=0.81 $Y2=0.216
r96 34 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.231 $X2=0.702
+ $Y2=0.231
r97 31 34 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.216 $X2=0.702 $Y2=0.216
r98 30 34 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.216 $X2=0.702 $Y2=0.216
r99 29 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.072 $X2=0.756
+ $Y2=0.072
r100 26 29 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.756 $Y2=0.0675
r101 25 29 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.756 $Y2=0.0675
r102 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.136 $X2=0.999 $Y2=0.2025
r103 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.136
r104 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.945
+ $Y=0.136 $X2=0.999 $Y2=0.136
r105 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.136 $X2=0.945 $Y2=0.2025
r106 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.0675 $X2=0.945 $Y2=0.136
r107 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.891
+ $Y=0.136 $X2=0.945 $Y2=0.136
r108 5 62 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.891 $Y=0.136 $X2=0.891
+ $Y2=0.136
r109 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.136 $X2=0.891 $Y2=0.2025
r110 2 5 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.0675 $X2=0.891 $Y2=0.136
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%GCLK 1 2 6 11 12 15 16 21 23 24 31 33 44 46 VSS
c18 48 VSS 4.30151e-19 $X=1.053 $Y=0.2155
c19 46 VSS 0.00228126f $X=1.053 $Y=0.1145
c20 45 VSS 8.85605e-19 $X=1.053 $Y=0.063
c21 44 VSS 0.00433352f $X=1.057 $Y=0.166
c22 42 VSS 4.55454e-19 $X=1.053 $Y=0.225
c23 33 VSS 0.00191952f $X=0.918 $Y=0.234
c24 31 VSS 0.0181449f $X=1.044 $Y=0.234
c25 30 VSS 0.00692279f $X=1.026 $Y=0.036
c26 24 VSS 0.0104348f $X=0.918 $Y=0.036
c27 23 VSS 0.0039905f $X=0.918 $Y=0.036
c28 21 VSS 0.0181177f $X=1.044 $Y=0.036
c29 19 VSS 0.00719225f $X=1.024 $Y=0.2025
c30 15 VSS 0.010473f $X=0.918 $Y=0.2025
c31 11 VSS 5.38922e-19 $X=0.935 $Y=0.2025
c32 9 VSS 2.69461e-19 $X=1.024 $Y=0.0675
c33 1 VSS 5.38922e-19 $X=0.935 $Y=0.0675
r34 47 48 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.206 $X2=1.053 $Y2=0.2155
r35 45 46 3.49691 $w=1.8e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.063 $X2=1.053 $Y2=0.1145
r36 44 47 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.166 $X2=1.053 $Y2=0.206
r37 44 46 3.49691 $w=1.8e-08 $l=5.15e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.166 $X2=1.053 $Y2=0.1145
r38 42 48 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.225 $X2=1.053 $Y2=0.2155
r39 41 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.045 $X2=1.053 $Y2=0.063
r40 33 39 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.234 $X2=1.026 $Y2=0.234
r41 31 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.234 $X2=1.053 $Y2=0.225
r42 31 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.234 $X2=1.026 $Y2=0.234
r43 29 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.036 $X2=1.026
+ $Y2=0.036
r44 23 29 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.036 $X2=1.026 $Y2=0.036
r45 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.036 $X2=0.918
+ $Y2=0.036
r46 21 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.036 $X2=1.053 $Y2=0.045
r47 21 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=1.026 $Y2=0.036
r48 19 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.234 $X2=1.026
+ $Y2=0.234
r49 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.2025 $X2=1.024 $Y2=0.2025
r50 15 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.234 $X2=0.918
+ $Y2=0.234
r51 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.2025 $X2=0.918 $Y2=0.2025
r52 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.935 $Y=0.2025 $X2=0.918 $Y2=0.2025
r53 9 30 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=1.026
+ $Y=0.0675 $X2=1.026 $Y2=0.036
r54 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=1.009
+ $Y=0.0675 $X2=1.024 $Y2=0.0675
r55 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.918
+ $Y=0.0675 $X2=0.918 $Y2=0.036
r56 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.901
+ $Y=0.0675 $X2=0.918 $Y2=0.0675
r57 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.935
+ $Y=0.0675 $X2=0.918 $Y2=0.0675
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%12 1 6 9 VSS
c9 9 VSS 0.0197042f $X=0.272 $Y=0.0675
c10 6 VSS 3.61939e-19 $X=0.287 $Y=0.0675
c11 4 VSS 3.25039e-19 $X=0.214 $Y=0.0675
r12 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.272 $Y2=0.0675
r13 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.214
+ $Y=0.0675 $X2=0.272 $Y2=0.0675
r14 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.214 $Y2=0.0675
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%13 1 2 5 VSS
c5 5 VSS 0.00678699f $X=0.216 $Y=0.2025
c6 1 VSS 6.50078e-19 $X=0.233 $Y=0.2025
r7 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.2025 $X2=0.216 $Y2=0.2025
r8 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.216 $Y2=0.2025
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%14 1 6 9 VSS
c10 9 VSS 0.018833f $X=0.38 $Y=0.2295
c11 6 VSS 3.72954e-19 $X=0.395 $Y=0.2295
c12 4 VSS 3.77944e-19 $X=0.322 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.2295 $X2=0.38 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.2295 $X2=0.38 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2295 $X2=0.322 $Y2=0.2295
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%15 1 2 5 VSS
c4 5 VSS 0.00485144f $X=0.378 $Y=0.0405
c5 1 VSS 6.8236e-19 $X=0.395 $Y=0.0405
r6 2 5 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.0405 $X2=0.378 $Y2=0.0405
r7 1 5 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0405 $X2=0.378 $Y2=0.0405
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%16 1 2 VSS
c1 1 VSS 0.00221026f $X=0.719 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0675 $X2=0.685 $Y2=0.0675
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%17 1 2 VSS
c2 1 VSS 0.00230546f $X=0.827 $Y=0.0675
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.827
+ $Y=0.0675 $X2=0.793 $Y2=0.0675
.ends

.subckt PM_ICGX3_ASAP7_75T_SRAM%18 1 2 VSS
c0 1 VSS 0.00242486f $X=0.125 $Y=0.216
r1 1 2 25.1852 $w=5.4e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.216 $X2=0.091 $Y2=0.216
.ends


* END of "./ICGx3_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt ICGx3_ASAP7_75t_SRAM  VSS VDD ENA SE CLK GCLK
* 
* GCLK	GCLK
* CLK	CLK
* SE	SE
* ENA	ENA
M0 N_5_M0_d N_ENA_M0_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 VSS N_SE_M1_g N_5_M1_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 N_12_M2_d N_5_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_9_M3_d N_7_M3_g N_12_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M4 N_15_M4_d N_CLK_M4_g N_9_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.341
+ $Y=0.027
M5 VSS N_8_M5_g N_15_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.395
+ $Y=0.027
M6 N_8_M6_d N_9_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449 $Y=0.027
M7 VSS N_CLK_M7_g N_7_M7_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M8 VSS N_9_M8_g N_16_M8_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M9 N_16_M9_d N_CLK_M9_g N_10_M9_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M10 N_17_M10_d N_CLK_M10_g N_10_M10_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.773 $Y=0.027
M11 VSS N_9_M11_g N_17_M11_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.027
M12 N_GCLK_M12_d N_10_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.027
M13 N_GCLK_M13_d N_10_M13_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.027
M14 N_GCLK_M14_d N_10_M14_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M15 N_18_M15_d N_ENA_M15_g N_5_M15_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2
+ $X=0.071 $Y=0.189
M16 VDD N_SE_M16_g N_18_M16_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M17 N_13_M17_d N_5_M17_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M18 N_9_M18_d N_CLK_M18_g N_13_M18_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M19 N_14_M19_d N_7_M19_g N_9_M19_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.287 $Y=0.216
M20 VDD N_8_M20_g N_14_M20_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.395
+ $Y=0.216
M21 N_8_M21_d N_9_M21_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.216
M22 VDD N_CLK_M22_g N_7_M22_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M23 N_10_M23_d N_9_M23_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.665
+ $Y=0.189
M24 VDD N_CLK_M24_g N_10_M24_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.719
+ $Y=0.189
M25 VDD N_CLK_M25_g N_10_M25_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.773
+ $Y=0.189
M26 N_10_M26_d N_9_M26_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.827
+ $Y=0.189
M27 N_GCLK_M27_d N_10_M27_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.162
M28 N_GCLK_M28_d N_10_M28_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.162
M29 N_GCLK_M29_d N_10_M29_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
*
* 
* .include "ICGx3_ASAP7_75t_SRAM.pex.sp.ICGX3_ASAP7_75T_SRAM.pxi"
* BEGIN of "./ICGx3_ASAP7_75t_SRAM.pex.sp.ICGX3_ASAP7_75T_SRAM.pxi"
* File: ICGx3_ASAP7_75t_SRAM.pex.sp.ICGX3_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:32:22 2017
* 
x_PM_ICGX3_ASAP7_75T_SRAM%ENA N_ENA_M0_g N_ENA_c_2_p N_ENA_M15_g ENA N_ENA_c_6_p
+ VSS PM_ICGX3_ASAP7_75T_SRAM%ENA
x_PM_ICGX3_ASAP7_75T_SRAM%SE N_SE_M1_g N_SE_c_10_n N_SE_M16_g SE VSS
+ PM_ICGX3_ASAP7_75T_SRAM%SE
x_PM_ICGX3_ASAP7_75T_SRAM%5 N_5_M2_g N_5_c_26_n N_5_M17_g N_5_M1_s N_5_M0_d
+ N_5_c_21_n N_5_M15_s N_5_c_22_n N_5_c_40_p N_5_c_23_n N_5_c_27_n N_5_c_41_p
+ N_5_c_29_n N_5_c_34_p N_5_c_37_p N_5_c_31_n N_5_c_38_p N_5_c_35_p N_5_c_39_p
+ VSS PM_ICGX3_ASAP7_75T_SRAM%5
x_PM_ICGX3_ASAP7_75T_SRAM%CLK N_CLK_c_43_n N_CLK_M18_g N_CLK_M4_g N_CLK_M7_g
+ N_CLK_c_84_p N_CLK_M22_g N_CLK_M9_g N_CLK_M24_g N_CLK_M10_g N_CLK_c_107_p
+ N_CLK_M25_g N_CLK_c_51_p N_CLK_c_117_p CLK N_CLK_c_83_p N_CLK_c_108_p
+ N_CLK_c_109_p N_CLK_c_110_p N_CLK_c_46_n N_CLK_c_56_p N_CLK_c_53_p
+ N_CLK_c_59_p N_CLK_c_52_p N_CLK_c_47_n N_CLK_c_66_p N_CLK_c_69_p N_CLK_c_62_p
+ VSS PM_ICGX3_ASAP7_75T_SRAM%CLK
x_PM_ICGX3_ASAP7_75T_SRAM%7 N_7_M3_g N_7_c_138_n N_7_M19_g N_7_M7_s N_7_c_140_n
+ N_7_M22_s N_7_c_141_n N_7_c_133_n N_7_c_146_n N_7_c_160_p N_7_c_147_n
+ N_7_c_190_p N_7_c_161_p N_7_c_148_n N_7_c_149_n N_7_c_151_n N_7_c_162_p
+ N_7_c_153_n N_7_c_155_n N_7_c_135_n VSS PM_ICGX3_ASAP7_75T_SRAM%7
x_PM_ICGX3_ASAP7_75T_SRAM%8 N_8_M5_g N_8_c_218_p N_8_M20_g N_8_M6_d N_8_c_196_n
+ N_8_M21_d N_8_c_206_n N_8_c_208_n N_8_c_197_n N_8_c_198_n N_8_c_200_n
+ N_8_c_209_n N_8_c_210_n N_8_c_201_n N_8_c_202_n N_8_c_212_n N_8_c_213_n
+ N_8_c_214_n N_8_c_215_n VSS PM_ICGX3_ASAP7_75T_SRAM%8
x_PM_ICGX3_ASAP7_75T_SRAM%9 N_9_M6_g N_9_c_264_n N_9_M21_g N_9_M8_g N_9_c_233_n
+ N_9_M23_g N_9_M11_g N_9_c_299_p N_9_M26_g N_9_M3_d N_9_M4_s N_9_M18_d
+ N_9_c_236_n N_9_M19_s N_9_c_266_n N_9_c_227_n N_9_c_267_n N_9_c_239_n
+ N_9_c_240_n N_9_c_272_n N_9_c_273_n N_9_c_241_n N_9_c_242_n N_9_c_247_n
+ N_9_c_322_p N_9_c_300_p N_9_c_325_p N_9_c_291_n N_9_c_248_n N_9_c_276_n
+ N_9_c_249_n N_9_c_279_n N_9_c_251_n N_9_c_253_n N_9_c_307_p N_9_c_282_n
+ N_9_c_301_p N_9_c_283_n N_9_c_328_p N_9_c_255_n N_9_c_258_n N_9_c_259_n
+ N_9_c_260_n N_9_c_326_p N_9_c_284_n N_9_c_262_n N_9_c_310_p N_9_c_309_p VSS
+ PM_ICGX3_ASAP7_75T_SRAM%9
x_PM_ICGX3_ASAP7_75T_SRAM%10 N_10_M12_g N_10_M27_g N_10_M13_g N_10_M28_g N_10_M14_g
+ N_10_c_341_n N_10_M29_g N_10_M10_s N_10_M9_s N_10_c_330_n N_10_M24_s
+ N_10_M23_d N_10_c_331_n N_10_M26_d N_10_M25_s N_10_c_333_n N_10_c_335_n
+ N_10_c_363_p N_10_c_337_n N_10_c_351_n N_10_c_352_n N_10_c_358_p N_10_c_353_n
+ N_10_c_354_n VSS PM_ICGX3_ASAP7_75T_SRAM%10
x_PM_ICGX3_ASAP7_75T_SRAM%GCLK N_GCLK_M13_d N_GCLK_M12_d N_GCLK_M14_d N_GCLK_M28_d
+ N_GCLK_M27_d N_GCLK_c_376_n N_GCLK_M29_d N_GCLK_c_378_n N_GCLK_c_380_n
+ N_GCLK_c_383_n N_GCLK_c_385_n N_GCLK_c_387_n GCLK N_GCLK_c_391_n VSS
+ PM_ICGX3_ASAP7_75T_SRAM%GCLK
x_PM_ICGX3_ASAP7_75T_SRAM%12 N_12_M2_d N_12_M3_s N_12_c_392_n VSS
+ PM_ICGX3_ASAP7_75T_SRAM%12
x_PM_ICGX3_ASAP7_75T_SRAM%13 N_13_M18_s N_13_M17_d N_13_c_401_n VSS
+ PM_ICGX3_ASAP7_75T_SRAM%13
x_PM_ICGX3_ASAP7_75T_SRAM%14 N_14_M19_d N_14_M20_s N_14_c_406_n VSS
+ PM_ICGX3_ASAP7_75T_SRAM%14
x_PM_ICGX3_ASAP7_75T_SRAM%15 N_15_M5_s N_15_M4_d N_15_c_416_n VSS
+ PM_ICGX3_ASAP7_75T_SRAM%15
x_PM_ICGX3_ASAP7_75T_SRAM%16 N_16_M9_d N_16_M8_s VSS PM_ICGX3_ASAP7_75T_SRAM%16
x_PM_ICGX3_ASAP7_75T_SRAM%17 N_17_M11_s N_17_M10_d VSS PM_ICGX3_ASAP7_75T_SRAM%17
x_PM_ICGX3_ASAP7_75T_SRAM%18 N_18_M16_s N_18_M15_d VSS PM_ICGX3_ASAP7_75T_SRAM%18
cc_1 N_ENA_M0_g N_SE_M1_g 0.00328721f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_ENA_c_2_p N_SE_c_10_n 9.35826e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 ENA SE 0.00588002f $X=0.082 $Y=0.125 $X2=0.135 $Y2=0.125
cc_4 N_ENA_M0_g N_5_M2_g 2.13359e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 ENA N_5_c_21_n 6.06976e-19 $X=0.082 $Y=0.125 $X2=0.135 $Y2=0.137
cc_6 N_ENA_c_6_p N_5_c_22_n 0.00174918f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_7 N_ENA_M0_g N_5_c_23_n 2.28086e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_8 N_ENA_c_6_p N_5_c_23_n 0.00499899f $X=0.081 $Y=0.137 $X2=0 $Y2=0
cc_9 N_SE_M1_g N_5_M2_g 0.00268443f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_10 N_SE_c_10_n N_5_c_26_n 9.11034e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_11 N_SE_M1_g N_5_c_27_n 2.59938e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_12 SE N_5_c_27_n 0.00123553f $X=0.135 $Y=0.125 $X2=0 $Y2=0
cc_13 N_SE_M1_g N_5_c_29_n 2.84283e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_14 SE N_5_c_29_n 0.001038f $X=0.135 $Y=0.125 $X2=0 $Y2=0
cc_15 SE N_5_c_31_n 0.00457266f $X=0.135 $Y=0.125 $X2=0 $Y2=0
cc_16 N_SE_M1_g N_CLK_c_43_n 2.13359e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_17 N_5_M2_g N_CLK_c_43_n 0.00341068f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_18 N_5_c_26_n N_CLK_c_43_n 8.10277e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.054
cc_19 N_5_c_34_p N_CLK_c_46_n 3.51913e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_20 N_5_c_35_p N_CLK_c_47_n 0.00253589f $X=0.189 $Y=0.127 $X2=0 $Y2=0
cc_21 N_5_M2_g N_7_M3_g 2.82885e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_22 N_5_c_37_p N_7_c_133_n 3.23824e-19 $X=0.189 $Y=0.076 $X2=0 $Y2=0
cc_23 N_5_c_38_p N_7_c_133_n 2.18117e-19 $X=0.189 $Y=0.119 $X2=0 $Y2=0
cc_24 N_5_c_39_p N_7_c_135_n 2.18117e-19 $X=0.189 $Y=0.198 $X2=0 $Y2=0
cc_25 N_5_c_40_p N_9_c_227_n 4.49022e-19 $X=0.18 $Y=0.233 $X2=0 $Y2=0
cc_26 N_5_c_41_p N_12_c_392_n 0.00246673f $X=0.18 $Y=0.036 $X2=0 $Y2=0
cc_27 N_5_c_34_p N_13_c_401_n 0.00182314f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_28 N_CLK_c_43_n N_7_M3_g 0.00355599f $X=0.243 $Y=0.1335 $X2=0.135 $Y2=0.054
cc_29 N_CLK_M4_g N_7_M3_g 0.00355599f $X=0.351 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_30 N_CLK_c_43_n N_7_c_138_n 8.50652e-19 $X=0.243 $Y=0.1335 $X2=0.135
+ $Y2=0.135
cc_31 N_CLK_c_51_p N_7_c_138_n 9.50591e-19 $X=0.3555 $Y=0.1335 $X2=0.135
+ $Y2=0.135
cc_32 N_CLK_c_52_p N_7_c_140_n 2.51466e-19 $X=0.6015 $Y=0.153 $X2=0.135
+ $Y2=0.137
cc_33 N_CLK_c_53_p N_7_c_141_n 6.1856e-19 $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_34 N_CLK_c_52_p N_7_c_141_n 2.98103e-19 $X=0.6015 $Y=0.153 $X2=0 $Y2=0
cc_35 N_CLK_c_46_n N_7_c_133_n 0.0010183f $X=0.296 $Y=0.153 $X2=0 $Y2=0
cc_36 N_CLK_c_56_p N_7_c_133_n 5.3655e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_37 N_CLK_c_47_n N_7_c_133_n 0.00252905f $X=0.243 $Y=0.133 $X2=0 $Y2=0
cc_38 N_CLK_c_52_p N_7_c_146_n 2.62247e-19 $X=0.6015 $Y=0.153 $X2=0 $Y2=0
cc_39 N_CLK_c_59_p N_7_c_147_n 2.62247e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_40 N_CLK_c_56_p N_7_c_148_n 2.46239e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_41 N_CLK_c_56_p N_7_c_149_n 0.0242262f $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_42 N_CLK_c_62_p N_7_c_149_n 4.84045e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_43 N_CLK_c_53_p N_7_c_151_n 0.0017697f $X=0.621 $Y=0.153 $X2=0 $Y2=0
cc_44 N_CLK_c_59_p N_7_c_151_n 4.75571e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_45 N_CLK_c_59_p N_7_c_153_n 3.96692e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_46 N_CLK_c_66_p N_7_c_153_n 0.00167205f $X=0.621 $Y=0.133 $X2=0 $Y2=0
cc_47 N_CLK_c_59_p N_7_c_155_n 2.46239e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_48 N_CLK_M4_g N_8_M5_g 0.00341068f $X=0.351 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_49 N_CLK_c_69_p N_8_M5_g 0.00207156f $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.054
cc_50 N_CLK_c_62_p N_8_M5_g 2.24185e-19 $X=0.405 $Y=0.134 $X2=0.135 $Y2=0.054
cc_51 N_CLK_c_59_p N_8_c_196_n 2.35254e-19 $X=0.582 $Y=0.153 $X2=0.135 $Y2=0.137
cc_52 N_CLK_c_62_p N_8_c_197_n 8.28523e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_53 N_CLK_c_59_p N_8_c_198_n 3.19268e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_54 N_CLK_c_62_p N_8_c_198_n 0.00100725f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_55 N_CLK_c_59_p N_8_c_200_n 9.01736e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_56 N_CLK_c_62_p N_8_c_201_n 3.5769e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_57 N_CLK_c_59_p N_8_c_202_n 6.41758e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_58 N_CLK_c_62_p N_8_c_202_n 4.93535e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_59 N_CLK_M4_g N_9_M6_g 2.13359e-19 $X=0.351 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_60 N_CLK_M7_g N_9_M8_g 0.00268443f $X=0.621 $Y=0.0675 $X2=0.135 $Y2=0.125
cc_61 N_CLK_M9_g N_9_M8_g 0.00328721f $X=0.729 $Y=0.0675 $X2=0.135 $Y2=0.125
cc_62 N_CLK_M10_g N_9_M8_g 2.48122e-19 $X=0.783 $Y=0.0675 $X2=0.135 $Y2=0.125
cc_63 N_CLK_c_83_p N_9_M8_g 3.92861e-19 $X=0.684 $Y=0.187 $X2=0.135 $Y2=0.125
cc_64 N_CLK_c_84_p N_9_c_233_n 9.91457e-19 $X=0.621 $Y=0.135 $X2=0.135 $Y2=0.137
cc_65 N_CLK_M9_g N_9_M11_g 2.48122e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_66 N_CLK_M10_g N_9_M11_g 0.00328721f $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_67 N_CLK_c_46_n N_9_c_236_n 3.0124e-19 $X=0.296 $Y=0.153 $X2=0 $Y2=0
cc_68 N_CLK_c_47_n N_9_c_236_n 5.62774e-19 $X=0.243 $Y=0.133 $X2=0 $Y2=0
cc_69 N_CLK_c_46_n N_9_c_227_n 3.44788e-19 $X=0.296 $Y=0.153 $X2=0 $Y2=0
cc_70 N_CLK_c_56_p N_9_c_239_n 4.44284e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_71 N_CLK_c_56_p N_9_c_240_n 2.54113e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_72 N_CLK_M4_g N_9_c_241_n 2.69763e-19 $X=0.351 $Y=0.0405 $X2=0 $Y2=0
cc_73 N_CLK_c_51_p N_9_c_242_n 5.33107e-19 $X=0.3555 $Y=0.1335 $X2=0 $Y2=0
cc_74 N_CLK_c_56_p N_9_c_242_n 4.41663e-19 $X=0.3595 $Y=0.153 $X2=0 $Y2=0
cc_75 N_CLK_c_59_p N_9_c_242_n 3.17785e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_76 N_CLK_c_69_p N_9_c_242_n 0.025735f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_77 N_CLK_c_62_p N_9_c_242_n 0.00252282f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_78 N_CLK_M4_g N_9_c_247_n 2.92102e-19 $X=0.351 $Y=0.0405 $X2=0 $Y2=0
cc_79 N_CLK_c_59_p N_9_c_248_n 6.2848e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_80 N_CLK_M7_g N_9_c_249_n 3.73075e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_81 N_CLK_c_66_p N_9_c_249_n 4.18576e-19 $X=0.621 $Y=0.133 $X2=0 $Y2=0
cc_82 N_CLK_c_59_p N_9_c_251_n 2.73788e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_83 N_CLK_c_69_p N_9_c_251_n 3.82241e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_84 N_CLK_c_59_p N_9_c_253_n 3.8223e-19 $X=0.582 $Y=0.153 $X2=0 $Y2=0
cc_85 N_CLK_c_62_p N_9_c_253_n 0.00487778f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_86 N_CLK_M9_g N_9_c_255_n 5.5355e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_87 N_CLK_c_107_p N_9_c_255_n 3.64914e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_88 N_CLK_c_108_p N_9_c_255_n 8.0008e-19 $X=0.688 $Y=0.187 $X2=0 $Y2=0
cc_89 N_CLK_c_109_p N_9_c_258_n 8.0008e-19 $X=0.6935 $Y=0.187 $X2=0 $Y2=0
cc_90 N_CLK_c_110_p N_9_c_259_n 0.00118098f $X=0.756 $Y=0.162 $X2=0 $Y2=0
cc_91 N_CLK_M10_g N_9_c_260_n 3.81593e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_92 N_CLK_c_107_p N_9_c_260_n 4.3841e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_93 N_CLK_c_83_p N_9_c_262_n 9.869e-19 $X=0.684 $Y=0.187 $X2=0 $Y2=0
cc_94 N_CLK_c_66_p N_9_c_262_n 0.00110905f $X=0.621 $Y=0.133 $X2=0 $Y2=0
cc_95 N_CLK_M10_g N_10_M12_g 2.13359e-19 $X=0.783 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_96 N_CLK_c_107_p N_10_c_330_n 3.02943e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_97 N_CLK_c_117_p N_10_c_331_n 0.049634f $X=0.747 $Y=0.187 $X2=0 $Y2=0
cc_98 N_CLK_c_109_p N_10_c_331_n 0.0086729f $X=0.6935 $Y=0.187 $X2=0 $Y2=0
cc_99 N_CLK_M9_g N_10_c_333_n 2.89162e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_100 N_CLK_c_109_p N_10_c_333_n 0.00454542f $X=0.6935 $Y=0.187 $X2=0 $Y2=0
cc_101 N_CLK_M10_g N_10_c_335_n 2.82957e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_102 N_CLK_c_107_p N_10_c_335_n 3.8451e-19 $X=0.783 $Y=0.162 $X2=0 $Y2=0
cc_103 N_CLK_M10_g N_10_c_337_n 3.96202e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_104 N_CLK_c_43_n N_12_c_392_n 0.00570295f $X=0.243 $Y=0.1335 $X2=0.135
+ $Y2=0.125
cc_105 N_CLK_c_46_n N_12_c_392_n 3.91758e-19 $X=0.296 $Y=0.153 $X2=0.135
+ $Y2=0.125
cc_106 N_CLK_c_47_n N_12_c_392_n 3.48512e-19 $X=0.243 $Y=0.133 $X2=0.135
+ $Y2=0.125
cc_107 N_CLK_c_47_n N_13_c_401_n 5.62774e-19 $X=0.243 $Y=0.133 $X2=0.135
+ $Y2=0.135
cc_108 N_CLK_M4_g N_14_c_406_n 0.00275062f $X=0.351 $Y=0.0405 $X2=0.135
+ $Y2=0.125
cc_109 N_CLK_c_51_p N_14_c_406_n 2.06383e-19 $X=0.3555 $Y=0.1335 $X2=0.135
+ $Y2=0.125
cc_110 N_CLK_c_69_p N_14_c_406_n 8.83266e-19 $X=0.405 $Y=0.134 $X2=0.135
+ $Y2=0.125
cc_111 N_CLK_c_69_p N_15_c_416_n 7.69733e-19 $X=0.405 $Y=0.134 $X2=0.135
+ $Y2=0.135
cc_112 N_7_M3_g N_8_M5_g 2.82885e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_113 N_7_c_140_n N_8_c_196_n 0.00109006f $X=0.596 $Y=0.0675 $X2=0 $Y2=0
cc_114 N_7_c_141_n N_8_c_206_n 4.54309e-19 $X=0.596 $Y=0.2025 $X2=0.056
+ $Y2=0.216
cc_115 N_7_c_149_n N_8_c_206_n 2.60284e-19 $X=0.568 $Y=0.189 $X2=0.056 $Y2=0.216
cc_116 N_7_c_160_p N_8_c_208_n 0.00134983f $X=0.577 $Y=0.086 $X2=0.18 $Y2=0.233
cc_117 N_7_c_161_p N_8_c_209_n 0.00134983f $X=0.577 $Y=0.232 $X2=0 $Y2=0
cc_118 N_7_c_162_p N_8_c_210_n 0.00134983f $X=0.568 $Y=0.116 $X2=0.126 $Y2=0.036
cc_119 N_7_c_153_n N_8_c_202_n 0.00134983f $X=0.568 $Y=0.1525 $X2=0.189
+ $Y2=0.045
cc_120 N_7_c_151_n N_8_c_212_n 0.00134983f $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.224
cc_121 N_7_c_149_n N_8_c_213_n 6.67324e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.135
cc_122 N_7_c_155_n N_8_c_214_n 0.00134983f $X=0.568 $Y=0.222 $X2=0.189 $Y2=0.135
cc_123 N_7_c_149_n N_8_c_215_n 5.91796e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.063
cc_124 N_7_c_141_n N_9_c_264_n 2.47747e-19 $X=0.596 $Y=0.2025 $X2=0.189
+ $Y2=0.135
cc_125 N_7_c_133_n N_9_c_236_n 0.00130909f $X=0.297 $Y=0.133 $X2=0.189 $Y2=0.045
cc_126 N_7_c_149_n N_9_c_266_n 5.00653e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.135
cc_127 N_7_M3_g N_9_c_267_n 2.70372e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.198
cc_128 N_7_c_148_n N_9_c_267_n 4.88088e-19 $X=0.31 $Y=0.189 $X2=0.189 $Y2=0.198
cc_129 N_7_c_149_n N_9_c_267_n 3.79017e-19 $X=0.568 $Y=0.189 $X2=0.189 $Y2=0.198
cc_130 N_7_c_135_n N_9_c_267_n 0.00265354f $X=0.306 $Y=0.189 $X2=0.189 $Y2=0.198
cc_131 N_7_c_133_n N_9_c_240_n 0.0011408f $X=0.297 $Y=0.133 $X2=0.189 $Y2=0.2235
cc_132 N_7_c_133_n N_9_c_272_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_133 N_7_c_133_n N_9_c_273_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_134 N_7_c_133_n N_9_c_241_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_135 N_7_c_133_n N_9_c_242_n 8.47314e-19 $X=0.297 $Y=0.133 $X2=0 $Y2=0
cc_136 N_7_M7_s N_9_c_276_n 3.12749e-19 $X=0.611 $Y=0.0675 $X2=0 $Y2=0
cc_137 N_7_c_140_n N_9_c_276_n 0.00290811f $X=0.596 $Y=0.0675 $X2=0 $Y2=0
cc_138 N_7_c_160_p N_9_c_276_n 0.0027674f $X=0.577 $Y=0.086 $X2=0 $Y2=0
cc_139 N_7_c_149_n N_9_c_279_n 2.35423e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_140 N_7_c_149_n N_9_c_251_n 3.37429e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_141 N_7_c_149_n N_9_c_253_n 6.95518e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_142 N_7_c_146_n N_9_c_282_n 3.43042e-19 $X=0.594 $Y=0.086 $X2=0 $Y2=0
cc_143 N_7_c_162_p N_9_c_283_n 2.65458e-19 $X=0.568 $Y=0.116 $X2=0 $Y2=0
cc_144 N_7_c_148_n N_9_c_284_n 0.00126174f $X=0.31 $Y=0.189 $X2=0 $Y2=0
cc_145 N_7_c_149_n N_9_c_284_n 4.35645e-19 $X=0.568 $Y=0.189 $X2=0 $Y2=0
cc_146 N_7_c_190_p N_10_c_333_n 2.63066e-19 $X=0.594 $Y=0.232 $X2=0.189
+ $Y2=0.184
cc_147 N_7_c_133_n N_12_c_392_n 0.00329939f $X=0.297 $Y=0.133 $X2=0.125
+ $Y2=0.054
cc_148 N_7_c_149_n N_14_c_406_n 3.19426e-19 $X=0.568 $Y=0.189 $X2=0.125
+ $Y2=0.054
cc_149 N_8_M5_g N_9_M6_g 0.00268443f $X=0.405 $Y=0.0405 $X2=0.243 $Y2=0.1335
cc_150 N_8_c_200_n N_9_M6_g 5.07993e-19 $X=0.473 $Y=0.082 $X2=0.243 $Y2=0.1335
cc_151 N_8_c_218_p N_9_c_240_n 5.2508e-19 $X=0.405 $Y=0.082 $X2=0.756 $Y2=0.162
cc_152 N_8_c_196_n N_9_c_240_n 3.84672e-19 $X=0.484 $Y=0.0405 $X2=0.756
+ $Y2=0.162
cc_153 N_8_c_197_n N_9_c_273_n 0.00112828f $X=0.406 $Y=0.082 $X2=0.243 $Y2=0.153
cc_154 N_8_M5_g N_9_c_291_n 2.1403e-19 $X=0.405 $Y=0.0405 $X2=0.621 $Y2=0.153
cc_155 N_8_c_196_n N_9_c_291_n 0.00315627f $X=0.484 $Y=0.0405 $X2=0.621
+ $Y2=0.153
cc_156 N_8_c_197_n N_9_c_291_n 0.00735876f $X=0.406 $Y=0.082 $X2=0.621 $Y2=0.153
cc_157 N_8_c_213_n N_9_c_279_n 9.42345e-19 $X=0.5125 $Y=0.199 $X2=0.243
+ $Y2=0.133
cc_158 N_8_c_215_n N_9_c_279_n 2.89066e-19 $X=0.486 $Y=0.233 $X2=0.243 $Y2=0.133
cc_159 N_8_M5_g N_9_c_253_n 5.18398e-19 $X=0.405 $Y=0.0405 $X2=0.621 $Y2=0.133
cc_160 N_9_M11_g N_10_M12_g 0.00268443f $X=0.837 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_161 N_9_M11_g N_10_M13_g 2.13359e-19 $X=0.837 $Y=0.0675 $X2=0.091 $Y2=0.054
cc_162 N_9_c_299_p N_10_c_341_n 9.44581e-19 $X=0.837 $Y=0.135 $X2=0.054
+ $Y2=0.233
cc_163 N_9_c_300_p N_10_c_330_n 6.30417e-19 $X=0.666 $Y=0.036 $X2=0.108
+ $Y2=0.036
cc_164 N_9_c_301_p N_10_c_330_n 2.62833e-19 $X=0.675 $Y=0.095 $X2=0.108
+ $Y2=0.036
cc_165 N_9_c_258_n N_10_c_330_n 5.00181e-19 $X=0.747 $Y=0.108 $X2=0.108
+ $Y2=0.036
cc_166 N_9_c_259_n N_10_c_330_n 0.00105563f $X=0.765 $Y=0.108 $X2=0.108
+ $Y2=0.036
cc_167 N_9_c_260_n N_10_c_330_n 5.00181e-19 $X=0.7965 $Y=0.108 $X2=0.108
+ $Y2=0.036
cc_168 N_9_c_255_n N_10_c_335_n 4.7805e-19 $X=0.742 $Y=0.108 $X2=0.189 $Y2=0.198
cc_169 N_9_M11_g N_10_c_337_n 3.37536e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_170 N_9_c_307_p N_10_c_337_n 5.50762e-19 $X=0.675 $Y=0.073 $X2=0 $Y2=0
cc_171 N_9_c_258_n N_10_c_337_n 0.00883267f $X=0.747 $Y=0.108 $X2=0 $Y2=0
cc_172 N_9_c_309_p N_10_c_351_n 0.00104987f $X=0.837 $Y=0.133 $X2=0 $Y2=0
cc_173 N_9_c_310_p N_10_c_352_n 0.00104987f $X=0.837 $Y=0.108 $X2=0 $Y2=0
cc_174 N_9_c_309_p N_10_c_353_n 8.04994e-19 $X=0.837 $Y=0.133 $X2=0 $Y2=0
cc_175 N_9_c_259_n N_10_c_354_n 4.7805e-19 $X=0.765 $Y=0.108 $X2=0 $Y2=0
cc_176 N_9_c_236_n N_12_c_392_n 0.00144308f $X=0.27 $Y=0.2025 $X2=0.125
+ $Y2=0.054
cc_177 N_9_c_239_n N_12_c_392_n 5.41912e-19 $X=0.349 $Y=0.036 $X2=0.125
+ $Y2=0.054
cc_178 N_9_c_240_n N_12_c_392_n 0.00295119f $X=0.324 $Y=0.036 $X2=0.125
+ $Y2=0.054
cc_179 N_9_c_236_n N_13_c_401_n 0.00390769f $X=0.27 $Y=0.2025 $X2=0.189
+ $Y2=0.135
cc_180 N_9_c_227_n N_13_c_401_n 3.96553e-19 $X=0.27 $Y=0.232 $X2=0.189 $Y2=0.135
cc_181 N_9_c_236_n N_14_c_406_n 0.00164257f $X=0.27 $Y=0.2025 $X2=0.125
+ $Y2=0.054
cc_182 N_9_c_266_n N_14_c_406_n 0.00263901f $X=0.349 $Y=0.232 $X2=0.125
+ $Y2=0.054
cc_183 N_9_c_267_n N_14_c_406_n 0.00102838f $X=0.324 $Y=0.232 $X2=0.125
+ $Y2=0.054
cc_184 N_9_c_240_n N_14_c_406_n 6.05863e-19 $X=0.324 $Y=0.036 $X2=0.125
+ $Y2=0.054
cc_185 N_9_c_322_p N_14_c_406_n 0.0127725f $X=0.358 $Y=0.223 $X2=0.125 $Y2=0.054
cc_186 N_9_c_251_n N_14_c_406_n 2.57332e-19 $X=0.392 $Y=0.19 $X2=0.125 $Y2=0.054
cc_187 N_9_c_240_n N_15_c_416_n 0.00179714f $X=0.324 $Y=0.036 $X2=0.189
+ $Y2=0.135
cc_188 N_9_c_325_p N_15_c_416_n 0.00159984f $X=0.392 $Y=0.036 $X2=0.189
+ $Y2=0.135
cc_189 N_9_c_326_p N_15_c_416_n 4.19603e-19 $X=0.358 $Y=0.036 $X2=0.189
+ $Y2=0.135
cc_190 N_9_c_255_n N_16_M9_d 5.62141e-19 $X=0.742 $Y=0.108 $X2=0.189 $Y2=0.0675
cc_191 N_9_c_328_p N_17_M11_s 4.38445e-19 $X=0.828 $Y=0.108 $X2=0.189 $Y2=0.0675
cc_192 N_10_c_341_n N_GCLK_M13_d 3.7444e-19 $X=0.999 $Y=0.136 $X2=0.243
+ $Y2=0.1335
cc_193 N_10_c_341_n N_GCLK_M28_d 3.87022e-19 $X=0.999 $Y=0.136 $X2=0.351
+ $Y2=0.1335
cc_194 N_10_c_341_n N_GCLK_c_376_n 8.43851e-19 $X=0.999 $Y=0.136 $X2=0 $Y2=0
cc_195 N_10_c_358_p N_GCLK_c_376_n 0.00158777f $X=0.891 $Y=0.1675 $X2=0 $Y2=0
cc_196 N_10_M13_g N_GCLK_c_378_n 4.61823e-19 $X=0.945 $Y=0.0675 $X2=0.729
+ $Y2=0.0675
cc_197 N_10_M14_g N_GCLK_c_378_n 4.61823e-19 $X=0.999 $Y=0.0675 $X2=0.729
+ $Y2=0.0675
cc_198 N_10_M12_g N_GCLK_c_380_n 2.25273e-19 $X=0.891 $Y=0.0675 $X2=0 $Y2=0
cc_199 N_10_c_341_n N_GCLK_c_380_n 0.00137255f $X=0.999 $Y=0.136 $X2=0 $Y2=0
cc_200 N_10_c_363_p N_GCLK_c_380_n 0.0022316f $X=0.882 $Y=0.072 $X2=0 $Y2=0
cc_201 N_10_c_341_n N_GCLK_c_383_n 7.60428e-19 $X=0.999 $Y=0.136 $X2=0.729
+ $Y2=0.162
cc_202 N_10_c_363_p N_GCLK_c_383_n 0.00163229f $X=0.882 $Y=0.072 $X2=0.729
+ $Y2=0.162
cc_203 N_10_M13_g N_GCLK_c_385_n 4.56718e-19 $X=0.945 $Y=0.0675 $X2=0 $Y2=0
cc_204 N_10_M14_g N_GCLK_c_385_n 4.56718e-19 $X=0.999 $Y=0.0675 $X2=0 $Y2=0
cc_205 N_10_c_341_n N_GCLK_c_387_n 0.00140068f $X=0.999 $Y=0.136 $X2=0.783
+ $Y2=0.162
cc_206 N_10_c_354_n N_GCLK_c_387_n 3.56146e-19 $X=0.837 $Y=0.228 $X2=0.783
+ $Y2=0.162
cc_207 N_10_c_341_n GCLK 2.12243e-19 $X=0.999 $Y=0.136 $X2=0.699 $Y2=0.187
cc_208 N_10_c_351_n GCLK 3.84006e-19 $X=0.891 $Y=0.136 $X2=0.699 $Y2=0.187
cc_209 N_10_c_363_p N_GCLK_c_391_n 3.84006e-19 $X=0.882 $Y=0.072 $X2=0.666
+ $Y2=0.187
cc_210 N_10_c_337_n N_17_M11_s 4.98974e-19 $X=0.846 $Y=0.072 $X2=0.243
+ $Y2=0.1335
cc_211 N_12_c_392_n N_13_c_401_n 9.62348e-19 $X=0.272 $Y=0.0675 $X2=0.189
+ $Y2=0.135

* END of "./ICGx3_ASAP7_75t_SRAM.pex.sp.ICGX3_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DHLx1_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:27:08 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DHLx1_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DHLx1_ASAP7_75t_SRAM.pex.sp.pex"
* File: DHLx1_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:27:08 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DHLX1_ASAP7_75T_SRAM%CLK 2 5 7 12 14 17 VSS
c18 17 VSS 5.41721e-21 $X=0.081 $Y=0.1305
c19 14 VSS 0.00699913f $X=0.081 $Y=0.135
c20 12 VSS 0.00699194f $X=0.08 $Y=0.119
c21 5 VSS 0.00183412f $X=0.081 $Y=0.135
c22 2 VSS 0.0642213f $X=0.081 $Y=0.054
r23 16 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r24 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r25 12 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.126
r26 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DHLX1_ASAP7_75T_SRAM%4 2 7 10 13 16 24 26 29 31 34 37 38 39 41 44 51 56
+ 58 59 65 66 69 76 83 84 85 87 89 90 108 109 123 VSS
c84 123 VSS 5.19505e-19 $X=0.18 $Y=0.189
c85 122 VSS 1.53285e-19 $X=0.189 $Y=0.189
c86 118 VSS 7.0154e-20 $X=0.03 $Y=0.189
c87 117 VSS 5.9624e-19 $X=0.027 $Y=0.189
c88 109 VSS 7.76097e-19 $X=0.513 $Y=0.18
c89 108 VSS 0.0574701f $X=0.513 $Y=0.18
c90 90 VSS 0.00123576f $X=0.45 $Y=0.189
c91 89 VSS 0.0038091f $X=0.414 $Y=0.189
c92 87 VSS 0.00305138f $X=0.513 $Y=0.189
c93 85 VSS 0.00251877f $X=0.29 $Y=0.189
c94 84 VSS 0.00700382f $X=0.229 $Y=0.189
c95 83 VSS 0.00149088f $X=0.351 $Y=0.189
c96 76 VSS 6.98042e-19 $X=0.033 $Y=0.189
c97 73 VSS 1.35996e-19 $X=0.351 $Y=0.18
c98 69 VSS 7.2814e-19 $X=0.351 $Y=0.134
c99 66 VSS 2.89511e-19 $X=0.189 $Y=0.1665
c100 65 VSS 3.97151e-19 $X=0.189 $Y=0.153
c101 64 VSS 1.55454e-19 $X=0.189 $Y=0.18
c102 59 VSS 0.00360014f $X=0.152 $Y=0.135
c103 58 VSS 4.22838e-19 $X=0.152 $Y=0.135
c104 56 VSS 0.00120122f $X=0.18 $Y=0.135
c105 54 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c106 53 VSS 0.00169428f $X=0.047 $Y=0.234
c107 51 VSS 0.00250477f $X=0.054 $Y=0.234
c108 49 VSS 0.00306385f $X=0.027 $Y=0.234
c109 47 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c110 46 VSS 0.00205521f $X=0.047 $Y=0.036
c111 44 VSS 0.00250477f $X=0.054 $Y=0.036
c112 42 VSS 0.00305101f $X=0.027 $Y=0.036
c113 41 VSS 0.00106422f $X=0.018 $Y=0.225
c114 39 VSS 0.00252163f $X=0.018 $Y=0.1305
c115 38 VSS 0.00142827f $X=0.018 $Y=0.081
c116 37 VSS 0.00214048f $X=0.018 $Y=0.18
c117 34 VSS 0.00507986f $X=0.056 $Y=0.216
c118 31 VSS 2.98509e-19 $X=0.071 $Y=0.216
c119 29 VSS 0.00454717f $X=0.056 $Y=0.054
c120 26 VSS 2.98509e-19 $X=0.071 $Y=0.054
c121 24 VSS 0.00218115f $X=0.464 $Y=0.179
c122 16 VSS 0.059523f $X=0.459 $Y=0.0405
c123 10 VSS 0.0605486f $X=0.351 $Y=0.134
c124 2 VSS 0.0639492f $X=0.135 $Y=0.054
r125 123 124 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.189 $X2=0.1845 $Y2=0.189
r126 122 124 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.189 $X2=0.1845 $Y2=0.189
r127 117 118 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.03 $Y2=0.189
r128 114 117 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.027 $Y2=0.189
r129 108 109 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r130 89 90 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.414
+ $Y=0.189 $X2=0.45 $Y2=0.189
r131 87 90 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.45 $Y2=0.189
r132 87 109 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r133 84 85 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.189 $X2=0.29 $Y2=0.189
r134 82 89 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.414 $Y2=0.189
r135 82 85 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.29 $Y2=0.189
r136 82 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.189 $X2=0.351
+ $Y2=0.189
r137 80 123 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.189 $X2=0.18 $Y2=0.189
r138 79 84 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.162
+ $Y=0.189 $X2=0.229 $Y2=0.189
r139 79 80 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.162 $Y=0.189 $X2=0.162
+ $Y2=0.189
r140 76 118 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.03 $Y2=0.189
r141 75 79 8.75926 $w=1.8e-08 $l=1.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.162 $Y2=0.189
r142 75 76 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.189 $X2=0.033
+ $Y2=0.189
r143 73 83 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.18 $X2=0.351 $Y2=0.189
r144 72 73 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.171 $X2=0.351 $Y2=0.18
r145 69 72 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.134 $X2=0.351 $Y2=0.171
r146 65 66 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.1665
r147 64 122 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.189
r148 64 66 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.1665
r149 63 65 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.153
r150 58 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.152 $Y=0.135 $X2=0.152
+ $Y2=0.135
r151 56 63 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r152 56 58 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.152 $Y2=0.135
r153 53 54 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r154 51 54 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r155 49 53 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r156 46 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r157 44 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r158 42 46 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r159 41 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r160 40 114 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.189
r161 40 41 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.225
r162 38 39 3.36111 $w=1.8e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.1305
r163 37 114 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.189
r164 37 39 3.36111 $w=1.8e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.1305
r165 36 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r166 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r167 34 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r168 31 34 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r169 29 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r170 26 29 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r171 24 108 42.2917 $w=2.4e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.179 $X2=0.513 $Y2=0.179
r172 19 24 3.57143 $w=2.8e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.179 $X2=0.464 $Y2=0.179
r173 16 19 518.891 $w=2e-08 $l=1.385e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.179
r174 10 69 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.134 $X2=0.351
+ $Y2=0.134
r175 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.134 $X2=0.351 $Y2=0.2025
r176 5 59 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.152 $Y2=0.135
r177 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r178 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DHLX1_ASAP7_75T_SRAM%D 2 5 7 11 15 VSS
c18 15 VSS 0.00225715f $X=0.297 $Y=0.135
c19 11 VSS 0.00893359f $X=0.297 $Y=0.1165
c20 5 VSS 0.00197947f $X=0.297 $Y=0.135
c21 2 VSS 0.0613821f $X=0.297 $Y=0.0675
r22 11 15 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1165 $X2=0.297 $Y2=0.135
r23 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r24 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r25 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DHLX1_ASAP7_75T_SRAM%6 2 5 7 9 14 17 19 24 26 31 32 34 37 40 45 55 56 58
+ VSS
c36 58 VSS 8.1019e-19 $X=0.243 $Y=0.2115
c37 56 VSS 4.07532e-19 $X=0.243 $Y=0.126
c38 55 VSS 0.00265408f $X=0.243 $Y=0.117
c39 45 VSS 0.00102494f $X=0.405 $Y=0.134
c40 40 VSS 0.00607715f $X=0.405 $Y=0.153
c41 37 VSS 0.00176992f $X=0.243 $Y=0.153
c42 34 VSS 5.5218e-19 $X=0.243 $Y=0.225
c43 32 VSS 0.00181981f $X=0.216 $Y=0.234
c44 31 VSS 0.0052254f $X=0.198 $Y=0.234
c45 26 VSS 0.00501032f $X=0.234 $Y=0.234
c46 25 VSS 0.00200074f $X=0.216 $Y=0.036
c47 24 VSS 0.00549661f $X=0.198 $Y=0.036
c48 19 VSS 0.00500597f $X=0.234 $Y=0.036
c49 17 VSS 0.00666939f $X=0.16 $Y=0.216
c50 12 VSS 0.00625354f $X=0.16 $Y=0.054
c51 5 VSS 0.0015003f $X=0.405 $Y=0.134
c52 2 VSS 0.059003f $X=0.405 $Y=0.0675
r53 57 58 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.198 $X2=0.243 $Y2=0.2115
r54 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.117 $X2=0.243 $Y2=0.126
r55 41 45 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.405 $Y2=0.134
r56 40 41 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r57 37 57 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.198
r58 37 56 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.126
r59 36 40 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.405 $Y2=0.153
r60 36 37 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.153 $X2=0.243
+ $Y2=0.153
r61 34 58 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.2115
r62 33 55 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.117
r63 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.216 $Y2=0.234
r64 28 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.198 $Y2=0.234
r65 26 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r66 26 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r67 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.216 $Y2=0.036
r68 21 24 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r69 19 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r70 19 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r71 17 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r72 14 17 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r73 12 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r74 9 12 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r75 5 45 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.134 $X2=0.405
+ $Y2=0.134
r76 5 7 357.791 $w=2e-08 $l=9.55e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.134 $X2=0.405 $Y2=0.2295
r77 2 5 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.134
.ends

.subckt PM_DHLX1_ASAP7_75T_SRAM%7 2 5 7 9 12 14 17 21 24 25 29 33 34 36 37 38 39 42
+ 47 48 VSS
c30 48 VSS 0.00241451f $X=0.612 $Y=0.234
c31 47 VSS 0.00236179f $X=0.621 $Y=0.234
c32 42 VSS 0.00170515f $X=0.594 $Y=0.234
c33 40 VSS 4.27948e-19 $X=0.621 $Y=0.216
c34 39 VSS 8.40068e-19 $X=0.621 $Y=0.207
c35 38 VSS 6.87809e-20 $X=0.621 $Y=0.167
c36 37 VSS 7.07046e-19 $X=0.621 $Y=0.164
c37 36 VSS 4.68234e-19 $X=0.621 $Y=0.139
c38 34 VSS 0.00113623f $X=0.621 $Y=0.121
c39 33 VSS 0.00164946f $X=0.621 $Y=0.096
c40 32 VSS 6.22949e-19 $X=0.621 $Y=0.225
c41 30 VSS 7.17067e-19 $X=0.5875 $Y=0.036
c42 29 VSS 0.00656714f $X=0.581 $Y=0.036
c43 25 VSS 0.00222389f $X=0.522 $Y=0.036
c44 24 VSS 0.00488919f $X=0.612 $Y=0.036
c45 21 VSS 5.75409e-19 $X=0.513 $Y=0.082
c46 17 VSS 0.0049422f $X=0.592 $Y=0.2295
c47 12 VSS 0.00511578f $X=0.592 $Y=0.0405
c48 5 VSS 0.00257008f $X=0.513 $Y=0.082
c49 2 VSS 0.058175f $X=0.513 $Y=0.0405
r50 48 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r51 47 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r52 42 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.612 $Y2=0.234
r53 39 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.207 $X2=0.621 $Y2=0.216
r54 38 39 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.207
r55 37 38 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.164 $X2=0.621 $Y2=0.167
r56 36 37 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.139 $X2=0.621 $Y2=0.164
r57 35 36 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.139
r58 34 35 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.121 $X2=0.621 $Y2=0.122
r59 33 34 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.096 $X2=0.621 $Y2=0.121
r60 32 47 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.234
r61 32 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.216
r62 31 33 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.096
r63 29 30 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.581
+ $Y=0.036 $X2=0.5875 $Y2=0.036
r64 27 30 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.5875 $Y2=0.036
r65 25 29 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.581 $Y2=0.036
r66 24 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r67 24 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.594 $Y2=0.036
r68 19 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.513 $Y=0.045 $X2=0.522 $Y2=0.036
r69 19 21 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.082
r70 17 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r71 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r72 12 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036 $X2=0.594
+ $Y2=0.036
r73 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.592 $Y2=0.0405
r74 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.082 $X2=0.513
+ $Y2=0.082
r75 5 7 552.609 $w=2e-08 $l=1.475e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.082 $X2=0.513 $Y2=0.2295
r76 2 5 155.48 $w=2e-08 $l=4.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.082
.ends

.subckt PM_DHLX1_ASAP7_75T_SRAM%8 2 7 10 15 17 22 25 29 30 33 38 39 40 41 42 45 48
+ 49 50 53 55 56 61 64 67 69 70 77 89 90 91 VSS
c61 91 VSS 3.47616e-19 $X=0.459 $Y=0.207
c62 90 VSS 3.33252e-19 $X=0.459 $Y=0.189
c63 89 VSS 1.82803e-20 $X=0.459 $Y=0.171
c64 77 VSS 0.00126446f $X=0.729 $Y=0.136
c65 70 VSS 0.0040364f $X=0.628 $Y=0.153
c66 69 VSS 0.00146526f $X=0.527 $Y=0.153
c67 67 VSS 0.00840598f $X=0.729 $Y=0.153
c68 64 VSS 4.02226e-19 $X=0.459 $Y=0.153
c69 61 VSS 5.11551e-19 $X=0.459 $Y=0.225
c70 60 VSS 2.42691e-19 $X=0.459 $Y=0.13
c71 56 VSS 3.63326e-20 $X=0.522 $Y=0.13
c72 55 VSS 0.00173658f $X=0.504 $Y=0.13
c73 53 VSS 0.00149487f $X=0.567 $Y=0.13
c74 50 VSS 2.19687e-19 $X=0.459 $Y=0.106
c75 49 VSS 3.06086e-19 $X=0.459 $Y=0.096
c76 48 VSS 1.63148e-19 $X=0.459 $Y=0.121
c77 45 VSS 0.00271748f $X=0.432 $Y=0.036
c78 42 VSS 0.00636114f $X=0.45 $Y=0.036
c79 41 VSS 0.00163742f $X=0.432 $Y=0.234
c80 40 VSS 0.00142296f $X=0.414 $Y=0.234
c81 39 VSS 0.00166696f $X=0.396 $Y=0.234
c82 38 VSS 0.00188233f $X=0.379 $Y=0.234
c83 33 VSS 0.00408073f $X=0.45 $Y=0.234
c84 32 VSS 5.7602e-19 $X=0.378 $Y=0.2295
c85 29 VSS 0.00367263f $X=0.378 $Y=0.2025
c86 26 VSS 3.44634e-20 $X=0.3735 $Y=0.216
c87 24 VSS 5.36734e-19 $X=0.432 $Y=0.0405
c88 13 VSS 0.00370005f $X=0.729 $Y=0.136
c89 10 VSS 0.0661232f $X=0.729 $Y=0.0675
c90 5 VSS 0.00267876f $X=0.567 $Y=0.13
c91 2 VSS 0.061627f $X=0.567 $Y=0.0405
r92 90 91 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.189 $X2=0.459 $Y2=0.207
r93 89 90 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.171 $X2=0.459 $Y2=0.189
r94 88 89 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.164 $X2=0.459 $Y2=0.171
r95 69 70 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.628 $Y2=0.153
r96 67 70 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M2 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.628 $Y2=0.153
r97 67 77 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.729 $Y=0.153 $X2=0.729
+ $Y2=0.153
r98 64 88 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.459 $Y2=0.164
r99 63 69 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.527 $Y2=0.153
r100 63 64 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.459 $Y=0.153 $X2=0.459
+ $Y2=0.153
r101 61 91 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.207
r102 59 64 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.139 $X2=0.459 $Y2=0.153
r103 59 60 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.139 $X2=0.459 $Y2=0.13
r104 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.13 $X2=0.522 $Y2=0.13
r105 53 56 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.13 $X2=0.522 $Y2=0.13
r106 51 60 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.13 $X2=0.459 $Y2=0.13
r107 51 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.13 $X2=0.504 $Y2=0.13
r108 49 50 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.096 $X2=0.459 $Y2=0.106
r109 48 60 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.121 $X2=0.459 $Y2=0.13
r110 48 50 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.121 $X2=0.459 $Y2=0.106
r111 47 49 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.096
r112 44 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r113 42 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r114 42 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.432 $Y2=0.036
r115 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.432 $Y2=0.234
r116 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r117 38 39 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.234 $X2=0.396 $Y2=0.234
r118 35 38 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.379 $Y2=0.234
r119 33 61 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r120 33 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.432 $Y2=0.234
r121 30 32 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r122 29 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r123 26 32 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r124 26 29 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r125 25 29 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r126 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r127 21 45 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r128 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r129 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r130 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r131 13 77 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.729 $Y=0.136 $X2=0.729
+ $Y2=0.136
r132 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.136 $X2=0.729 $Y2=0.2025
r133 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.136
r134 5 53 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.13 $X2=0.567
+ $Y2=0.13
r135 5 7 372.777 $w=2e-08 $l=9.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.13 $X2=0.567 $Y2=0.2295
r136 2 5 335.312 $w=2e-08 $l=8.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.13
.ends

.subckt PM_DHLX1_ASAP7_75T_SRAM%Q 1 6 12 14 16 22 30 VSS
c6 30 VSS 0.00433882f $X=0.774 $Y=0.234
c7 29 VSS 0.00278493f $X=0.783 $Y=0.234
c8 22 VSS 0.00433882f $X=0.774 $Y=0.036
c9 21 VSS 0.00278493f $X=0.783 $Y=0.036
c10 19 VSS 0.00641332f $X=0.756 $Y=0.036
c11 16 VSS 0.00208871f $X=0.783 $Y=0.167
c12 14 VSS 0.00372956f $X=0.783 $Y=0.081
c13 12 VSS 0.002726f $X=0.783 $Y=0.225
c14 9 VSS 0.00703052f $X=0.754 $Y=0.2025
c15 4 VSS 3.77696e-19 $X=0.754 $Y=0.0675
r16 30 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.234 $X2=0.7785 $Y2=0.234
r17 29 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.234 $X2=0.7785 $Y2=0.234
r18 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.774 $Y2=0.234
r19 22 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.036 $X2=0.7785 $Y2=0.036
r20 21 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.036 $X2=0.7785 $Y2=0.036
r21 18 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.774 $Y2=0.036
r22 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r23 15 16 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.122 $X2=0.783 $Y2=0.167
r24 14 15 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.081 $X2=0.783 $Y2=0.122
r25 12 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.225 $X2=0.783 $Y2=0.234
r26 12 16 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.225 $X2=0.783 $Y2=0.167
r27 11 21 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.036
r28 11 14 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.081
r29 9 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234 $X2=0.756
+ $Y2=0.234
r30 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.2025 $X2=0.754 $Y2=0.2025
r31 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.756
+ $Y=0.0675 $X2=0.756 $Y2=0.036
r32 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.0675 $X2=0.754 $Y2=0.0675
.ends

.subckt PM_DHLX1_ASAP7_75T_SRAM%10 1 6 9 VSS
c7 9 VSS 0.0266194f $X=0.38 $Y=0.0675
c8 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c9 4 VSS 3.9325e-19 $X=0.322 $Y=0.0675
r10 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r12 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DHLX1_ASAP7_75T_SRAM%11 1 6 9 VSS
c10 9 VSS 0.0211086f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.84146e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DHLX1_ASAP7_75T_SRAM%12 1 2 VSS
c0 1 VSS 0.00220425f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DHLX1_ASAP7_75T_SRAM%13 1 2 VSS
c0 1 VSS 0.00221026f $X=0.341 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends


* END of "./DHLx1_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DHLx1_ASAP7_75t_SRAM  VSS VDD CLK D Q
* 
* Q	Q
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_10_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_6_M3_g N_10_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_12_M4_d N_4_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_12_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_Q_M7_d N_8_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M8 VDD N_CLK_M8_g N_4_M8_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M9 N_6_M9_d N_4_M9_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
M10 N_13_M10_d N_D_M10_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_8_M11_d N_4_M11_g N_13_M11_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M12 N_11_M12_d N_6_M12_g N_8_M12_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M13 VDD N_7_M13_g N_11_M13_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M14 N_7_M14_d N_8_M14_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M15 N_Q_M15_d N_8_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
*
* 
* .include "DHLx1_ASAP7_75t_SRAM.pex.sp.DHLX1_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DHLx1_ASAP7_75t_SRAM.pex.sp.DHLX1_ASAP7_75T_SRAM.pxi"
* File: DHLx1_ASAP7_75t_SRAM.pex.sp.DHLX1_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:27:08 2017
* 
x_PM_DHLX1_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_11_p N_CLK_M8_g CLK N_CLK_c_3_p
+ N_CLK_c_10_p VSS PM_DHLX1_ASAP7_75T_SRAM%CLK
x_PM_DHLX1_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M9_g N_4_c_34_p N_4_M11_g N_4_M4_g
+ N_4_c_88_p N_4_M0_s N_4_c_20_n N_4_M8_s N_4_c_21_n N_4_c_22_n N_4_c_23_n
+ N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_49_p N_4_c_28_n N_4_c_29_n
+ N_4_c_51_p N_4_c_30_n N_4_c_36_p N_4_c_31_n N_4_c_37_p N_4_c_32_n N_4_c_38_p
+ N_4_c_84_p N_4_c_39_p N_4_c_74_p N_4_c_58_p N_4_c_59_p N_4_c_33_n VSS
+ PM_DHLX1_ASAP7_75T_SRAM%4
x_PM_DHLX1_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_104_n N_D_M10_g D N_D_c_111_p VSS
+ PM_DHLX1_ASAP7_75T_SRAM%D
x_PM_DHLX1_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_126_n N_6_M12_g N_6_M1_d N_6_M9_d
+ N_6_c_127_n N_6_c_142_n N_6_c_121_n N_6_c_129_n N_6_c_122_n N_6_c_132_n
+ N_6_c_143_n N_6_c_133_n N_6_c_135_n N_6_c_139_n N_6_c_123_n N_6_c_147_n
+ N_6_c_148_n VSS PM_DHLX1_ASAP7_75T_SRAM%6
x_PM_DHLX1_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_160_n N_7_M13_g N_7_M6_d N_7_c_161_n
+ N_7_M14_d N_7_c_162_n N_7_c_172_p N_7_c_185_p N_7_c_171_p N_7_c_170_p
+ N_7_c_184_p N_7_c_173_p N_7_c_175_p N_7_c_178_p N_7_c_163_n N_7_c_165_n
+ N_7_c_166_n N_7_c_186_p N_7_c_167_n VSS PM_DHLX1_ASAP7_75T_SRAM%7
x_PM_DHLX1_ASAP7_75T_SRAM%8 N_8_M6_g N_8_M14_g N_8_M7_g N_8_M15_g N_8_M3_d N_8_M4_s
+ N_8_M11_d N_8_c_189_n N_8_M12_s N_8_c_244_p N_8_c_191_n N_8_c_192_n
+ N_8_c_219_n N_8_c_193_n N_8_c_194_n N_8_c_195_n N_8_c_196_n N_8_c_197_n
+ N_8_c_198_n N_8_c_199_n N_8_c_200_n N_8_c_201_n N_8_c_247_p N_8_c_202_n
+ N_8_c_233_n N_8_c_204_n N_8_c_234_n N_8_c_237_n N_8_c_207_n N_8_c_209_n
+ N_8_c_212_n VSS PM_DHLX1_ASAP7_75T_SRAM%8
x_PM_DHLX1_ASAP7_75T_SRAM%Q N_Q_M7_d N_Q_M15_d N_Q_c_248_n Q N_Q_c_252_n
+ N_Q_c_250_n N_Q_c_251_n VSS PM_DHLX1_ASAP7_75T_SRAM%Q
x_PM_DHLX1_ASAP7_75T_SRAM%10 N_10_M2_d N_10_M3_s N_10_c_254_n VSS
+ PM_DHLX1_ASAP7_75T_SRAM%10
x_PM_DHLX1_ASAP7_75T_SRAM%11 N_11_M12_d N_11_M13_s N_11_c_262_n VSS
+ PM_DHLX1_ASAP7_75T_SRAM%11
x_PM_DHLX1_ASAP7_75T_SRAM%12 N_12_M5_s N_12_M4_d VSS PM_DHLX1_ASAP7_75T_SRAM%12
x_PM_DHLX1_ASAP7_75T_SRAM%13 N_13_M11_s N_13_M10_d VSS PM_DHLX1_ASAP7_75T_SRAM%13
cc_1 N_CLK_M0_g N_4_M1_g 0.0027643f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_20_n 2.66516e-19 $X=0.08 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 N_CLK_c_3_p N_4_c_21_n 2.48575e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.216
cc_4 N_CLK_c_3_p N_4_c_22_n 0.0020081f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.18
cc_5 CLK N_4_c_23_n 3.98992e-19 $X=0.08 $Y=0.119 $X2=0.018 $Y2=0.081
cc_6 CLK N_4_c_24_n 0.0020081f $X=0.08 $Y=0.119 $X2=0.018 $Y2=0.1305
cc_7 N_CLK_c_3_p N_4_c_25_n 3.00513e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.225
cc_8 CLK N_4_c_26_n 4.98319e-19 $X=0.08 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_3_p N_4_c_27_n 4.98319e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_10_p N_4_c_28_n 4.17e-19 $X=0.081 $Y=0.1305 $X2=0.152 $Y2=0.135
cc_11 N_CLK_c_11_p N_4_c_29_n 0.00111278f $X=0.081 $Y=0.135 $X2=0.152 $Y2=0.135
cc_12 N_CLK_c_3_p N_4_c_30_n 9.46659e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.1665
cc_13 N_CLK_c_3_p N_4_c_31_n 8.7692e-19 $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.189
cc_14 N_CLK_c_3_p N_4_c_32_n 0.00163094f $X=0.081 $Y=0.135 $X2=0.229 $Y2=0.189
cc_15 N_CLK_c_3_p N_4_c_33_n 9.73303e-19 $X=0.081 $Y=0.135 $X2=0.18 $Y2=0.189
cc_16 CLK N_6_c_121_n 6.45949e-19 $X=0.08 $Y=0.119 $X2=0.464 $Y2=0.179
cc_17 N_CLK_c_3_p N_6_c_122_n 6.45949e-19 $X=0.081 $Y=0.135 $X2=0.071 $Y2=0.216
cc_18 CLK N_6_c_123_n 7.98675e-19 $X=0.08 $Y=0.119 $X2=0 $Y2=0
cc_19 N_4_c_34_p N_D_M2_g 0.00341068f $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.054
cc_20 N_4_c_34_p N_D_c_104_n 9.3313e-19 $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.135
cc_21 N_4_c_36_p D 0.00227186f $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.119
cc_22 N_4_c_37_p D 0.00227186f $X=0.351 $Y=0.189 $X2=0.081 $Y2=0.119
cc_23 N_4_c_38_p D 2.29805e-19 $X=0.29 $Y=0.189 $X2=0.081 $Y2=0.119
cc_24 N_4_c_39_p D 6.20826e-19 $X=0.414 $Y=0.189 $X2=0.081 $Y2=0.119
cc_25 N_4_c_34_p N_6_M3_g 0.00355599f $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.054
cc_26 N_4_M4_g N_6_M3_g 0.00355599f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_27 N_4_c_34_p N_6_c_126_n 9.75871e-19 $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.135
cc_28 N_4_c_33_n N_6_c_127_n 0.00154329f $X=0.18 $Y=0.189 $X2=0.081 $Y2=0.1305
cc_29 N_4_c_28_n N_6_c_121_n 9.9131e-19 $X=0.152 $Y=0.135 $X2=0 $Y2=0
cc_30 N_4_c_38_p N_6_c_129_n 4.24027e-19 $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_31 N_4_c_32_n N_6_c_122_n 6.5319e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_32 N_4_c_33_n N_6_c_122_n 0.00305813f $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_33 N_4_c_32_n N_6_c_132_n 4.24027e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_34 N_4_c_49_p N_6_c_133_n 0.00351161f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_35 N_4_c_38_p N_6_c_133_n 0.00102041f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_36 N_4_c_51_p N_6_c_135_n 3.48096e-19 $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_37 N_4_c_36_p N_6_c_135_n 8.9767e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_38 N_4_c_37_p N_6_c_135_n 3.61885e-19 $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_39 N_4_c_38_p N_6_c_135_n 0.0160071f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_40 N_4_c_36_p N_6_c_139_n 0.00286743f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_41 N_4_c_39_p N_6_c_139_n 2.98086e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_42 N_4_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_43 N_4_c_58_p N_7_M5_g 0.00199227f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_44 N_4_c_59_p N_7_M5_g 5.16754e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_45 N_4_c_58_p N_7_c_160_n 4.44235e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.135
cc_46 N_4_c_58_p N_7_c_161_n 5.31675e-19 $X=0.513 $Y=0.18 $X2=0.08 $Y2=0.119
cc_47 N_4_c_58_p N_7_c_162_n 0.00169036f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.1305
cc_48 N_4_c_58_p N_7_c_163_n 6.34096e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_49 N_4_c_59_p N_7_c_163_n 7.16706e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_50 N_4_c_58_p N_7_c_165_n 0.0026997f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_51 N_4_c_58_p N_7_c_166_n 3.09575e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_52 N_4_c_58_p N_7_c_167_n 2.32568e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_53 N_4_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_54 N_4_c_58_p N_8_M6_g 0.00305656f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_55 N_4_c_36_p N_8_c_189_n 9.02348e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_56 N_4_c_37_p N_8_c_189_n 0.00144031f $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_57 N_4_c_37_p N_8_c_191_n 0.00138499f $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_58 N_4_c_39_p N_8_c_192_n 6.75805e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_59 N_4_c_74_p N_8_c_193_n 6.75805e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_60 N_4_c_74_p N_8_c_194_n 3.48842e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_61 N_4_c_74_p N_8_c_195_n 2.01793e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_62 N_4_M4_g N_8_c_196_n 2.73971e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_63 N_4_M4_g N_8_c_197_n 3.60498e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_64 N_4_M4_g N_8_c_198_n 2.06358e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_65 N_4_c_58_p N_8_c_199_n 4.82796e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_66 N_4_c_58_p N_8_c_200_n 7.81688e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_67 N_4_c_59_p N_8_c_201_n 0.001012f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_68 N_4_M4_g N_8_c_202_n 2.17193e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_69 N_4_c_84_p N_8_c_202_n 2.46239e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_70 N_4_c_84_p N_8_c_204_n 0.00694522f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_71 N_4_c_58_p N_8_c_204_n 0.00195859f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_72 N_4_c_59_p N_8_c_204_n 2.84813e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_73 N_4_c_88_p N_8_c_207_n 0.00127126f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_74 N_4_c_59_p N_8_c_207_n 0.00199566f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_75 N_4_c_88_p N_8_c_209_n 0.0011121f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_76 N_4_c_84_p N_8_c_209_n 3.67862e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_77 N_4_c_58_p N_8_c_209_n 4.28262e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_78 N_4_c_88_p N_8_c_212_n 7.05645e-19 $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_79 N_4_c_37_p N_8_c_212_n 2.96264e-19 $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_80 N_4_c_84_p N_8_c_212_n 3.05556e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_81 N_4_c_34_p N_10_c_254_n 0.00650944f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_82 N_4_c_36_p N_10_c_254_n 0.00135463f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_83 N_4_c_58_p N_11_M13_s 2.34172e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.216
cc_84 N_4_M4_g N_11_c_262_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_85 N_4_c_88_p N_11_c_262_n 0.0013957f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_86 N_4_c_74_p N_11_c_262_n 7.09553e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_87 N_4_c_58_p N_11_c_262_n 0.00230217f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_88 N_D_M2_g N_6_M3_g 2.82885e-19 $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_89 D N_6_c_142_n 0.00128741f $X=0.297 $Y=0.1165 $X2=0.459 $Y2=0.179
cc_90 N_D_c_111_p N_6_c_143_n 0.00128741f $X=0.297 $Y=0.135 $X2=0.056 $Y2=0.216
cc_91 D N_6_c_133_n 0.00138082f $X=0.297 $Y=0.1165 $X2=0.018 $Y2=0.18
cc_92 D N_6_c_135_n 0.0012236f $X=0.297 $Y=0.1165 $X2=0.018 $Y2=0.198
cc_93 D N_6_c_123_n 0.00128741f $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_94 D N_6_c_147_n 0.00128741f $X=0.297 $Y=0.1165 $X2=0.18 $Y2=0.135
cc_95 N_D_c_111_p N_6_c_148_n 0.00128741f $X=0.297 $Y=0.135 $X2=0.152 $Y2=0.135
cc_96 N_D_c_111_p N_8_c_189_n 3.23895e-19 $X=0.297 $Y=0.135 $X2=0.056 $Y2=0.054
cc_97 N_D_c_111_p N_8_c_191_n 3.35757e-19 $X=0.297 $Y=0.135 $X2=0.018 $Y2=0.081
cc_98 D N_8_c_194_n 2.05539e-19 $X=0.297 $Y=0.1165 $X2=0.027 $Y2=0.036
cc_99 D N_10_c_254_n 0.00445409f $X=0.297 $Y=0.1165 $X2=0.351 $Y2=0.134
cc_100 N_6_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_101 N_6_c_139_n N_8_c_189_n 4.65343e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_102 N_6_M3_g N_8_c_219_n 3.33314e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_103 N_6_c_139_n N_8_c_219_n 4.18821e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_104 N_6_c_139_n N_8_c_196_n 0.00307076f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_105 N_6_c_139_n N_8_c_202_n 2.60642e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_106 N_6_c_135_n N_8_c_204_n 8.88396e-19 $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_107 N_6_c_135_n N_10_c_254_n 8.35084e-19 $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_108 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_109 N_7_c_170_p N_8_M6_g 3.83894e-19 $X=0.581 $Y=0.036 $X2=0.135 $Y2=0.054
cc_110 N_7_c_171_p N_8_c_194_n 0.0017541f $X=0.522 $Y=0.036 $X2=0.027 $Y2=0.036
cc_111 N_7_c_172_p N_8_c_197_n 0.0017541f $X=0.513 $Y=0.082 $X2=0.027 $Y2=0.234
cc_112 N_7_c_173_p N_8_c_198_n 2.88106e-19 $X=0.621 $Y=0.121 $X2=0.054 $Y2=0.234
cc_113 N_7_c_170_p N_8_c_199_n 7.32482e-19 $X=0.581 $Y=0.036 $X2=0.047 $Y2=0.234
cc_114 N_7_c_175_p N_8_c_199_n 9.52305e-19 $X=0.621 $Y=0.139 $X2=0.047 $Y2=0.234
cc_115 N_7_M5_g N_8_c_201_n 4.16078e-19 $X=0.513 $Y=0.0405 $X2=0.18 $Y2=0.135
cc_116 N_7_c_172_p N_8_c_201_n 0.00115865f $X=0.513 $Y=0.082 $X2=0.18 $Y2=0.135
cc_117 N_7_c_178_p N_8_c_233_n 3.90412e-19 $X=0.621 $Y=0.164 $X2=0.351 $Y2=0.189
cc_118 N_7_c_161_n N_8_c_234_n 2.11538e-19 $X=0.592 $Y=0.0405 $X2=0.351
+ $Y2=0.134
cc_119 N_7_c_178_p N_8_c_234_n 8.8208e-19 $X=0.621 $Y=0.164 $X2=0.351 $Y2=0.134
cc_120 N_7_c_166_n N_8_c_234_n 5.92034e-19 $X=0.594 $Y=0.234 $X2=0.351 $Y2=0.134
cc_121 N_7_c_175_p N_8_c_237_n 6.03721e-19 $X=0.621 $Y=0.139 $X2=0 $Y2=0
cc_122 N_7_c_165_n N_Q_c_248_n 3.1718e-19 $X=0.621 $Y=0.207 $X2=0.351 $Y2=0.2025
cc_123 N_7_c_184_p Q 3.1718e-19 $X=0.621 $Y=0.096 $X2=0 $Y2=0
cc_124 N_7_c_185_p N_Q_c_250_n 2.22376e-19 $X=0.612 $Y=0.036 $X2=0 $Y2=0
cc_125 N_7_c_186_p N_Q_c_251_n 2.15386e-19 $X=0.621 $Y=0.234 $X2=0 $Y2=0
cc_126 N_8_c_233_n N_Q_c_252_n 2.31367e-19 $X=0.729 $Y=0.153 $X2=0.459
+ $Y2=0.0405
cc_127 N_8_c_237_n N_Q_c_252_n 0.00212036f $X=0.729 $Y=0.136 $X2=0.459
+ $Y2=0.0405
cc_128 N_8_c_189_n N_10_c_254_n 0.00119601f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.134
cc_129 N_8_c_194_n N_10_c_254_n 4.50844e-19 $X=0.45 $Y=0.036 $X2=0.351 $Y2=0.134
cc_130 N_8_c_195_n N_10_c_254_n 0.00394776f $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.134
cc_131 N_8_c_189_n N_11_c_262_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.134
cc_132 N_8_c_244_p N_11_c_262_n 0.00222776f $X=0.45 $Y=0.234 $X2=0.351 $Y2=0.134
cc_133 N_8_c_193_n N_11_c_262_n 0.00118584f $X=0.432 $Y=0.234 $X2=0.351
+ $Y2=0.134
cc_134 N_8_c_195_n N_11_c_262_n 5.72355e-19 $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.134
cc_135 N_8_c_247_p N_11_c_262_n 0.00116187f $X=0.459 $Y=0.225 $X2=0.351
+ $Y2=0.134

* END of "./DHLx1_ASAP7_75t_SRAM.pex.sp.DHLX1_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DHLx2_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:27:30 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DHLx2_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DHLx2_ASAP7_75t_SRAM.pex.sp.pex"
* File: DHLx2_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:27:30 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DHLX2_ASAP7_75T_SRAM%CLK 2 5 7 12 14 17 VSS
c18 17 VSS 5.41721e-21 $X=0.081 $Y=0.1305
c19 14 VSS 0.00699913f $X=0.081 $Y=0.135
c20 12 VSS 0.00699194f $X=0.08 $Y=0.119
c21 5 VSS 0.00183412f $X=0.081 $Y=0.135
c22 2 VSS 0.062963f $X=0.081 $Y=0.054
r23 16 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r24 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r25 12 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.126
r26 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DHLX2_ASAP7_75T_SRAM%4 2 7 10 13 16 24 26 29 31 34 37 38 39 41 44 51 56
+ 58 59 65 66 69 76 83 84 85 87 89 90 108 109 123 VSS
c83 123 VSS 5.19505e-19 $X=0.18 $Y=0.189
c84 122 VSS 1.53285e-19 $X=0.189 $Y=0.189
c85 118 VSS 7.0154e-20 $X=0.03 $Y=0.189
c86 117 VSS 5.9624e-19 $X=0.027 $Y=0.189
c87 109 VSS 7.76097e-19 $X=0.513 $Y=0.18
c88 108 VSS 0.0574514f $X=0.513 $Y=0.18
c89 90 VSS 0.00123576f $X=0.45 $Y=0.189
c90 89 VSS 0.0038091f $X=0.414 $Y=0.189
c91 87 VSS 0.00305138f $X=0.513 $Y=0.189
c92 85 VSS 0.00251877f $X=0.29 $Y=0.189
c93 84 VSS 0.00700382f $X=0.229 $Y=0.189
c94 83 VSS 0.00149088f $X=0.351 $Y=0.189
c95 76 VSS 6.98042e-19 $X=0.033 $Y=0.189
c96 73 VSS 1.35996e-19 $X=0.351 $Y=0.18
c97 69 VSS 7.2814e-19 $X=0.351 $Y=0.134
c98 66 VSS 2.89511e-19 $X=0.189 $Y=0.1665
c99 65 VSS 3.97151e-19 $X=0.189 $Y=0.153
c100 64 VSS 1.55454e-19 $X=0.189 $Y=0.18
c101 59 VSS 0.00360014f $X=0.152 $Y=0.135
c102 58 VSS 4.22838e-19 $X=0.152 $Y=0.135
c103 56 VSS 0.00120122f $X=0.18 $Y=0.135
c104 54 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c105 53 VSS 0.00169428f $X=0.047 $Y=0.234
c106 51 VSS 0.00250477f $X=0.054 $Y=0.234
c107 49 VSS 0.00306385f $X=0.027 $Y=0.234
c108 47 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c109 46 VSS 0.00205521f $X=0.047 $Y=0.036
c110 44 VSS 0.00250477f $X=0.054 $Y=0.036
c111 42 VSS 0.00305101f $X=0.027 $Y=0.036
c112 41 VSS 0.00106422f $X=0.018 $Y=0.225
c113 39 VSS 0.00252163f $X=0.018 $Y=0.1305
c114 38 VSS 0.00142827f $X=0.018 $Y=0.081
c115 37 VSS 0.00214048f $X=0.018 $Y=0.18
c116 34 VSS 0.00507986f $X=0.056 $Y=0.216
c117 31 VSS 2.98509e-19 $X=0.071 $Y=0.216
c118 29 VSS 0.00454717f $X=0.056 $Y=0.054
c119 26 VSS 2.98509e-19 $X=0.071 $Y=0.054
c120 24 VSS 0.00218115f $X=0.464 $Y=0.179
c121 16 VSS 0.059523f $X=0.459 $Y=0.0405
c122 10 VSS 0.0605486f $X=0.351 $Y=0.134
c123 2 VSS 0.0627154f $X=0.135 $Y=0.054
r124 123 124 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.189 $X2=0.1845 $Y2=0.189
r125 122 124 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.189 $X2=0.1845 $Y2=0.189
r126 117 118 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.03 $Y2=0.189
r127 114 117 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.027 $Y2=0.189
r128 108 109 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r129 89 90 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.414
+ $Y=0.189 $X2=0.45 $Y2=0.189
r130 87 90 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.45 $Y2=0.189
r131 87 109 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r132 84 85 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.189 $X2=0.29 $Y2=0.189
r133 82 89 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.414 $Y2=0.189
r134 82 85 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.29 $Y2=0.189
r135 82 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.189 $X2=0.351
+ $Y2=0.189
r136 80 123 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.189 $X2=0.18 $Y2=0.189
r137 79 84 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.162
+ $Y=0.189 $X2=0.229 $Y2=0.189
r138 79 80 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.162 $Y=0.189 $X2=0.162
+ $Y2=0.189
r139 76 118 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.03 $Y2=0.189
r140 75 79 8.75926 $w=1.8e-08 $l=1.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.162 $Y2=0.189
r141 75 76 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.189 $X2=0.033
+ $Y2=0.189
r142 73 83 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.18 $X2=0.351 $Y2=0.189
r143 72 73 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.171 $X2=0.351 $Y2=0.18
r144 69 72 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.134 $X2=0.351 $Y2=0.171
r145 65 66 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.1665
r146 64 122 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.189
r147 64 66 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.1665
r148 63 65 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.153
r149 58 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.152 $Y=0.135 $X2=0.152
+ $Y2=0.135
r150 56 63 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r151 56 58 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.152 $Y2=0.135
r152 53 54 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r153 51 54 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r154 49 53 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r155 46 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r156 44 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r157 42 46 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r158 41 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r159 40 114 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.189
r160 40 41 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.225
r161 38 39 3.36111 $w=1.8e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.1305
r162 37 114 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.189
r163 37 39 3.36111 $w=1.8e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.1305
r164 36 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r165 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r166 34 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r167 31 34 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r168 29 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r169 26 29 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r170 24 108 42.2917 $w=2.4e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.179 $X2=0.513 $Y2=0.179
r171 19 24 3.57143 $w=2.8e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.179 $X2=0.464 $Y2=0.179
r172 16 19 518.891 $w=2e-08 $l=1.385e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.179
r173 10 69 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.134 $X2=0.351
+ $Y2=0.134
r174 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.134 $X2=0.351 $Y2=0.2025
r175 5 59 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.152 $Y2=0.135
r176 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r177 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DHLX2_ASAP7_75T_SRAM%D 2 5 7 11 15 VSS
c18 15 VSS 0.00225715f $X=0.297 $Y=0.135
c19 11 VSS 0.00893359f $X=0.297 $Y=0.1165
c20 5 VSS 0.00197947f $X=0.297 $Y=0.135
c21 2 VSS 0.0613821f $X=0.297 $Y=0.0675
r22 11 15 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1165 $X2=0.297 $Y2=0.135
r23 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r24 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r25 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DHLX2_ASAP7_75T_SRAM%6 2 5 7 9 14 17 19 24 26 31 32 34 37 40 45 55 56 58
+ VSS
c36 58 VSS 8.1019e-19 $X=0.243 $Y=0.2115
c37 56 VSS 4.07532e-19 $X=0.243 $Y=0.126
c38 55 VSS 0.00265408f $X=0.243 $Y=0.117
c39 45 VSS 0.00102515f $X=0.405 $Y=0.134
c40 40 VSS 0.00607715f $X=0.405 $Y=0.153
c41 37 VSS 0.00176992f $X=0.243 $Y=0.153
c42 34 VSS 5.5218e-19 $X=0.243 $Y=0.225
c43 32 VSS 0.00181981f $X=0.216 $Y=0.234
c44 31 VSS 0.0052254f $X=0.198 $Y=0.234
c45 26 VSS 0.00501032f $X=0.234 $Y=0.234
c46 25 VSS 0.00200074f $X=0.216 $Y=0.036
c47 24 VSS 0.00549661f $X=0.198 $Y=0.036
c48 19 VSS 0.00500597f $X=0.234 $Y=0.036
c49 17 VSS 0.00666939f $X=0.16 $Y=0.216
c50 12 VSS 0.00625354f $X=0.16 $Y=0.054
c51 5 VSS 0.0015003f $X=0.405 $Y=0.134
c52 2 VSS 0.059003f $X=0.405 $Y=0.0675
r53 57 58 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.198 $X2=0.243 $Y2=0.2115
r54 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.117 $X2=0.243 $Y2=0.126
r55 41 45 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.405 $Y2=0.134
r56 40 41 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r57 37 57 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.198
r58 37 56 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.126
r59 36 40 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.405 $Y2=0.153
r60 36 37 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.153 $X2=0.243
+ $Y2=0.153
r61 34 58 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.2115
r62 33 55 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.117
r63 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.216 $Y2=0.234
r64 28 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.198 $Y2=0.234
r65 26 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r66 26 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r67 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.216 $Y2=0.036
r68 21 24 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r69 19 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r70 19 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r71 17 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r72 14 17 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r73 12 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r74 9 12 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r75 5 45 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.134 $X2=0.405
+ $Y2=0.134
r76 5 7 357.791 $w=2e-08 $l=9.55e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.134 $X2=0.405 $Y2=0.2295
r77 2 5 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.134
.ends

.subckt PM_DHLX2_ASAP7_75T_SRAM%7 2 5 7 9 12 14 17 21 25 29 35 36 37 38 39 40 44 50
+ VSS
c25 50 VSS 0.00241451f $X=0.612 $Y=0.234
c26 49 VSS 0.00242518f $X=0.621 $Y=0.234
c27 44 VSS 0.00170515f $X=0.594 $Y=0.234
c28 42 VSS 4.20115e-19 $X=0.621 $Y=0.2205
c29 41 VSS 3.42267e-19 $X=0.621 $Y=0.216
c30 40 VSS 0.00103787f $X=0.621 $Y=0.207
c31 39 VSS 5.73174e-20 $X=0.621 $Y=0.167
c32 38 VSS 7.19987e-19 $X=0.621 $Y=0.164
c33 37 VSS 4.79275e-19 $X=0.621 $Y=0.139
c34 36 VSS 0.00102697f $X=0.621 $Y=0.121
c35 35 VSS 1.81917e-19 $X=0.621 $Y=0.096
c36 34 VSS 0.0014183f $X=0.621 $Y=0.09
c37 33 VSS 2.06522e-19 $X=0.621 $Y=0.054
c38 32 VSS 4.87482e-19 $X=0.621 $Y=0.225
c39 30 VSS 7.17067e-19 $X=0.5875 $Y=0.036
c40 29 VSS 0.00656714f $X=0.581 $Y=0.036
c41 25 VSS 0.00222389f $X=0.522 $Y=0.036
c42 24 VSS 0.00513623f $X=0.612 $Y=0.036
c43 21 VSS 5.75409e-19 $X=0.513 $Y=0.082
c44 17 VSS 0.00494219f $X=0.592 $Y=0.2295
c45 12 VSS 0.00511578f $X=0.592 $Y=0.0405
c46 5 VSS 0.00257008f $X=0.513 $Y=0.082
c47 2 VSS 0.058175f $X=0.513 $Y=0.0405
r48 50 51 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r49 49 51 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r50 44 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.612 $Y2=0.234
r51 41 42 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.216 $X2=0.621 $Y2=0.2205
r52 40 41 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.207 $X2=0.621 $Y2=0.216
r53 39 40 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.207
r54 38 39 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.164 $X2=0.621 $Y2=0.167
r55 37 38 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.139 $X2=0.621 $Y2=0.164
r56 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.121 $X2=0.621 $Y2=0.139
r57 35 36 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.096 $X2=0.621 $Y2=0.121
r58 34 35 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.621 $Y2=0.096
r59 33 34 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.054 $X2=0.621 $Y2=0.09
r60 32 49 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.234
r61 32 42 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.2205
r62 31 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.054
r63 29 30 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.581
+ $Y=0.036 $X2=0.5875 $Y2=0.036
r64 27 30 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.5875 $Y2=0.036
r65 25 29 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.581 $Y2=0.036
r66 24 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r67 24 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.594 $Y2=0.036
r68 19 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.513 $Y=0.045 $X2=0.522 $Y2=0.036
r69 19 21 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.082
r70 17 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r71 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r72 12 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036 $X2=0.594
+ $Y2=0.036
r73 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.592 $Y2=0.0405
r74 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.082 $X2=0.513
+ $Y2=0.082
r75 5 7 552.609 $w=2e-08 $l=1.475e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.082 $X2=0.513 $Y2=0.2295
r76 2 5 155.48 $w=2e-08 $l=4.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.082
.ends

.subckt PM_DHLX2_ASAP7_75T_SRAM%8 2 7 10 15 18 23 25 30 33 37 38 41 46 47 48 49 50
+ 53 56 57 58 61 63 64 69 72 77 78 80 88 93 105 106 107 VSS
c71 107 VSS 3.47616e-19 $X=0.459 $Y=0.207
c72 106 VSS 3.33252e-19 $X=0.459 $Y=0.189
c73 105 VSS 1.82803e-20 $X=0.459 $Y=0.171
c74 93 VSS 0.00121597f $X=0.783 $Y=0.136
c75 88 VSS 0.00219093f $X=0.729 $Y=0.136
c76 80 VSS 0.00985038f $X=0.783 $Y=0.153
c77 78 VSS 0.0040364f $X=0.628 $Y=0.153
c78 77 VSS 0.00146547f $X=0.527 $Y=0.153
c79 72 VSS 4.01751e-19 $X=0.459 $Y=0.153
c80 69 VSS 5.11076e-19 $X=0.459 $Y=0.225
c81 68 VSS 2.42691e-19 $X=0.459 $Y=0.13
c82 64 VSS 3.63326e-20 $X=0.522 $Y=0.13
c83 63 VSS 0.00173658f $X=0.504 $Y=0.13
c84 61 VSS 0.00150363f $X=0.567 $Y=0.13
c85 58 VSS 2.19687e-19 $X=0.459 $Y=0.106
c86 57 VSS 3.06086e-19 $X=0.459 $Y=0.096
c87 56 VSS 1.63148e-19 $X=0.459 $Y=0.121
c88 53 VSS 0.00271748f $X=0.432 $Y=0.036
c89 50 VSS 0.00636114f $X=0.45 $Y=0.036
c90 49 VSS 0.00163742f $X=0.432 $Y=0.234
c91 48 VSS 0.00142296f $X=0.414 $Y=0.234
c92 47 VSS 0.00166696f $X=0.396 $Y=0.234
c93 46 VSS 0.00188233f $X=0.379 $Y=0.234
c94 41 VSS 0.00408073f $X=0.45 $Y=0.234
c95 40 VSS 5.7602e-19 $X=0.378 $Y=0.2295
c96 37 VSS 0.00367263f $X=0.378 $Y=0.2025
c97 34 VSS 3.44634e-20 $X=0.3735 $Y=0.216
c98 32 VSS 5.36734e-19 $X=0.432 $Y=0.0405
c99 21 VSS 0.00232571f $X=0.783 $Y=0.136
c100 18 VSS 0.0609548f $X=0.783 $Y=0.0675
c101 13 VSS 0.00318825f $X=0.729 $Y=0.136
c102 10 VSS 0.0612321f $X=0.729 $Y=0.0675
c103 5 VSS 0.00268089f $X=0.567 $Y=0.13
c104 2 VSS 0.061627f $X=0.567 $Y=0.0405
r105 106 107 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.189 $X2=0.459 $Y2=0.207
r106 105 106 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.171 $X2=0.459 $Y2=0.189
r107 104 105 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.164 $X2=0.459 $Y2=0.171
r108 80 93 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.783 $Y=0.153 $X2=0.783
+ $Y2=0.153
r109 77 78 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.628 $Y2=0.153
r110 75 80 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.783 $Y2=0.153
r111 75 78 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M2 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.628 $Y2=0.153
r112 75 88 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.729 $Y=0.153 $X2=0.729
+ $Y2=0.153
r113 72 104 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.459 $Y2=0.164
r114 71 77 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.527 $Y2=0.153
r115 71 72 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.459 $Y=0.153 $X2=0.459
+ $Y2=0.153
r116 69 107 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.207
r117 67 72 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.139 $X2=0.459 $Y2=0.153
r118 67 68 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.139 $X2=0.459 $Y2=0.13
r119 63 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.13 $X2=0.522 $Y2=0.13
r120 61 64 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.13 $X2=0.522 $Y2=0.13
r121 59 68 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.13 $X2=0.459 $Y2=0.13
r122 59 63 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.13 $X2=0.504 $Y2=0.13
r123 57 58 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.096 $X2=0.459 $Y2=0.106
r124 56 68 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.121 $X2=0.459 $Y2=0.13
r125 56 58 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.121 $X2=0.459 $Y2=0.106
r126 55 57 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.096
r127 52 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r128 50 55 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r129 50 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.432 $Y2=0.036
r130 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.432 $Y2=0.234
r131 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r132 46 47 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.234 $X2=0.396 $Y2=0.234
r133 43 46 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.379 $Y2=0.234
r134 41 69 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r135 41 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.432 $Y2=0.234
r136 38 40 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r137 37 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r138 34 40 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r139 34 37 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r140 33 37 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r141 30 32 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r142 29 53 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r143 26 32 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r144 26 29 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r145 25 29 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r146 21 93 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.136 $X2=0.783
+ $Y2=0.136
r147 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.136 $X2=0.783 $Y2=0.2025
r148 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.136
r149 13 88 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.729 $Y=0.136 $X2=0.729
+ $Y2=0.136
r150 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.136 $X2=0.729 $Y2=0.2025
r151 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.136
r152 5 61 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.13 $X2=0.567
+ $Y2=0.13
r153 5 7 372.777 $w=2e-08 $l=9.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.13 $X2=0.567 $Y2=0.2295
r154 2 5 335.312 $w=2e-08 $l=8.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.13
.ends

.subckt PM_DHLX2_ASAP7_75T_SRAM%Q 1 2 6 7 10 13 19 23 25 26 30 32 VSS
c12 34 VSS 0.00149303f $X=0.841 $Y=0.1915
c13 32 VSS 6.40338e-19 $X=0.841 $Y=0.103
c14 31 VSS 0.00187702f $X=0.841 $Y=0.09
c15 30 VSS 0.00318964f $X=0.841 $Y=0.116
c16 28 VSS 0.00116885f $X=0.841 $Y=0.216
c17 26 VSS 9.95001e-19 $X=0.792 $Y=0.045
c18 25 VSS 0.00317904f $X=0.774 $Y=0.045
c19 23 VSS 0.00776403f $X=0.756 $Y=0.045
c20 20 VSS 0.00817147f $X=0.832 $Y=0.045
c21 19 VSS 9.93081e-19 $X=0.792 $Y=0.225
c22 18 VSS 0.00169843f $X=0.774 $Y=0.225
c23 13 VSS 0.00145993f $X=0.756 $Y=0.225
c24 11 VSS 0.00819723f $X=0.832 $Y=0.225
c25 10 VSS 0.00750057f $X=0.756 $Y=0.2025
c26 6 VSS 7.42424e-19 $X=0.773 $Y=0.2025
c27 1 VSS 7.38823e-19 $X=0.773 $Y=0.0675
r28 33 34 1.66358 $w=1.8e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.841
+ $Y=0.167 $X2=0.841 $Y2=0.1915
r29 31 32 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.841
+ $Y=0.09 $X2=0.841 $Y2=0.103
r30 30 33 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.841
+ $Y=0.116 $X2=0.841 $Y2=0.167
r31 30 32 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.841
+ $Y=0.116 $X2=0.841 $Y2=0.103
r32 28 34 1.66358 $w=1.8e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.841
+ $Y=0.216 $X2=0.841 $Y2=0.1915
r33 27 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.841
+ $Y=0.054 $X2=0.841 $Y2=0.09
r34 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.045 $X2=0.792 $Y2=0.045
r35 22 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.045 $X2=0.774 $Y2=0.045
r36 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.045 $X2=0.756
+ $Y2=0.045
r37 20 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.832 $Y=0.045 $X2=0.841 $Y2=0.054
r38 20 26 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.832
+ $Y=0.045 $X2=0.792 $Y2=0.045
r39 18 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.225 $X2=0.792 $Y2=0.225
r40 13 18 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.225 $X2=0.774 $Y2=0.225
r41 11 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.832 $Y=0.225 $X2=0.841 $Y2=0.216
r42 11 19 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.832
+ $Y=0.225 $X2=0.792 $Y2=0.225
r43 10 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.225 $X2=0.756
+ $Y2=0.225
r44 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r45 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r46 5 23 19.4196 $w=2.4e-08 $l=2.25e-08 $layer=LISD $thickness=2.8e-08 $X=0.756
+ $Y=0.0675 $X2=0.756 $Y2=0.045
r47 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
r48 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
.ends

.subckt PM_DHLX2_ASAP7_75T_SRAM%10 1 6 9 VSS
c7 9 VSS 0.0266194f $X=0.38 $Y=0.0675
c8 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c9 4 VSS 3.9325e-19 $X=0.322 $Y=0.0675
r10 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r12 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DHLX2_ASAP7_75T_SRAM%11 1 6 9 VSS
c10 9 VSS 0.0211086f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.84146e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DHLX2_ASAP7_75T_SRAM%12 1 2 VSS
c0 1 VSS 0.00220425f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DHLX2_ASAP7_75T_SRAM%13 1 2 VSS
c0 1 VSS 0.00221026f $X=0.341 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends


* END of "./DHLx2_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DHLx2_ASAP7_75t_SRAM  VSS VDD CLK D Q
* 
* Q	Q
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_10_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_6_M3_g N_10_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_12_M4_d N_4_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_12_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_Q_M7_d N_8_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M8 N_Q_M8_d N_8_M8_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773 $Y=0.027
M9 VDD N_CLK_M9_g N_4_M9_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M10 N_6_M10_d N_4_M10_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M11 N_13_M11_d N_D_M11_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M12 N_8_M12_d N_4_M12_g N_13_M12_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M13 N_11_M13_d N_6_M13_g N_8_M13_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M14 VDD N_7_M14_g N_11_M14_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M15 N_7_M15_d N_8_M15_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M16 N_Q_M16_d N_8_M16_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M17 N_Q_M17_d N_8_M17_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
*
* 
* .include "DHLx2_ASAP7_75t_SRAM.pex.sp.DHLX2_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DHLx2_ASAP7_75t_SRAM.pex.sp.DHLX2_ASAP7_75T_SRAM.pxi"
* File: DHLx2_ASAP7_75t_SRAM.pex.sp.DHLX2_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:27:30 2017
* 
x_PM_DHLX2_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_11_p N_CLK_M9_g CLK N_CLK_c_3_p
+ N_CLK_c_10_p VSS PM_DHLX2_ASAP7_75T_SRAM%CLK
x_PM_DHLX2_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M10_g N_4_c_34_p N_4_M12_g N_4_M4_g
+ N_4_c_87_p N_4_M0_s N_4_c_20_n N_4_M9_s N_4_c_21_n N_4_c_22_n N_4_c_23_n
+ N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_49_p N_4_c_28_n N_4_c_29_n
+ N_4_c_51_p N_4_c_30_n N_4_c_36_p N_4_c_31_n N_4_c_37_p N_4_c_32_n N_4_c_38_p
+ N_4_c_83_p N_4_c_39_p N_4_c_73_p N_4_c_58_p N_4_c_59_p N_4_c_33_n VSS
+ PM_DHLX2_ASAP7_75T_SRAM%4
x_PM_DHLX2_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_103_n N_D_M11_g D N_D_c_110_p VSS
+ PM_DHLX2_ASAP7_75T_SRAM%D
x_PM_DHLX2_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_125_n N_6_M13_g N_6_M1_d N_6_M10_d
+ N_6_c_126_n N_6_c_141_n N_6_c_120_n N_6_c_128_n N_6_c_121_n N_6_c_131_n
+ N_6_c_142_n N_6_c_132_n N_6_c_134_n N_6_c_138_n N_6_c_122_n N_6_c_146_n
+ N_6_c_147_n VSS PM_DHLX2_ASAP7_75T_SRAM%6
x_PM_DHLX2_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_159_n N_7_M14_g N_7_M6_d N_7_c_160_n
+ N_7_M15_d N_7_c_161_n N_7_c_170_p N_7_c_169_p N_7_c_168_p N_7_c_180_p
+ N_7_c_171_p N_7_c_173_p N_7_c_177_p N_7_c_162_n N_7_c_163_n N_7_c_164_n
+ N_7_c_165_n VSS PM_DHLX2_ASAP7_75T_SRAM%7
x_PM_DHLX2_ASAP7_75T_SRAM%8 N_8_M6_g N_8_M15_g N_8_M7_g N_8_M16_g N_8_M8_g
+ N_8_M17_g N_8_M3_d N_8_M4_s N_8_M12_d N_8_c_183_n N_8_M13_s N_8_c_248_p
+ N_8_c_185_n N_8_c_186_n N_8_c_213_n N_8_c_187_n N_8_c_188_n N_8_c_189_n
+ N_8_c_190_n N_8_c_191_n N_8_c_192_n N_8_c_193_n N_8_c_194_n N_8_c_195_n
+ N_8_c_251_p N_8_c_196_n N_8_c_198_n N_8_c_227_n N_8_c_230_n N_8_c_231_n
+ N_8_c_235_p N_8_c_201_n N_8_c_203_n N_8_c_206_n VSS PM_DHLX2_ASAP7_75T_SRAM%8
x_PM_DHLX2_ASAP7_75T_SRAM%Q N_Q_M8_d N_Q_M7_d N_Q_M17_d N_Q_M16_d N_Q_c_252_n
+ N_Q_c_253_n N_Q_c_254_n N_Q_c_256_n N_Q_c_259_n N_Q_c_260_n Q N_Q_c_263_n VSS
+ PM_DHLX2_ASAP7_75T_SRAM%Q
x_PM_DHLX2_ASAP7_75T_SRAM%10 N_10_M2_d N_10_M3_s N_10_c_264_n VSS
+ PM_DHLX2_ASAP7_75T_SRAM%10
x_PM_DHLX2_ASAP7_75T_SRAM%11 N_11_M13_d N_11_M14_s N_11_c_272_n VSS
+ PM_DHLX2_ASAP7_75T_SRAM%11
x_PM_DHLX2_ASAP7_75T_SRAM%12 N_12_M5_s N_12_M4_d VSS PM_DHLX2_ASAP7_75T_SRAM%12
x_PM_DHLX2_ASAP7_75T_SRAM%13 N_13_M12_s N_13_M11_d VSS PM_DHLX2_ASAP7_75T_SRAM%13
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_20_n 2.66516e-19 $X=0.08 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 N_CLK_c_3_p N_4_c_21_n 2.48575e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.216
cc_4 N_CLK_c_3_p N_4_c_22_n 0.0020081f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.18
cc_5 CLK N_4_c_23_n 3.98992e-19 $X=0.08 $Y=0.119 $X2=0.018 $Y2=0.081
cc_6 CLK N_4_c_24_n 0.0020081f $X=0.08 $Y=0.119 $X2=0.018 $Y2=0.1305
cc_7 N_CLK_c_3_p N_4_c_25_n 3.00513e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.225
cc_8 CLK N_4_c_26_n 4.98319e-19 $X=0.08 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_3_p N_4_c_27_n 4.98319e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_10_p N_4_c_28_n 4.17e-19 $X=0.081 $Y=0.1305 $X2=0.152 $Y2=0.135
cc_11 N_CLK_c_11_p N_4_c_29_n 0.00111278f $X=0.081 $Y=0.135 $X2=0.152 $Y2=0.135
cc_12 N_CLK_c_3_p N_4_c_30_n 9.46659e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.1665
cc_13 N_CLK_c_3_p N_4_c_31_n 8.7692e-19 $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.189
cc_14 N_CLK_c_3_p N_4_c_32_n 0.00163094f $X=0.081 $Y=0.135 $X2=0.229 $Y2=0.189
cc_15 N_CLK_c_3_p N_4_c_33_n 9.73303e-19 $X=0.081 $Y=0.135 $X2=0.18 $Y2=0.189
cc_16 CLK N_6_c_120_n 6.45949e-19 $X=0.08 $Y=0.119 $X2=0.464 $Y2=0.179
cc_17 N_CLK_c_3_p N_6_c_121_n 6.45949e-19 $X=0.081 $Y=0.135 $X2=0.071 $Y2=0.216
cc_18 CLK N_6_c_122_n 7.98675e-19 $X=0.08 $Y=0.119 $X2=0 $Y2=0
cc_19 N_4_c_34_p N_D_M2_g 0.00341068f $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.054
cc_20 N_4_c_34_p N_D_c_103_n 9.3313e-19 $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.135
cc_21 N_4_c_36_p D 0.00227186f $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.119
cc_22 N_4_c_37_p D 0.00227186f $X=0.351 $Y=0.189 $X2=0.081 $Y2=0.119
cc_23 N_4_c_38_p D 2.29805e-19 $X=0.29 $Y=0.189 $X2=0.081 $Y2=0.119
cc_24 N_4_c_39_p D 6.20826e-19 $X=0.414 $Y=0.189 $X2=0.081 $Y2=0.119
cc_25 N_4_c_34_p N_6_M3_g 0.00355599f $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.054
cc_26 N_4_M4_g N_6_M3_g 0.00355599f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_27 N_4_c_34_p N_6_c_125_n 9.75871e-19 $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.135
cc_28 N_4_c_33_n N_6_c_126_n 0.00154329f $X=0.18 $Y=0.189 $X2=0.081 $Y2=0.1305
cc_29 N_4_c_28_n N_6_c_120_n 9.9131e-19 $X=0.152 $Y=0.135 $X2=0 $Y2=0
cc_30 N_4_c_38_p N_6_c_128_n 4.24027e-19 $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_31 N_4_c_32_n N_6_c_121_n 6.5319e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_32 N_4_c_33_n N_6_c_121_n 0.00305813f $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_33 N_4_c_32_n N_6_c_131_n 4.24027e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_34 N_4_c_49_p N_6_c_132_n 0.00351161f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_35 N_4_c_38_p N_6_c_132_n 0.00102041f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_36 N_4_c_51_p N_6_c_134_n 3.48096e-19 $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_37 N_4_c_36_p N_6_c_134_n 8.9767e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_38 N_4_c_37_p N_6_c_134_n 3.61885e-19 $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_39 N_4_c_38_p N_6_c_134_n 0.0160071f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_40 N_4_c_36_p N_6_c_138_n 0.00286743f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_41 N_4_c_39_p N_6_c_138_n 2.98086e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_42 N_4_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_43 N_4_c_58_p N_7_M5_g 0.00199227f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_44 N_4_c_59_p N_7_M5_g 5.16754e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_45 N_4_c_58_p N_7_c_159_n 4.44235e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.135
cc_46 N_4_c_58_p N_7_c_160_n 5.31675e-19 $X=0.513 $Y=0.18 $X2=0.08 $Y2=0.119
cc_47 N_4_c_58_p N_7_c_161_n 0.00169036f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.1305
cc_48 N_4_c_59_p N_7_c_162_n 7.15747e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_49 N_4_c_58_p N_7_c_163_n 0.00330898f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_50 N_4_c_58_p N_7_c_164_n 3.09575e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_51 N_4_c_58_p N_7_c_165_n 2.32568e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_52 N_4_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_53 N_4_c_58_p N_8_M6_g 0.00305656f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_54 N_4_c_36_p N_8_c_183_n 9.02348e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_55 N_4_c_37_p N_8_c_183_n 0.00144031f $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_56 N_4_c_37_p N_8_c_185_n 0.00138499f $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_57 N_4_c_39_p N_8_c_186_n 6.75805e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_58 N_4_c_73_p N_8_c_187_n 6.75805e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_59 N_4_c_73_p N_8_c_188_n 3.48842e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_60 N_4_c_73_p N_8_c_189_n 2.01793e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_61 N_4_M4_g N_8_c_190_n 2.73971e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_62 N_4_M4_g N_8_c_191_n 3.60498e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_63 N_4_M4_g N_8_c_192_n 2.06358e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_64 N_4_c_58_p N_8_c_193_n 4.82796e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_65 N_4_c_58_p N_8_c_194_n 7.81688e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_66 N_4_c_59_p N_8_c_195_n 0.001012f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_67 N_4_M4_g N_8_c_196_n 2.17193e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_68 N_4_c_83_p N_8_c_196_n 2.46239e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_69 N_4_c_83_p N_8_c_198_n 0.00694522f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_70 N_4_c_58_p N_8_c_198_n 0.00195859f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_71 N_4_c_59_p N_8_c_198_n 2.84813e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_72 N_4_c_87_p N_8_c_201_n 0.00127126f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_73 N_4_c_59_p N_8_c_201_n 0.00199566f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_74 N_4_c_87_p N_8_c_203_n 0.0011121f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_75 N_4_c_83_p N_8_c_203_n 3.67862e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_76 N_4_c_58_p N_8_c_203_n 4.28262e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_77 N_4_c_87_p N_8_c_206_n 7.05645e-19 $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_78 N_4_c_37_p N_8_c_206_n 2.96264e-19 $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_79 N_4_c_83_p N_8_c_206_n 3.05556e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_80 N_4_c_34_p N_10_c_264_n 0.00650944f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_81 N_4_c_36_p N_10_c_264_n 0.00135463f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_82 N_4_c_58_p N_11_M14_s 2.34172e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.216
cc_83 N_4_M4_g N_11_c_272_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_84 N_4_c_87_p N_11_c_272_n 0.0013957f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_85 N_4_c_73_p N_11_c_272_n 7.09553e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_86 N_4_c_58_p N_11_c_272_n 0.00230217f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_87 N_D_M2_g N_6_M3_g 2.82885e-19 $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_88 D N_6_c_141_n 0.00128741f $X=0.297 $Y=0.1165 $X2=0.459 $Y2=0.179
cc_89 N_D_c_110_p N_6_c_142_n 0.00128741f $X=0.297 $Y=0.135 $X2=0.056 $Y2=0.216
cc_90 D N_6_c_132_n 0.00138082f $X=0.297 $Y=0.1165 $X2=0.018 $Y2=0.18
cc_91 D N_6_c_134_n 0.0012236f $X=0.297 $Y=0.1165 $X2=0.018 $Y2=0.198
cc_92 D N_6_c_122_n 0.00128741f $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_93 D N_6_c_146_n 0.00128741f $X=0.297 $Y=0.1165 $X2=0.18 $Y2=0.135
cc_94 N_D_c_110_p N_6_c_147_n 0.00128741f $X=0.297 $Y=0.135 $X2=0.152 $Y2=0.135
cc_95 N_D_c_110_p N_8_c_183_n 3.23895e-19 $X=0.297 $Y=0.135 $X2=0.018 $Y2=0.18
cc_96 N_D_c_110_p N_8_c_185_n 3.35757e-19 $X=0.297 $Y=0.135 $X2=0.047 $Y2=0.036
cc_97 D N_8_c_188_n 2.05539e-19 $X=0.297 $Y=0.1165 $X2=0.054 $Y2=0.234
cc_98 D N_10_c_264_n 0.00445409f $X=0.297 $Y=0.1165 $X2=0.351 $Y2=0.134
cc_99 N_6_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_100 N_6_c_138_n N_8_c_183_n 4.65343e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_101 N_6_M3_g N_8_c_213_n 3.33314e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_102 N_6_c_138_n N_8_c_213_n 4.18821e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_103 N_6_c_138_n N_8_c_190_n 0.00307076f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_104 N_6_c_138_n N_8_c_196_n 2.60642e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_105 N_6_c_134_n N_8_c_198_n 8.94731e-19 $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_106 N_6_c_134_n N_10_c_264_n 8.35084e-19 $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_107 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_108 N_7_c_168_p N_8_M6_g 3.83894e-19 $X=0.581 $Y=0.036 $X2=0.135 $Y2=0.054
cc_109 N_7_c_169_p N_8_c_188_n 0.0017541f $X=0.522 $Y=0.036 $X2=0.054 $Y2=0.234
cc_110 N_7_c_170_p N_8_c_191_n 0.0017541f $X=0.513 $Y=0.082 $X2=0.152 $Y2=0.135
cc_111 N_7_c_171_p N_8_c_192_n 2.88106e-19 $X=0.621 $Y=0.121 $X2=0.152 $Y2=0.135
cc_112 N_7_c_168_p N_8_c_193_n 7.32482e-19 $X=0.581 $Y=0.036 $X2=0 $Y2=0
cc_113 N_7_c_173_p N_8_c_193_n 9.65274e-19 $X=0.621 $Y=0.139 $X2=0 $Y2=0
cc_114 N_7_M5_g N_8_c_195_n 4.16078e-19 $X=0.513 $Y=0.0405 $X2=0.189 $Y2=0.18
cc_115 N_7_c_170_p N_8_c_195_n 0.00115865f $X=0.513 $Y=0.082 $X2=0.189 $Y2=0.18
cc_116 N_7_c_160_n N_8_c_227_n 2.11538e-19 $X=0.592 $Y=0.0405 $X2=0.162
+ $Y2=0.189
cc_117 N_7_c_177_p N_8_c_227_n 8.8208e-19 $X=0.621 $Y=0.164 $X2=0.162 $Y2=0.189
cc_118 N_7_c_164_n N_8_c_227_n 5.92034e-19 $X=0.594 $Y=0.234 $X2=0.162 $Y2=0.189
cc_119 N_7_c_177_p N_8_c_230_n 3.90412e-19 $X=0.621 $Y=0.164 $X2=0.162 $Y2=0.189
cc_120 N_7_c_180_p N_8_c_231_n 0.00102407f $X=0.621 $Y=0.096 $X2=0.513 $Y2=0.189
cc_121 N_8_c_230_n N_Q_c_252_n 3.0124e-19 $X=0.783 $Y=0.153 $X2=0.351 $Y2=0.134
cc_122 N_8_c_230_n N_Q_c_253_n 3.84808e-19 $X=0.783 $Y=0.153 $X2=0.351
+ $Y2=0.2025
cc_123 N_8_M8_g N_Q_c_254_n 3.55084e-19 $X=0.783 $Y=0.0675 $X2=0.459 $Y2=0.179
cc_124 N_8_c_235_p N_Q_c_254_n 6.56888e-19 $X=0.783 $Y=0.136 $X2=0.459 $Y2=0.179
cc_125 N_8_c_230_n N_Q_c_256_n 2.54113e-19 $X=0.783 $Y=0.153 $X2=0.464 $Y2=0.179
cc_126 N_8_c_231_n N_Q_c_256_n 5.42522e-19 $X=0.729 $Y=0.136 $X2=0.464 $Y2=0.179
cc_127 N_8_c_235_p N_Q_c_256_n 5.42522e-19 $X=0.783 $Y=0.136 $X2=0.464 $Y2=0.179
cc_128 N_8_c_230_n N_Q_c_259_n 4.00565e-19 $X=0.783 $Y=0.153 $X2=0 $Y2=0
cc_129 N_8_M8_g N_Q_c_260_n 3.25912e-19 $X=0.783 $Y=0.0675 $X2=0.071 $Y2=0.054
cc_130 N_8_c_235_p N_Q_c_260_n 8.86582e-19 $X=0.783 $Y=0.136 $X2=0.071 $Y2=0.054
cc_131 N_8_c_230_n Q 2.27402e-19 $X=0.783 $Y=0.153 $X2=0 $Y2=0
cc_132 N_8_c_235_p N_Q_c_263_n 0.0028735f $X=0.783 $Y=0.136 $X2=0.056 $Y2=0.216
cc_133 N_8_c_183_n N_10_c_264_n 0.00119601f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.134
cc_134 N_8_c_188_n N_10_c_264_n 4.50844e-19 $X=0.45 $Y=0.036 $X2=0.351 $Y2=0.134
cc_135 N_8_c_189_n N_10_c_264_n 0.00394776f $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.134
cc_136 N_8_c_183_n N_11_c_272_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.134
cc_137 N_8_c_248_p N_11_c_272_n 0.00222776f $X=0.45 $Y=0.234 $X2=0.351 $Y2=0.134
cc_138 N_8_c_187_n N_11_c_272_n 0.00118584f $X=0.432 $Y=0.234 $X2=0.351
+ $Y2=0.134
cc_139 N_8_c_189_n N_11_c_272_n 5.72355e-19 $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.134
cc_140 N_8_c_251_p N_11_c_272_n 0.00116187f $X=0.459 $Y=0.225 $X2=0.351
+ $Y2=0.134

* END of "./DHLx2_ASAP7_75t_SRAM.pex.sp.DHLX2_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DHLx3_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:27:53 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DHLx3_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DHLx3_ASAP7_75t_SRAM.pex.sp.pex"
* File: DHLx3_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:27:53 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DHLX3_ASAP7_75T_SRAM%CLK 2 5 7 12 14 17 VSS
c18 17 VSS 5.41721e-21 $X=0.081 $Y=0.1305
c19 14 VSS 0.00699913f $X=0.081 $Y=0.135
c20 12 VSS 0.00699194f $X=0.08 $Y=0.119
c21 5 VSS 0.00183412f $X=0.081 $Y=0.135
c22 2 VSS 0.062963f $X=0.081 $Y=0.054
r23 16 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r24 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r25 12 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.126
r26 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DHLX3_ASAP7_75T_SRAM%4 2 7 10 13 16 24 26 29 31 34 37 38 39 41 44 51 56
+ 58 59 65 66 69 76 83 84 85 87 89 90 108 109 123 VSS
c85 123 VSS 5.19505e-19 $X=0.18 $Y=0.189
c86 122 VSS 1.53285e-19 $X=0.189 $Y=0.189
c87 118 VSS 7.0154e-20 $X=0.03 $Y=0.189
c88 117 VSS 5.9624e-19 $X=0.027 $Y=0.189
c89 109 VSS 7.76097e-19 $X=0.513 $Y=0.18
c90 108 VSS 0.05629f $X=0.513 $Y=0.18
c91 90 VSS 0.00123576f $X=0.45 $Y=0.189
c92 89 VSS 0.0038091f $X=0.414 $Y=0.189
c93 87 VSS 0.00305138f $X=0.513 $Y=0.189
c94 85 VSS 0.00251877f $X=0.29 $Y=0.189
c95 84 VSS 0.00700382f $X=0.229 $Y=0.189
c96 83 VSS 0.00149088f $X=0.351 $Y=0.189
c97 76 VSS 6.98042e-19 $X=0.033 $Y=0.189
c98 73 VSS 1.35996e-19 $X=0.351 $Y=0.18
c99 69 VSS 7.2814e-19 $X=0.351 $Y=0.134
c100 66 VSS 2.89511e-19 $X=0.189 $Y=0.1665
c101 65 VSS 3.97151e-19 $X=0.189 $Y=0.153
c102 64 VSS 1.55454e-19 $X=0.189 $Y=0.18
c103 59 VSS 0.00360014f $X=0.152 $Y=0.135
c104 58 VSS 4.22838e-19 $X=0.152 $Y=0.135
c105 56 VSS 0.00120122f $X=0.18 $Y=0.135
c106 54 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c107 53 VSS 0.00169428f $X=0.047 $Y=0.234
c108 51 VSS 0.00250477f $X=0.054 $Y=0.234
c109 49 VSS 0.00306385f $X=0.027 $Y=0.234
c110 47 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c111 46 VSS 0.00205521f $X=0.047 $Y=0.036
c112 44 VSS 0.00250477f $X=0.054 $Y=0.036
c113 42 VSS 0.00305101f $X=0.027 $Y=0.036
c114 41 VSS 0.00106422f $X=0.018 $Y=0.225
c115 39 VSS 0.00252163f $X=0.018 $Y=0.1305
c116 38 VSS 0.00142827f $X=0.018 $Y=0.081
c117 37 VSS 0.00214048f $X=0.018 $Y=0.18
c118 34 VSS 0.00507986f $X=0.056 $Y=0.216
c119 31 VSS 2.98509e-19 $X=0.071 $Y=0.216
c120 29 VSS 0.00454717f $X=0.056 $Y=0.054
c121 26 VSS 2.98509e-19 $X=0.071 $Y=0.054
c122 24 VSS 0.00218115f $X=0.464 $Y=0.179
c123 16 VSS 0.059523f $X=0.459 $Y=0.0405
c124 10 VSS 0.0605486f $X=0.351 $Y=0.134
c125 2 VSS 0.0627154f $X=0.135 $Y=0.054
r126 123 124 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.189 $X2=0.1845 $Y2=0.189
r127 122 124 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.189 $X2=0.1845 $Y2=0.189
r128 117 118 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.03 $Y2=0.189
r129 114 117 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.027 $Y2=0.189
r130 108 109 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18
+ $X2=0.513 $Y2=0.18
r131 89 90 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.414
+ $Y=0.189 $X2=0.45 $Y2=0.189
r132 87 90 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.45 $Y2=0.189
r133 87 109 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r134 84 85 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.189 $X2=0.29 $Y2=0.189
r135 82 89 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.414 $Y2=0.189
r136 82 85 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.29 $Y2=0.189
r137 82 83 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.189 $X2=0.351
+ $Y2=0.189
r138 80 123 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.189 $X2=0.18 $Y2=0.189
r139 79 84 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M2 $thickness=3.6e-08 $X=0.162
+ $Y=0.189 $X2=0.229 $Y2=0.189
r140 79 80 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.162 $Y=0.189 $X2=0.162
+ $Y2=0.189
r141 76 118 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.03 $Y2=0.189
r142 75 79 8.75926 $w=1.8e-08 $l=1.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.189 $X2=0.162 $Y2=0.189
r143 75 76 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.189 $X2=0.033
+ $Y2=0.189
r144 73 83 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.18 $X2=0.351 $Y2=0.189
r145 72 73 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.171 $X2=0.351 $Y2=0.18
r146 69 72 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.134 $X2=0.351 $Y2=0.171
r147 65 66 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.189 $Y2=0.1665
r148 64 122 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.189
r149 64 66 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.18 $X2=0.189 $Y2=0.1665
r150 63 65 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.153
r151 58 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.152 $Y=0.135 $X2=0.152
+ $Y2=0.135
r152 56 63 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r153 56 58 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.152 $Y2=0.135
r154 53 54 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r155 51 54 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r156 49 53 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r157 46 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r158 44 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r159 42 46 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r160 41 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r161 40 114 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.189
r162 40 41 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.198 $X2=0.018 $Y2=0.225
r163 38 39 3.36111 $w=1.8e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.1305
r164 37 114 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.189
r165 37 39 3.36111 $w=1.8e-08 $l=4.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.18 $X2=0.018 $Y2=0.1305
r166 36 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r167 36 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r168 34 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r169 31 34 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r170 29 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r171 26 29 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r172 24 108 42.2917 $w=2.4e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.464 $Y=0.179 $X2=0.513 $Y2=0.179
r173 19 24 3.57143 $w=2.8e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.179 $X2=0.464 $Y2=0.179
r174 16 19 518.891 $w=2e-08 $l=1.385e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.179
r175 10 69 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.134 $X2=0.351
+ $Y2=0.134
r176 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.134 $X2=0.351 $Y2=0.2025
r177 5 59 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.152 $Y2=0.135
r178 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r179 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DHLX3_ASAP7_75T_SRAM%D 2 5 7 11 15 VSS
c18 15 VSS 0.00225715f $X=0.297 $Y=0.135
c19 11 VSS 0.00893359f $X=0.297 $Y=0.1165
c20 5 VSS 0.00197947f $X=0.297 $Y=0.135
c21 2 VSS 0.0613821f $X=0.297 $Y=0.0675
r22 11 15 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1165 $X2=0.297 $Y2=0.135
r23 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r24 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r25 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DHLX3_ASAP7_75T_SRAM%6 2 5 7 9 14 17 19 24 26 31 32 34 37 40 45 55 56 58
+ VSS
c36 58 VSS 8.1019e-19 $X=0.243 $Y=0.2115
c37 56 VSS 4.07532e-19 $X=0.243 $Y=0.126
c38 55 VSS 0.00265408f $X=0.243 $Y=0.117
c39 45 VSS 0.00102533f $X=0.405 $Y=0.134
c40 40 VSS 0.00607715f $X=0.405 $Y=0.153
c41 37 VSS 0.00176992f $X=0.243 $Y=0.153
c42 34 VSS 5.5218e-19 $X=0.243 $Y=0.225
c43 32 VSS 0.00181981f $X=0.216 $Y=0.234
c44 31 VSS 0.0052254f $X=0.198 $Y=0.234
c45 26 VSS 0.00501032f $X=0.234 $Y=0.234
c46 25 VSS 0.00200074f $X=0.216 $Y=0.036
c47 24 VSS 0.00549661f $X=0.198 $Y=0.036
c48 19 VSS 0.00500597f $X=0.234 $Y=0.036
c49 17 VSS 0.00666939f $X=0.16 $Y=0.216
c50 12 VSS 0.00625354f $X=0.16 $Y=0.054
c51 5 VSS 0.0015003f $X=0.405 $Y=0.134
c52 2 VSS 0.059003f $X=0.405 $Y=0.0675
r53 57 58 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.198 $X2=0.243 $Y2=0.2115
r54 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.117 $X2=0.243 $Y2=0.126
r55 41 45 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.405 $Y2=0.134
r56 40 41 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r57 37 57 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.198
r58 37 56 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.126
r59 36 40 11 $w=1.8e-08 $l=1.62e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.405 $Y2=0.153
r60 36 37 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.153 $X2=0.243
+ $Y2=0.153
r61 34 58 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.2115
r62 33 55 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.117
r63 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.216 $Y2=0.234
r64 28 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.198 $Y2=0.234
r65 26 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r66 26 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r67 24 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.216 $Y2=0.036
r68 21 24 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r69 19 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r70 19 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r71 17 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r72 14 17 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r73 12 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r74 9 12 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r75 5 45 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.134 $X2=0.405
+ $Y2=0.134
r76 5 7 357.791 $w=2e-08 $l=9.55e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.134 $X2=0.405 $Y2=0.2295
r77 2 5 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.134
.ends

.subckt PM_DHLX3_ASAP7_75T_SRAM%7 2 5 7 9 12 14 17 21 24 25 29 33 34 35 36 37 38 39
+ 42 47 48 VSS
c32 48 VSS 0.00241451f $X=0.612 $Y=0.234
c33 47 VSS 0.00208935f $X=0.621 $Y=0.234
c34 42 VSS 0.00170515f $X=0.594 $Y=0.234
c35 40 VSS 3.06787e-19 $X=0.621 $Y=0.216
c36 39 VSS 3.9255e-19 $X=0.621 $Y=0.207
c37 38 VSS 4.86711e-20 $X=0.621 $Y=0.167
c38 37 VSS 7.79237e-19 $X=0.621 $Y=0.164
c39 36 VSS 4.90317e-19 $X=0.621 $Y=0.139
c40 35 VSS 9.27636e-19 $X=0.621 $Y=0.121
c41 34 VSS 1.31821e-19 $X=0.621 $Y=0.096
c42 33 VSS 5.42108e-19 $X=0.621 $Y=0.09
c43 32 VSS 4.22112e-19 $X=0.621 $Y=0.225
c44 30 VSS 7.17067e-19 $X=0.5875 $Y=0.036
c45 29 VSS 0.00656714f $X=0.581 $Y=0.036
c46 25 VSS 0.00222389f $X=0.522 $Y=0.036
c47 24 VSS 0.00460947f $X=0.612 $Y=0.036
c48 21 VSS 5.75409e-19 $X=0.513 $Y=0.082
c49 17 VSS 0.00441196f $X=0.592 $Y=0.2295
c50 12 VSS 0.00458554f $X=0.592 $Y=0.0405
c51 5 VSS 0.00257008f $X=0.513 $Y=0.082
c52 2 VSS 0.058175f $X=0.513 $Y=0.0405
r53 48 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r54 47 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r55 42 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.612 $Y2=0.234
r56 39 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.207 $X2=0.621 $Y2=0.216
r57 38 39 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.207
r58 37 38 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.164 $X2=0.621 $Y2=0.167
r59 36 37 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.139 $X2=0.621 $Y2=0.164
r60 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.121 $X2=0.621 $Y2=0.139
r61 34 35 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.096 $X2=0.621 $Y2=0.121
r62 33 34 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.621 $Y2=0.096
r63 32 47 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.234
r64 32 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.216
r65 31 33 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.09
r66 29 30 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.581
+ $Y=0.036 $X2=0.5875 $Y2=0.036
r67 27 30 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.5875 $Y2=0.036
r68 25 29 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.581 $Y2=0.036
r69 24 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r70 24 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.594 $Y2=0.036
r71 19 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.513 $Y=0.045 $X2=0.522 $Y2=0.036
r72 19 21 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.082
r73 17 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r74 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r75 12 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036 $X2=0.594
+ $Y2=0.036
r76 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.592 $Y2=0.0405
r77 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.082 $X2=0.513
+ $Y2=0.082
r78 5 7 552.609 $w=2e-08 $l=1.475e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.082 $X2=0.513 $Y2=0.2295
r79 2 5 155.48 $w=2e-08 $l=4.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.082
.ends

.subckt PM_DHLX3_ASAP7_75T_SRAM%8 2 7 10 15 18 23 26 31 33 38 41 45 46 49 54 55 56
+ 57 58 61 64 65 66 69 71 72 77 80 85 86 91 99 104 109 121 122 123 VSS
c86 123 VSS 3.47616e-19 $X=0.459 $Y=0.207
c87 122 VSS 3.33252e-19 $X=0.459 $Y=0.189
c88 121 VSS 1.82803e-20 $X=0.459 $Y=0.171
c89 109 VSS 0.00125596f $X=0.837 $Y=0.136
c90 104 VSS 0.00102119f $X=0.783 $Y=0.136
c91 99 VSS 0.00127432f $X=0.729 $Y=0.136
c92 91 VSS 0.00987939f $X=0.837 $Y=0.153
c93 86 VSS 0.0040364f $X=0.628 $Y=0.153
c94 85 VSS 0.00146565f $X=0.527 $Y=0.153
c95 80 VSS 4.02226e-19 $X=0.459 $Y=0.153
c96 77 VSS 5.11551e-19 $X=0.459 $Y=0.225
c97 76 VSS 2.42691e-19 $X=0.459 $Y=0.13
c98 72 VSS 3.63326e-20 $X=0.522 $Y=0.13
c99 71 VSS 0.00173658f $X=0.504 $Y=0.13
c100 69 VSS 0.00150363f $X=0.567 $Y=0.13
c101 66 VSS 2.19687e-19 $X=0.459 $Y=0.106
c102 65 VSS 3.06086e-19 $X=0.459 $Y=0.096
c103 64 VSS 1.63148e-19 $X=0.459 $Y=0.121
c104 61 VSS 0.00271748f $X=0.432 $Y=0.036
c105 58 VSS 0.00636114f $X=0.45 $Y=0.036
c106 57 VSS 0.00163742f $X=0.432 $Y=0.234
c107 56 VSS 0.00142296f $X=0.414 $Y=0.234
c108 55 VSS 0.00166696f $X=0.396 $Y=0.234
c109 54 VSS 0.00188233f $X=0.379 $Y=0.234
c110 49 VSS 0.00408073f $X=0.45 $Y=0.234
c111 48 VSS 5.7602e-19 $X=0.378 $Y=0.2295
c112 45 VSS 0.00367263f $X=0.378 $Y=0.2025
c113 42 VSS 3.44634e-20 $X=0.3735 $Y=0.216
c114 40 VSS 5.36734e-19 $X=0.432 $Y=0.0405
c115 29 VSS 0.00216451f $X=0.837 $Y=0.136
c116 26 VSS 0.06069f $X=0.837 $Y=0.0675
c117 21 VSS 0.00190168f $X=0.783 $Y=0.136
c118 18 VSS 0.0608917f $X=0.783 $Y=0.0675
c119 13 VSS 0.00281985f $X=0.729 $Y=0.136
c120 10 VSS 0.0638816f $X=0.729 $Y=0.0675
c121 5 VSS 0.00267415f $X=0.567 $Y=0.13
c122 2 VSS 0.0627953f $X=0.567 $Y=0.0405
r123 122 123 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.189 $X2=0.459 $Y2=0.207
r124 121 122 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.171 $X2=0.459 $Y2=0.189
r125 120 121 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.164 $X2=0.459 $Y2=0.171
r126 91 109 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.837 $Y=0.153 $X2=0.837
+ $Y2=0.153
r127 88 91 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.783
+ $Y=0.153 $X2=0.837 $Y2=0.153
r128 88 104 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.783 $Y=0.153 $X2=0.783
+ $Y2=0.153
r129 85 86 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.628 $Y2=0.153
r130 83 88 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.783 $Y2=0.153
r131 83 86 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M2 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.628 $Y2=0.153
r132 83 99 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.729 $Y=0.153 $X2=0.729
+ $Y2=0.153
r133 80 120 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.459 $Y2=0.164
r134 79 85 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.527 $Y2=0.153
r135 79 80 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.459 $Y=0.153 $X2=0.459
+ $Y2=0.153
r136 77 123 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.207
r137 75 80 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.139 $X2=0.459 $Y2=0.153
r138 75 76 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.139 $X2=0.459 $Y2=0.13
r139 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.13 $X2=0.522 $Y2=0.13
r140 69 72 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.13 $X2=0.522 $Y2=0.13
r141 67 76 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.13 $X2=0.459 $Y2=0.13
r142 67 71 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.13 $X2=0.504 $Y2=0.13
r143 65 66 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.096 $X2=0.459 $Y2=0.106
r144 64 76 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.121 $X2=0.459 $Y2=0.13
r145 64 66 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.121 $X2=0.459 $Y2=0.106
r146 63 65 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.096
r147 60 61 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r148 58 63 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r149 58 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.432 $Y2=0.036
r150 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.432 $Y2=0.234
r151 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r152 54 55 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.379
+ $Y=0.234 $X2=0.396 $Y2=0.234
r153 51 54 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.379 $Y2=0.234
r154 49 77 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r155 49 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.432 $Y2=0.234
r156 46 48 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r157 45 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r158 42 48 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r159 42 45 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r160 41 45 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r161 38 40 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r162 37 61 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r163 34 40 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r164 34 37 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r165 33 37 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r166 29 109 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.837 $Y=0.136
+ $X2=0.837 $Y2=0.136
r167 29 31 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.136 $X2=0.837 $Y2=0.2025
r168 26 29 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0675 $X2=0.837 $Y2=0.136
r169 21 104 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.136
+ $X2=0.783 $Y2=0.136
r170 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.136 $X2=0.783 $Y2=0.2025
r171 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.136
r172 13 99 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.729 $Y=0.136 $X2=0.729
+ $Y2=0.136
r173 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.136 $X2=0.729 $Y2=0.2025
r174 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.136
r175 5 69 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.13 $X2=0.567
+ $Y2=0.13
r176 5 7 372.777 $w=2e-08 $l=9.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.13 $X2=0.567 $Y2=0.2295
r177 2 5 335.312 $w=2e-08 $l=8.95e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.13
.ends

.subckt PM_DHLX3_ASAP7_75T_SRAM%Q 1 6 7 11 14 16 17 20 24 28 29 30 31 32 33 34 43
+ 44 45 46 47 48 52 54 VSS
c34 56 VSS 0.00207706f $X=0.891 $Y=0.196
c35 54 VSS 0.00149295f $X=0.891 $Y=0.1215
c36 53 VSS 0.00272046f $X=0.891 $Y=0.09
c37 52 VSS 0.00221453f $X=0.893 $Y=0.153
c38 50 VSS 0.00156747f $X=0.891 $Y=0.225
c39 48 VSS 0.00146362f $X=0.846 $Y=0.234
c40 47 VSS 0.00311681f $X=0.828 $Y=0.234
c41 46 VSS 0.00146362f $X=0.792 $Y=0.234
c42 45 VSS 0.00596994f $X=0.774 $Y=0.234
c43 44 VSS 0.00146362f $X=0.738 $Y=0.234
c44 43 VSS 0.00361142f $X=0.72 $Y=0.234
c45 35 VSS 0.00935225f $X=0.882 $Y=0.234
c46 34 VSS 0.00146362f $X=0.846 $Y=0.036
c47 33 VSS 0.00311891f $X=0.828 $Y=0.036
c48 32 VSS 0.00146362f $X=0.792 $Y=0.036
c49 31 VSS 0.00597353f $X=0.774 $Y=0.036
c50 30 VSS 0.00146362f $X=0.738 $Y=0.036
c51 29 VSS 0.00361553f $X=0.72 $Y=0.036
c52 28 VSS 0.0097069f $X=0.81 $Y=0.036
c53 24 VSS 0.00585995f $X=0.702 $Y=0.036
c54 21 VSS 0.00933023f $X=0.882 $Y=0.036
c55 20 VSS 0.00935224f $X=0.81 $Y=0.2025
c56 16 VSS 6.15431e-19 $X=0.827 $Y=0.2025
c57 14 VSS 0.00596555f $X=0.704 $Y=0.2025
c58 11 VSS 3.4597e-19 $X=0.719 $Y=0.2025
c59 6 VSS 6.1381e-19 $X=0.827 $Y=0.0675
c60 1 VSS 3.44349e-19 $X=0.719 $Y=0.0675
r61 55 56 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.167 $X2=0.891 $Y2=0.196
r62 53 54 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.09 $X2=0.891 $Y2=0.1215
r63 52 55 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.891 $Y2=0.167
r64 52 54 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.153 $X2=0.891 $Y2=0.1215
r65 50 56 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.225 $X2=0.891 $Y2=0.196
r66 49 53 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.045 $X2=0.891 $Y2=0.09
r67 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.846 $Y2=0.234
r68 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.234 $X2=0.792 $Y2=0.234
r69 44 45 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.234 $X2=0.774 $Y2=0.234
r70 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.234 $X2=0.738 $Y2=0.234
r71 41 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.234 $X2=0.828 $Y2=0.234
r72 41 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.234 $X2=0.792 $Y2=0.234
r73 37 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.234 $X2=0.72 $Y2=0.234
r74 35 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.234 $X2=0.891 $Y2=0.225
r75 35 48 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.234 $X2=0.846 $Y2=0.234
r76 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.846 $Y2=0.036
r77 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.036 $X2=0.792 $Y2=0.036
r78 30 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.738
+ $Y=0.036 $X2=0.774 $Y2=0.036
r79 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.738 $Y2=0.036
r80 27 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.036 $X2=0.828 $Y2=0.036
r81 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.036 $X2=0.792 $Y2=0.036
r82 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.036 $X2=0.81
+ $Y2=0.036
r83 23 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.036 $X2=0.72 $Y2=0.036
r84 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.036 $X2=0.702
+ $Y2=0.036
r85 21 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.036 $X2=0.891 $Y2=0.045
r86 21 34 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.846 $Y2=0.036
r87 20 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.234 $X2=0.81
+ $Y2=0.234
r88 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2025 $X2=0.81 $Y2=0.2025
r89 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.2025 $X2=0.81 $Y2=0.2025
r90 14 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.234 $X2=0.702
+ $Y2=0.234
r91 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2025 $X2=0.704 $Y2=0.2025
r92 10 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.81
+ $Y=0.0675 $X2=0.81 $Y2=0.036
r93 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.0675 $X2=0.81 $Y2=0.0675
r94 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.0675 $X2=0.81 $Y2=0.0675
r95 4 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.702
+ $Y=0.0675 $X2=0.702 $Y2=0.036
r96 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0675 $X2=0.704 $Y2=0.0675
.ends

.subckt PM_DHLX3_ASAP7_75T_SRAM%10 1 6 9 VSS
c7 9 VSS 0.0266194f $X=0.38 $Y=0.0675
c8 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c9 4 VSS 3.9325e-19 $X=0.322 $Y=0.0675
r10 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r12 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DHLX3_ASAP7_75T_SRAM%11 1 6 9 VSS
c10 9 VSS 0.0211086f $X=0.488 $Y=0.2295
c11 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c12 4 VSS 2.84146e-19 $X=0.43 $Y=0.2295
r13 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r15 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DHLX3_ASAP7_75T_SRAM%12 1 2 VSS
c0 1 VSS 0.00220425f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DHLX3_ASAP7_75T_SRAM%13 1 2 VSS
c0 1 VSS 0.00221026f $X=0.341 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends


* END of "./DHLx3_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DHLx3_ASAP7_75t_SRAM  VSS VDD CLK D Q
* 
* Q	Q
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_10_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_6_M3_g N_10_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_12_M4_d N_4_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_12_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 VSS N_8_M7_g N_Q_M7_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M8 VSS N_8_M8_g N_Q_M8_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773 $Y=0.027
M9 VSS N_8_M9_g N_Q_M9_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827 $Y=0.027
M10 VDD N_CLK_M10_g N_4_M10_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M11 N_6_M11_d N_4_M11_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M12 N_13_M12_d N_D_M12_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M13 N_8_M13_d N_4_M13_g N_13_M13_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M14 N_11_M14_d N_6_M14_g N_8_M14_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M15 VDD N_7_M15_g N_11_M15_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M16 N_7_M16_d N_8_M16_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M17 VDD N_8_M17_g N_Q_M17_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M18 VDD N_8_M18_g N_Q_M18_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
M19 VDD N_8_M19_g N_Q_M19_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.162
*
* 
* .include "DHLx3_ASAP7_75t_SRAM.pex.sp.DHLX3_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DHLx3_ASAP7_75t_SRAM.pex.sp.DHLX3_ASAP7_75T_SRAM.pxi"
* File: DHLx3_ASAP7_75t_SRAM.pex.sp.DHLX3_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:27:53 2017
* 
x_PM_DHLX3_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_11_p N_CLK_M10_g CLK N_CLK_c_3_p
+ N_CLK_c_10_p VSS PM_DHLX3_ASAP7_75T_SRAM%CLK
x_PM_DHLX3_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M11_g N_4_c_34_p N_4_M13_g N_4_M4_g
+ N_4_c_88_p N_4_M0_s N_4_c_20_n N_4_M10_s N_4_c_21_n N_4_c_22_n N_4_c_23_n
+ N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_49_p N_4_c_28_n N_4_c_29_n
+ N_4_c_51_p N_4_c_30_n N_4_c_36_p N_4_c_31_n N_4_c_37_p N_4_c_32_n N_4_c_38_p
+ N_4_c_84_p N_4_c_39_p N_4_c_74_p N_4_c_58_p N_4_c_59_p N_4_c_33_n VSS
+ PM_DHLX3_ASAP7_75T_SRAM%4
x_PM_DHLX3_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_105_n N_D_M12_g D N_D_c_112_p VSS
+ PM_DHLX3_ASAP7_75T_SRAM%D
x_PM_DHLX3_ASAP7_75T_SRAM%6 N_6_M3_g N_6_c_127_n N_6_M14_g N_6_M1_d N_6_M11_d
+ N_6_c_128_n N_6_c_143_n N_6_c_122_n N_6_c_130_n N_6_c_123_n N_6_c_133_n
+ N_6_c_144_n N_6_c_134_n N_6_c_136_n N_6_c_140_n N_6_c_124_n N_6_c_148_n
+ N_6_c_149_n VSS PM_DHLX3_ASAP7_75T_SRAM%6
x_PM_DHLX3_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_161_n N_7_M15_g N_7_M6_d N_7_c_162_n
+ N_7_M16_d N_7_c_163_n N_7_c_173_p N_7_c_188_p N_7_c_172_p N_7_c_171_p
+ N_7_c_187_p N_7_c_183_p N_7_c_174_p N_7_c_176_p N_7_c_180_p N_7_c_164_n
+ N_7_c_166_n N_7_c_167_n N_7_c_189_p N_7_c_168_n VSS PM_DHLX3_ASAP7_75T_SRAM%7
x_PM_DHLX3_ASAP7_75T_SRAM%8 N_8_M6_g N_8_M16_g N_8_M7_g N_8_M17_g N_8_M8_g
+ N_8_M18_g N_8_M9_g N_8_M19_g N_8_M3_d N_8_M4_s N_8_M13_d N_8_c_192_n N_8_M14_s
+ N_8_c_272_p N_8_c_194_n N_8_c_195_n N_8_c_222_n N_8_c_196_n N_8_c_197_n
+ N_8_c_198_n N_8_c_199_n N_8_c_200_n N_8_c_201_n N_8_c_202_n N_8_c_203_n
+ N_8_c_204_n N_8_c_275_p N_8_c_205_n N_8_c_207_n N_8_c_236_n N_8_c_239_n
+ N_8_c_240_n N_8_c_246_p N_8_c_247_p N_8_c_210_n N_8_c_212_n N_8_c_215_n VSS
+ PM_DHLX3_ASAP7_75T_SRAM%8
x_PM_DHLX3_ASAP7_75T_SRAM%Q N_Q_M7_s N_Q_M9_s N_Q_M8_s N_Q_M17_s N_Q_c_276_n
+ N_Q_M19_s N_Q_M18_s N_Q_c_284_n N_Q_c_279_n N_Q_c_287_n N_Q_c_281_n
+ N_Q_c_291_n N_Q_c_293_n N_Q_c_294_n N_Q_c_296_n N_Q_c_297_n N_Q_c_282_n
+ N_Q_c_300_n N_Q_c_302_n N_Q_c_303_n N_Q_c_305_n N_Q_c_306_n Q N_Q_c_309_n VSS
+ PM_DHLX3_ASAP7_75T_SRAM%Q
x_PM_DHLX3_ASAP7_75T_SRAM%10 N_10_M2_d N_10_M3_s N_10_c_310_n VSS
+ PM_DHLX3_ASAP7_75T_SRAM%10
x_PM_DHLX3_ASAP7_75T_SRAM%11 N_11_M14_d N_11_M15_s N_11_c_318_n VSS
+ PM_DHLX3_ASAP7_75T_SRAM%11
x_PM_DHLX3_ASAP7_75T_SRAM%12 N_12_M5_s N_12_M4_d VSS PM_DHLX3_ASAP7_75T_SRAM%12
x_PM_DHLX3_ASAP7_75T_SRAM%13 N_13_M13_s N_13_M12_d VSS PM_DHLX3_ASAP7_75T_SRAM%13
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_20_n 2.66516e-19 $X=0.08 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 N_CLK_c_3_p N_4_c_21_n 2.48575e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.216
cc_4 N_CLK_c_3_p N_4_c_22_n 0.0020081f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.18
cc_5 CLK N_4_c_23_n 3.98992e-19 $X=0.08 $Y=0.119 $X2=0.018 $Y2=0.081
cc_6 CLK N_4_c_24_n 0.0020081f $X=0.08 $Y=0.119 $X2=0.018 $Y2=0.1305
cc_7 N_CLK_c_3_p N_4_c_25_n 3.00513e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.225
cc_8 CLK N_4_c_26_n 4.98319e-19 $X=0.08 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_3_p N_4_c_27_n 4.98319e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_10_p N_4_c_28_n 4.17e-19 $X=0.081 $Y=0.1305 $X2=0.152 $Y2=0.135
cc_11 N_CLK_c_11_p N_4_c_29_n 0.00111278f $X=0.081 $Y=0.135 $X2=0.152 $Y2=0.135
cc_12 N_CLK_c_3_p N_4_c_30_n 9.46659e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.1665
cc_13 N_CLK_c_3_p N_4_c_31_n 8.7692e-19 $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.189
cc_14 N_CLK_c_3_p N_4_c_32_n 0.00163094f $X=0.081 $Y=0.135 $X2=0.229 $Y2=0.189
cc_15 N_CLK_c_3_p N_4_c_33_n 9.73303e-19 $X=0.081 $Y=0.135 $X2=0.18 $Y2=0.189
cc_16 CLK N_6_c_122_n 6.45949e-19 $X=0.08 $Y=0.119 $X2=0.464 $Y2=0.179
cc_17 N_CLK_c_3_p N_6_c_123_n 6.45949e-19 $X=0.081 $Y=0.135 $X2=0.071 $Y2=0.216
cc_18 CLK N_6_c_124_n 7.98675e-19 $X=0.08 $Y=0.119 $X2=0 $Y2=0
cc_19 N_4_c_34_p N_D_M2_g 0.00341068f $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.054
cc_20 N_4_c_34_p N_D_c_105_n 9.3313e-19 $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.135
cc_21 N_4_c_36_p D 0.00227186f $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.119
cc_22 N_4_c_37_p D 0.00227186f $X=0.351 $Y=0.189 $X2=0.081 $Y2=0.119
cc_23 N_4_c_38_p D 2.29805e-19 $X=0.29 $Y=0.189 $X2=0.081 $Y2=0.119
cc_24 N_4_c_39_p D 6.20826e-19 $X=0.414 $Y=0.189 $X2=0.081 $Y2=0.119
cc_25 N_4_c_34_p N_6_M3_g 0.00355599f $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.054
cc_26 N_4_M4_g N_6_M3_g 0.00355599f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_27 N_4_c_34_p N_6_c_127_n 9.75871e-19 $X=0.351 $Y=0.134 $X2=0.081 $Y2=0.135
cc_28 N_4_c_33_n N_6_c_128_n 0.00154329f $X=0.18 $Y=0.189 $X2=0.081 $Y2=0.1305
cc_29 N_4_c_28_n N_6_c_122_n 9.9131e-19 $X=0.152 $Y=0.135 $X2=0 $Y2=0
cc_30 N_4_c_38_p N_6_c_130_n 4.24027e-19 $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_31 N_4_c_32_n N_6_c_123_n 6.5319e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_32 N_4_c_33_n N_6_c_123_n 0.00305813f $X=0.18 $Y=0.189 $X2=0 $Y2=0
cc_33 N_4_c_32_n N_6_c_133_n 4.24027e-19 $X=0.229 $Y=0.189 $X2=0 $Y2=0
cc_34 N_4_c_49_p N_6_c_134_n 0.00351161f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_35 N_4_c_38_p N_6_c_134_n 0.00102041f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_36 N_4_c_51_p N_6_c_136_n 3.48096e-19 $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_37 N_4_c_36_p N_6_c_136_n 8.9767e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_38 N_4_c_37_p N_6_c_136_n 3.61885e-19 $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_39 N_4_c_38_p N_6_c_136_n 0.0160071f $X=0.29 $Y=0.189 $X2=0 $Y2=0
cc_40 N_4_c_36_p N_6_c_140_n 0.00286743f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_41 N_4_c_39_p N_6_c_140_n 2.98086e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_42 N_4_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_43 N_4_c_58_p N_7_M5_g 0.00199227f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_44 N_4_c_59_p N_7_M5_g 5.16754e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_45 N_4_c_58_p N_7_c_161_n 4.44235e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.135
cc_46 N_4_c_58_p N_7_c_162_n 5.31675e-19 $X=0.513 $Y=0.18 $X2=0.08 $Y2=0.119
cc_47 N_4_c_58_p N_7_c_163_n 0.00169036f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.1305
cc_48 N_4_c_58_p N_7_c_164_n 6.34096e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_49 N_4_c_59_p N_7_c_164_n 7.16706e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_50 N_4_c_58_p N_7_c_166_n 0.00238219f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_51 N_4_c_58_p N_7_c_167_n 3.09575e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_52 N_4_c_58_p N_7_c_168_n 2.32568e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_53 N_4_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_54 N_4_c_58_p N_8_M6_g 0.00305656f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_55 N_4_c_36_p N_8_c_192_n 9.02348e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_56 N_4_c_37_p N_8_c_192_n 0.00144031f $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_57 N_4_c_37_p N_8_c_194_n 0.00138499f $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_58 N_4_c_39_p N_8_c_195_n 6.75805e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_59 N_4_c_74_p N_8_c_196_n 6.75805e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_60 N_4_c_74_p N_8_c_197_n 3.48842e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_61 N_4_c_74_p N_8_c_198_n 2.01793e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_62 N_4_M4_g N_8_c_199_n 2.73971e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_63 N_4_M4_g N_8_c_200_n 3.60498e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_64 N_4_M4_g N_8_c_201_n 2.06358e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_65 N_4_c_58_p N_8_c_202_n 4.82796e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_66 N_4_c_58_p N_8_c_203_n 7.81688e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_67 N_4_c_59_p N_8_c_204_n 0.001012f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_68 N_4_M4_g N_8_c_205_n 2.17193e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_69 N_4_c_84_p N_8_c_205_n 2.46239e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_70 N_4_c_84_p N_8_c_207_n 0.00694522f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_71 N_4_c_58_p N_8_c_207_n 0.00195859f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_72 N_4_c_59_p N_8_c_207_n 2.84813e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_73 N_4_c_88_p N_8_c_210_n 0.00127126f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_74 N_4_c_59_p N_8_c_210_n 0.00199566f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_75 N_4_c_88_p N_8_c_212_n 0.0011121f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_76 N_4_c_84_p N_8_c_212_n 3.67862e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_77 N_4_c_58_p N_8_c_212_n 4.28262e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_78 N_4_c_88_p N_8_c_215_n 7.05645e-19 $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_79 N_4_c_37_p N_8_c_215_n 2.96264e-19 $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_80 N_4_c_84_p N_8_c_215_n 3.05556e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_81 N_4_c_58_p N_Q_c_276_n 0.00114499f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.135
cc_82 N_4_c_34_p N_10_c_310_n 0.00650944f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_83 N_4_c_36_p N_10_c_310_n 0.00135463f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_84 N_4_c_58_p N_11_M15_s 2.34172e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.216
cc_85 N_4_M4_g N_11_c_318_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_86 N_4_c_88_p N_11_c_318_n 0.0013957f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_87 N_4_c_74_p N_11_c_318_n 7.09553e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_88 N_4_c_58_p N_11_c_318_n 0.00230217f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_89 N_D_M2_g N_6_M3_g 2.82885e-19 $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_90 D N_6_c_143_n 0.00128741f $X=0.297 $Y=0.1165 $X2=0.459 $Y2=0.179
cc_91 N_D_c_112_p N_6_c_144_n 0.00128741f $X=0.297 $Y=0.135 $X2=0.056 $Y2=0.216
cc_92 D N_6_c_134_n 0.00138082f $X=0.297 $Y=0.1165 $X2=0.018 $Y2=0.18
cc_93 D N_6_c_136_n 0.0012236f $X=0.297 $Y=0.1165 $X2=0.018 $Y2=0.198
cc_94 D N_6_c_124_n 0.00128741f $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_95 D N_6_c_148_n 0.00128741f $X=0.297 $Y=0.1165 $X2=0.18 $Y2=0.135
cc_96 N_D_c_112_p N_6_c_149_n 0.00128741f $X=0.297 $Y=0.135 $X2=0.152 $Y2=0.135
cc_97 N_D_c_112_p N_8_c_192_n 3.23895e-19 $X=0.297 $Y=0.135 $X2=0.054 $Y2=0.036
cc_98 N_D_c_112_p N_8_c_194_n 3.35757e-19 $X=0.297 $Y=0.135 $X2=0.0505 $Y2=0.234
cc_99 D N_8_c_197_n 2.05539e-19 $X=0.297 $Y=0.1165 $X2=0.152 $Y2=0.135
cc_100 D N_10_c_310_n 0.00445409f $X=0.297 $Y=0.1165 $X2=0.351 $Y2=0.134
cc_101 N_6_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_102 N_6_c_140_n N_8_c_192_n 4.65343e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_103 N_6_M3_g N_8_c_222_n 3.33314e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_104 N_6_c_140_n N_8_c_222_n 4.18821e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_105 N_6_c_140_n N_8_c_199_n 0.00307076f $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_106 N_6_c_140_n N_8_c_205_n 2.60642e-19 $X=0.405 $Y=0.134 $X2=0 $Y2=0
cc_107 N_6_c_136_n N_8_c_207_n 9.00219e-19 $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_108 N_6_c_136_n N_10_c_310_n 8.35084e-19 $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_109 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_110 N_7_c_171_p N_8_M6_g 3.83894e-19 $X=0.581 $Y=0.036 $X2=0.135 $Y2=0.054
cc_111 N_7_c_172_p N_8_c_197_n 0.0017541f $X=0.522 $Y=0.036 $X2=0.152 $Y2=0.135
cc_112 N_7_c_173_p N_8_c_200_n 0.0017541f $X=0.513 $Y=0.082 $X2=0.189 $Y2=0.153
cc_113 N_7_c_174_p N_8_c_201_n 2.86032e-19 $X=0.621 $Y=0.121 $X2=0.189
+ $Y2=0.1665
cc_114 N_7_c_171_p N_8_c_202_n 7.32482e-19 $X=0.581 $Y=0.036 $X2=0.351 $Y2=0.134
cc_115 N_7_c_176_p N_8_c_202_n 9.78244e-19 $X=0.621 $Y=0.139 $X2=0.351 $Y2=0.134
cc_116 N_7_M5_g N_8_c_204_n 4.16078e-19 $X=0.513 $Y=0.0405 $X2=0.351 $Y2=0.171
cc_117 N_7_c_173_p N_8_c_204_n 0.00115865f $X=0.513 $Y=0.082 $X2=0.351 $Y2=0.171
cc_118 N_7_c_162_n N_8_c_236_n 2.11538e-19 $X=0.592 $Y=0.0405 $X2=0.513
+ $Y2=0.189
cc_119 N_7_c_180_p N_8_c_236_n 8.8208e-19 $X=0.621 $Y=0.164 $X2=0.513 $Y2=0.189
cc_120 N_7_c_167_n N_8_c_236_n 5.92034e-19 $X=0.594 $Y=0.234 $X2=0.513 $Y2=0.189
cc_121 N_7_c_180_p N_8_c_239_n 3.90412e-19 $X=0.621 $Y=0.164 $X2=0 $Y2=0
cc_122 N_7_c_183_p N_8_c_240_n 0.00102774f $X=0.621 $Y=0.096 $X2=0 $Y2=0
cc_123 N_7_c_163_n N_Q_c_276_n 4.7734e-19 $X=0.592 $Y=0.2295 $X2=0 $Y2=0
cc_124 N_7_c_166_n N_Q_c_276_n 8.1674e-19 $X=0.621 $Y=0.207 $X2=0 $Y2=0
cc_125 N_7_c_162_n N_Q_c_279_n 4.7734e-19 $X=0.592 $Y=0.0405 $X2=0.464 $Y2=0.179
cc_126 N_7_c_187_p N_Q_c_279_n 0.00145282f $X=0.621 $Y=0.09 $X2=0.464 $Y2=0.179
cc_127 N_7_c_188_p N_Q_c_281_n 8.40653e-19 $X=0.612 $Y=0.036 $X2=0.056 $Y2=0.054
cc_128 N_7_c_189_p N_Q_c_282_n 7.85494e-19 $X=0.621 $Y=0.234 $X2=0.054 $Y2=0.036
cc_129 N_8_c_239_n N_Q_c_276_n 3.0124e-19 $X=0.837 $Y=0.153 $X2=0 $Y2=0
cc_130 N_8_c_239_n N_Q_c_284_n 3.0124e-19 $X=0.837 $Y=0.153 $X2=0 $Y2=0
cc_131 N_8_c_239_n N_Q_c_279_n 2.54113e-19 $X=0.837 $Y=0.153 $X2=0.464 $Y2=0.179
cc_132 N_8_c_240_n N_Q_c_279_n 6.27401e-19 $X=0.729 $Y=0.136 $X2=0.464 $Y2=0.179
cc_133 N_8_c_239_n N_Q_c_287_n 2.54113e-19 $X=0.837 $Y=0.153 $X2=0 $Y2=0
cc_134 N_8_c_246_p N_Q_c_287_n 5.42522e-19 $X=0.783 $Y=0.136 $X2=0 $Y2=0
cc_135 N_8_c_247_p N_Q_c_287_n 5.42522e-19 $X=0.837 $Y=0.136 $X2=0 $Y2=0
cc_136 N_8_c_239_n N_Q_c_281_n 3.83933e-19 $X=0.837 $Y=0.153 $X2=0.056 $Y2=0.054
cc_137 N_8_M7_g N_Q_c_291_n 3.24181e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_138 N_8_c_240_n N_Q_c_291_n 7.27236e-19 $X=0.729 $Y=0.136 $X2=0 $Y2=0
cc_139 N_8_c_239_n N_Q_c_293_n 4.26451e-19 $X=0.837 $Y=0.153 $X2=0.071 $Y2=0.216
cc_140 N_8_M8_g N_Q_c_294_n 3.24181e-19 $X=0.783 $Y=0.0675 $X2=0.056 $Y2=0.216
cc_141 N_8_c_246_p N_Q_c_294_n 7.27236e-19 $X=0.783 $Y=0.136 $X2=0.056 $Y2=0.216
cc_142 N_8_c_239_n N_Q_c_296_n 4.26451e-19 $X=0.837 $Y=0.153 $X2=0 $Y2=0
cc_143 N_8_M9_g N_Q_c_297_n 3.24181e-19 $X=0.837 $Y=0.0675 $X2=0.056 $Y2=0.216
cc_144 N_8_c_247_p N_Q_c_297_n 7.27236e-19 $X=0.837 $Y=0.136 $X2=0.056 $Y2=0.216
cc_145 N_8_c_239_n N_Q_c_282_n 3.65259e-19 $X=0.837 $Y=0.153 $X2=0.054 $Y2=0.036
cc_146 N_8_M7_g N_Q_c_300_n 3.50534e-19 $X=0.729 $Y=0.0675 $X2=0.054 $Y2=0.036
cc_147 N_8_c_240_n N_Q_c_300_n 5.44675e-19 $X=0.729 $Y=0.136 $X2=0.054 $Y2=0.036
cc_148 N_8_c_239_n N_Q_c_302_n 4.25288e-19 $X=0.837 $Y=0.153 $X2=0.054 $Y2=0.036
cc_149 N_8_M8_g N_Q_c_303_n 3.50534e-19 $X=0.783 $Y=0.0675 $X2=0.047 $Y2=0.036
cc_150 N_8_c_246_p N_Q_c_303_n 5.44675e-19 $X=0.783 $Y=0.136 $X2=0.047 $Y2=0.036
cc_151 N_8_c_239_n N_Q_c_305_n 4.25288e-19 $X=0.837 $Y=0.153 $X2=0.0505
+ $Y2=0.036
cc_152 N_8_M9_g N_Q_c_306_n 3.50534e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_153 N_8_c_247_p N_Q_c_306_n 5.44675e-19 $X=0.837 $Y=0.136 $X2=0 $Y2=0
cc_154 N_8_c_239_n Q 2.32153e-19 $X=0.837 $Y=0.153 $X2=0.054 $Y2=0.234
cc_155 N_8_c_247_p N_Q_c_309_n 0.00321652f $X=0.837 $Y=0.136 $X2=0.0505
+ $Y2=0.234
cc_156 N_8_c_192_n N_10_c_310_n 0.00119601f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.134
cc_157 N_8_c_197_n N_10_c_310_n 4.50844e-19 $X=0.45 $Y=0.036 $X2=0.351 $Y2=0.134
cc_158 N_8_c_198_n N_10_c_310_n 0.00394776f $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.134
cc_159 N_8_c_192_n N_11_c_318_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.134
cc_160 N_8_c_272_p N_11_c_318_n 0.00222776f $X=0.45 $Y=0.234 $X2=0.351 $Y2=0.134
cc_161 N_8_c_196_n N_11_c_318_n 0.00118584f $X=0.432 $Y=0.234 $X2=0.351
+ $Y2=0.134
cc_162 N_8_c_198_n N_11_c_318_n 5.72355e-19 $X=0.432 $Y=0.036 $X2=0.351
+ $Y2=0.134
cc_163 N_8_c_275_p N_11_c_318_n 0.00116187f $X=0.459 $Y=0.225 $X2=0.351
+ $Y2=0.134

* END of "./DHLx3_ASAP7_75t_SRAM.pex.sp.DHLX3_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DLLx1_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:28:15 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DLLx1_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DLLx1_ASAP7_75t_SRAM.pex.sp.pex"
* File: DLLx1_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:28:15 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DLLX1_ASAP7_75T_SRAM%CLK 2 5 7 12 14 17 VSS
c18 17 VSS 5.41721e-21 $X=0.081 $Y=0.1305
c19 14 VSS 0.00732563f $X=0.081 $Y=0.135
c20 12 VSS 0.00698013f $X=0.082 $Y=0.119
c21 5 VSS 0.0020626f $X=0.081 $Y=0.135
c22 2 VSS 0.0642213f $X=0.081 $Y=0.054
r23 16 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r24 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r25 12 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.126
r26 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DLLX1_ASAP7_75T_SRAM%4 2 7 10 13 15 17 20 22 25 28 29 30 33 37 44 49 51
+ 52 62 66 68 70 71 79 VSS
c44 96 VSS 1.06551e-19 $X=0.03 $Y=0.153
c45 95 VSS 6.89947e-19 $X=0.027 $Y=0.153
c46 79 VSS 0.00117224f $X=0.405 $Y=0.135
c47 71 VSS 0.0029117f $X=0.317 $Y=0.153
c48 70 VSS 0.00767547f $X=0.229 $Y=0.153
c49 68 VSS 0.00297348f $X=0.405 $Y=0.153
c50 66 VSS 0.00148441f $X=0.189 $Y=0.153
c51 62 VSS 9.21052e-19 $X=0.033 $Y=0.153
c52 52 VSS 0.00385436f $X=0.152 $Y=0.135
c53 51 VSS 4.1341e-19 $X=0.152 $Y=0.135
c54 49 VSS 0.00125241f $X=0.18 $Y=0.135
c55 47 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c56 46 VSS 0.00180216f $X=0.047 $Y=0.234
c57 44 VSS 0.00250477f $X=0.054 $Y=0.234
c58 42 VSS 0.00305101f $X=0.027 $Y=0.234
c59 40 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c60 39 VSS 0.00199699f $X=0.047 $Y=0.036
c61 37 VSS 0.00250477f $X=0.054 $Y=0.036
c62 35 VSS 0.00305101f $X=0.027 $Y=0.036
c63 34 VSS 9.44133e-19 $X=0.018 $Y=0.207
c64 33 VSS 0.00134027f $X=0.018 $Y=0.189
c65 32 VSS 8.82937e-19 $X=0.018 $Y=0.225
c66 30 VSS 0.00159315f $X=0.018 $Y=0.1125
c67 29 VSS 0.00142827f $X=0.018 $Y=0.081
c68 28 VSS 0.00144655f $X=0.018 $Y=0.144
c69 25 VSS 0.00453739f $X=0.056 $Y=0.216
c70 22 VSS 2.98509e-19 $X=0.071 $Y=0.216
c71 20 VSS 0.00456252f $X=0.056 $Y=0.054
c72 17 VSS 2.98509e-19 $X=0.071 $Y=0.054
c73 13 VSS 0.0015517f $X=0.405 $Y=0.135
c74 10 VSS 0.059003f $X=0.405 $Y=0.0675
c75 2 VSS 0.0639492f $X=0.135 $Y=0.054
r76 95 96 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r77 92 95 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r78 70 71 5.97531 $w=1.8e-08 $l=8.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.153 $X2=0.317 $Y2=0.153
r79 68 71 5.97531 $w=1.8e-08 $l=8.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.317 $Y2=0.153
r80 68 79 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r81 65 70 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.229 $Y2=0.153
r82 65 66 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.153 $X2=0.189
+ $Y2=0.153
r83 62 96 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r84 61 65 10.5926 $w=1.8e-08 $l=1.56e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.189 $Y2=0.153
r85 61 62 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r86 59 66 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.153
r87 51 52 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.152 $Y=0.135 $X2=0.152
+ $Y2=0.135
r88 49 59 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r89 49 51 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.152 $Y2=0.135
r90 46 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r91 44 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r92 42 46 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r93 39 40 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r94 37 40 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r95 35 39 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r96 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.207
r97 32 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r98 32 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.207
r99 31 92 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r100 31 33 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.189
r101 29 30 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.1125
r102 28 92 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r103 28 30 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1125
r104 27 35 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r105 27 29 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r106 25 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r107 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r108 20 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r109 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r110 13 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r111 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2295
r112 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r113 5 52 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.152 $Y2=0.135
r114 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r115 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DLLX1_ASAP7_75T_SRAM%D 2 5 7 12 16 VSS
c21 16 VSS 0.00596102f $X=0.297 $Y=0.135
c22 12 VSS 0.00848689f $X=0.297 $Y=0.1165
c23 5 VSS 0.0019062f $X=0.297 $Y=0.135
c24 2 VSS 0.061556f $X=0.297 $Y=0.0675
r25 12 16 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1165 $X2=0.297 $Y2=0.135
r26 5 16 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r27 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r28 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DLLX1_ASAP7_75T_SRAM%6 2 5 8 16 18 23 26 28 33 34 35 40 41 43 46 50 52
+ 54 55 59 71 72 75 76 78 VSS
c72 78 VSS 3.82279e-19 $X=0.243 $Y=0.216
c73 76 VSS 4.13588e-19 $X=0.243 $Y=0.126
c74 75 VSS 0.00265408f $X=0.243 $Y=0.117
c75 72 VSS 6.04312e-19 $X=0.513 $Y=0.18
c76 71 VSS 0.0601752f $X=0.513 $Y=0.18
c77 59 VSS 8.58425e-19 $X=0.351 $Y=0.135
c78 55 VSS 0.00132732f $X=0.45 $Y=0.189
c79 54 VSS 0.0053562f $X=0.414 $Y=0.189
c80 52 VSS 0.00307895f $X=0.513 $Y=0.189
c81 50 VSS 6.50668e-19 $X=0.351 $Y=0.189
c82 46 VSS 0.00221329f $X=0.243 $Y=0.189
c83 43 VSS 3.61041e-19 $X=0.243 $Y=0.225
c84 41 VSS 0.0018377f $X=0.216 $Y=0.234
c85 40 VSS 0.0051665f $X=0.198 $Y=0.234
c86 35 VSS 0.00483896f $X=0.234 $Y=0.234
c87 34 VSS 0.00184198f $X=0.216 $Y=0.036
c88 33 VSS 0.00552625f $X=0.198 $Y=0.036
c89 28 VSS 0.00484739f $X=0.234 $Y=0.036
c90 26 VSS 0.00641989f $X=0.16 $Y=0.216
c91 21 VSS 0.00625354f $X=0.16 $Y=0.054
c92 16 VSS 0.00212305f $X=0.464 $Y=0.179
c93 8 VSS 0.059718f $X=0.459 $Y=0.0405
c94 2 VSS 0.060362f $X=0.351 $Y=0.135
r95 77 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.207 $X2=0.243 $Y2=0.216
r96 75 76 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.117 $X2=0.243 $Y2=0.126
r97 71 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18 $X2=0.513
+ $Y2=0.18
r98 54 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.414
+ $Y=0.189 $X2=0.45 $Y2=0.189
r99 52 55 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.45 $Y2=0.189
r100 52 72 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r101 50 59 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.135
r102 49 54 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.414 $Y2=0.189
r103 49 50 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.189 $X2=0.351
+ $Y2=0.189
r104 46 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.207
r105 46 76 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.126
r106 45 49 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.351 $Y2=0.189
r107 45 46 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.189 $X2=0.243
+ $Y2=0.189
r108 43 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.216
r109 42 75 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.117
r110 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.216 $Y2=0.234
r111 37 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.198 $Y2=0.234
r112 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r113 35 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r114 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.216 $Y2=0.036
r115 30 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r116 28 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r117 28 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r118 26 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r119 23 26 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r120 21 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r121 18 21 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r122 16 71 42.2917 $w=2.4e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08 $X=0.464
+ $Y=0.179 $X2=0.513 $Y2=0.179
r123 11 16 3.57143 $w=2.8e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.179 $X2=0.464 $Y2=0.179
r124 8 11 518.891 $w=2e-08 $l=1.385e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.179
r125 2 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r126 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
.ends

.subckt PM_DLLX1_ASAP7_75T_SRAM%7 2 5 7 9 12 14 17 21 24 25 29 35 36 37 38 45 46
+ VSS
c25 46 VSS 0.00411848f $X=0.612 $Y=0.234
c26 45 VSS 0.00236179f $X=0.621 $Y=0.234
c27 40 VSS 4.66533e-19 $X=0.621 $Y=0.214
c28 39 VSS 2.58319e-19 $X=0.621 $Y=0.203
c29 38 VSS 6.12455e-19 $X=0.621 $Y=0.2
c30 37 VSS 6.7107e-19 $X=0.621 $Y=0.165
c31 36 VSS 4.81665e-19 $X=0.621 $Y=0.14
c32 35 VSS 8.07335e-19 $X=0.621 $Y=0.122
c33 34 VSS 5.25258e-19 $X=0.621 $Y=0.106
c34 33 VSS 0.00187639f $X=0.621 $Y=0.097
c35 32 VSS 7.90142e-19 $X=0.621 $Y=0.225
c36 30 VSS 8.17537e-19 $X=0.587 $Y=0.036
c37 29 VSS 0.00649884f $X=0.58 $Y=0.036
c38 25 VSS 0.0022245f $X=0.522 $Y=0.036
c39 24 VSS 0.00491847f $X=0.612 $Y=0.036
c40 21 VSS 5.81526e-19 $X=0.513 $Y=0.082
c41 17 VSS 0.00494953f $X=0.592 $Y=0.2295
c42 12 VSS 0.00511574f $X=0.592 $Y=0.0405
c43 5 VSS 0.00256679f $X=0.513 $Y=0.082
c44 2 VSS 0.0581876f $X=0.513 $Y=0.0405
r45 46 47 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r46 45 47 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r47 42 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.612 $Y2=0.234
r48 39 40 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.214
r49 38 39 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.2 $X2=0.621 $Y2=0.203
r50 37 38 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.2
r51 36 37 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r52 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r53 34 35 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.106 $X2=0.621 $Y2=0.122
r54 33 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.097 $X2=0.621 $Y2=0.106
r55 32 45 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.234
r56 32 40 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.214
r57 31 33 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.097
r58 29 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.58
+ $Y=0.036 $X2=0.587 $Y2=0.036
r59 27 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.587 $Y2=0.036
r60 25 29 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.58 $Y2=0.036
r61 24 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r62 24 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.594 $Y2=0.036
r63 19 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.513 $Y=0.045 $X2=0.522 $Y2=0.036
r64 19 21 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.082
r65 17 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r66 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r67 12 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036 $X2=0.594
+ $Y2=0.036
r68 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.592 $Y2=0.0405
r69 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.082 $X2=0.513
+ $Y2=0.082
r70 5 7 552.609 $w=2e-08 $l=1.475e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.082 $X2=0.513 $Y2=0.2295
r71 2 5 155.48 $w=2e-08 $l=4.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.082
.ends

.subckt PM_DLLX1_ASAP7_75T_SRAM%8 2 7 10 15 17 22 25 29 30 33 38 39 40 43 46 47 51
+ 53 54 58 61 64 66 67 74 86 VSS
c55 88 VSS 4.52133e-19 $X=0.459 $Y=0.214
c56 87 VSS 5.73001e-20 $X=0.459 $Y=0.203
c57 86 VSS 2.69603e-19 $X=0.459 $Y=0.2
c58 74 VSS 0.00254734f $X=0.729 $Y=0.136
c59 67 VSS 0.00410379f $X=0.628 $Y=0.153
c60 66 VSS 0.0014648f $X=0.527 $Y=0.153
c61 64 VSS 0.0083017f $X=0.729 $Y=0.153
c62 61 VSS 3.75508e-19 $X=0.459 $Y=0.153
c63 58 VSS 3.21606e-19 $X=0.459 $Y=0.225
c64 57 VSS 2.32827e-19 $X=0.459 $Y=0.131
c65 54 VSS 3.60459e-20 $X=0.522 $Y=0.131
c66 53 VSS 0.00173419f $X=0.504 $Y=0.131
c67 51 VSS 0.00147804f $X=0.566 $Y=0.131
c68 48 VSS 5.04027e-19 $X=0.459 $Y=0.106
c69 47 VSS 2.74504e-19 $X=0.459 $Y=0.097
c70 46 VSS 3.18939e-19 $X=0.459 $Y=0.122
c71 43 VSS 0.00271748f $X=0.432 $Y=0.036
c72 40 VSS 0.00636101f $X=0.45 $Y=0.036
c73 39 VSS 0.00146362f $X=0.414 $Y=0.234
c74 38 VSS 0.00368178f $X=0.396 $Y=0.234
c75 33 VSS 0.00571919f $X=0.45 $Y=0.234
c76 32 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c77 29 VSS 0.00348747f $X=0.378 $Y=0.2025
c78 24 VSS 5.36734e-19 $X=0.432 $Y=0.0405
c79 13 VSS 0.00369274f $X=0.729 $Y=0.136
c80 10 VSS 0.0655607f $X=0.729 $Y=0.0675
c81 5 VSS 0.00312272f $X=0.567 $Y=0.131
c82 2 VSS 0.0616253f $X=0.567 $Y=0.0405
r83 87 88 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.203 $X2=0.459 $Y2=0.214
r84 86 87 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.2 $X2=0.459 $Y2=0.203
r85 85 86 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.2
r86 66 67 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.628 $Y2=0.153
r87 64 67 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M2 $thickness=3.6e-08 $X=0.729
+ $Y=0.153 $X2=0.628 $Y2=0.153
r88 64 74 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.729 $Y=0.153 $X2=0.729
+ $Y2=0.153
r89 61 85 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.459 $Y2=0.165
r90 60 66 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.527 $Y2=0.153
r91 60 61 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.459 $Y=0.153 $X2=0.459
+ $Y2=0.153
r92 58 88 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r93 56 61 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.153
r94 56 57 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r95 53 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r96 51 54 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.566
+ $Y=0.131 $X2=0.522 $Y2=0.131
r97 49 57 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r98 49 53 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.504 $Y2=0.131
r99 47 48 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.097 $X2=0.459 $Y2=0.106
r100 46 57 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r101 46 48 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.106
r102 45 47 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.097
r103 42 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r104 40 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r105 40 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.432 $Y2=0.036
r106 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r107 35 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r108 33 58 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r109 33 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.414 $Y2=0.234
r110 30 32 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r111 29 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r112 26 32 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r113 26 29 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r114 25 29 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r115 22 24 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r116 21 43 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r117 18 24 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r118 18 21 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r119 17 21 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r120 13 74 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.729 $Y=0.136 $X2=0.729
+ $Y2=0.136
r121 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.136 $X2=0.729 $Y2=0.2025
r122 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.136
r123 5 51 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.566 $Y=0.131 $X2=0.566
+ $Y2=0.131
r124 5 7 369.03 $w=2e-08 $l=9.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.131 $X2=0.567 $Y2=0.2295
r125 2 5 339.058 $w=2e-08 $l=9.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.131
.ends

.subckt PM_DLLX1_ASAP7_75T_SRAM%Q 1 6 9 13 21 23 29 VSS
c6 29 VSS 0.00433882f $X=0.774 $Y=0.234
c7 28 VSS 0.00278493f $X=0.783 $Y=0.234
c8 23 VSS 0.00419073f $X=0.783 $Y=0.2
c9 21 VSS 0.00259959f $X=0.783 $Y=0.081
c10 19 VSS 0.00149091f $X=0.783 $Y=0.225
c11 14 VSS 0.00648051f $X=0.756 $Y=0.036
c12 13 VSS 0.00167221f $X=0.756 $Y=0.036
c13 11 VSS 0.00666612f $X=0.774 $Y=0.036
c14 9 VSS 0.0070175f $X=0.754 $Y=0.2025
c15 4 VSS 3.30876e-19 $X=0.754 $Y=0.0675
r16 29 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.234 $X2=0.7785 $Y2=0.234
r17 28 30 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.234 $X2=0.7785 $Y2=0.234
r18 25 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.774 $Y2=0.234
r19 22 23 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.106 $X2=0.783 $Y2=0.2
r20 21 22 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.081 $X2=0.783 $Y2=0.106
r21 19 28 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.225 $X2=0.783 $Y2=0.234
r22 19 23 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.225 $X2=0.783 $Y2=0.2
r23 18 21 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.045 $X2=0.783 $Y2=0.081
r24 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r25 11 18 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.774 $Y=0.036 $X2=0.783 $Y2=0.045
r26 11 13 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.036 $X2=0.756 $Y2=0.036
r27 9 25 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234 $X2=0.756
+ $Y2=0.234
r28 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.2025 $X2=0.754 $Y2=0.2025
r29 4 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.756
+ $Y=0.0675 $X2=0.756 $Y2=0.036
r30 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.0675 $X2=0.754 $Y2=0.0675
.ends

.subckt PM_DLLX1_ASAP7_75T_SRAM%10 1 6 9 VSS
c7 9 VSS 0.0266424f $X=0.38 $Y=0.0675
c8 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c9 4 VSS 3.22674e-19 $X=0.322 $Y=0.0675
r10 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r12 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DLLX1_ASAP7_75T_SRAM%11 1 6 9 VSS
c9 9 VSS 0.0211025f $X=0.488 $Y=0.2295
c10 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c11 4 VSS 2.84146e-19 $X=0.43 $Y=0.2295
r12 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r13 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DLLX1_ASAP7_75T_SRAM%12 1 2 VSS
c0 1 VSS 0.00220425f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DLLX1_ASAP7_75T_SRAM%13 1 2 VSS
c1 1 VSS 0.00201018f $X=0.341 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends


* END of "./DLLx1_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DLLx1_ASAP7_75t_SRAM  VSS VDD CLK D Q
* 
* Q	Q
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_10_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_4_M3_g N_10_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_12_M4_d N_6_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_12_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_Q_M7_d N_8_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M8 VDD N_CLK_M8_g N_4_M8_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M9 N_6_M9_d N_4_M9_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
M10 N_13_M10_d N_D_M10_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_8_M11_d N_6_M11_g N_13_M11_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M12 N_11_M12_d N_4_M12_g N_8_M12_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M13 VDD N_7_M13_g N_11_M13_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M14 N_7_M14_d N_8_M14_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M15 N_Q_M15_d N_8_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
*
* 
* .include "DLLx1_ASAP7_75t_SRAM.pex.sp.DLLX1_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DLLx1_ASAP7_75t_SRAM.pex.sp.DLLX1_ASAP7_75T_SRAM.pxi"
* File: DLLx1_ASAP7_75t_SRAM.pex.sp.DLLX1_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:28:15 2017
* 
x_PM_DLLX1_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_11_p N_CLK_M8_g CLK N_CLK_c_3_p
+ N_CLK_c_4_p VSS PM_DLLX1_ASAP7_75T_SRAM%CLK
x_PM_DLLX1_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M9_g N_4_M3_g N_4_c_38_p N_4_M12_g
+ N_4_M0_s N_4_c_20_n N_4_M8_s N_4_c_21_n N_4_c_22_n N_4_c_23_n N_4_c_24_n
+ N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_48_p N_4_c_28_n N_4_c_29_n N_4_c_30_n
+ N_4_c_31_n N_4_c_53_p N_4_c_32_n N_4_c_36_p N_4_c_40_p VSS
+ PM_DLLX1_ASAP7_75T_SRAM%4
x_PM_DLLX1_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_64_n N_D_M10_g D N_D_c_69_p VSS
+ PM_DLLX1_ASAP7_75T_SRAM%D
x_PM_DLLX1_ASAP7_75T_SRAM%6 N_6_c_87_n N_6_M11_g N_6_M4_g N_6_c_90_n N_6_M1_d
+ N_6_M9_d N_6_c_91_n N_6_c_92_n N_6_c_84_n N_6_c_94_n N_6_c_95_n N_6_c_85_n
+ N_6_c_97_n N_6_c_109_n N_6_c_98_n N_6_c_111_n N_6_c_141_p N_6_c_100_n
+ N_6_c_131_p N_6_c_103_n N_6_c_119_p N_6_c_120_p N_6_c_86_n N_6_c_116_n
+ N_6_c_117_n VSS PM_DLLX1_ASAP7_75T_SRAM%6
x_PM_DLLX1_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_160_n N_7_M13_g N_7_M6_d N_7_c_161_n
+ N_7_M14_d N_7_c_162_n N_7_c_169_p N_7_c_179_p N_7_c_168_p N_7_c_167_p
+ N_7_c_178_p N_7_c_171_p N_7_c_174_p N_7_c_163_n N_7_c_180_p N_7_c_165_n VSS
+ PM_DLLX1_ASAP7_75T_SRAM%7
x_PM_DLLX1_ASAP7_75T_SRAM%8 N_8_M6_g N_8_M14_g N_8_M7_g N_8_M15_g N_8_M3_d N_8_M4_s
+ N_8_M11_d N_8_c_181_n N_8_M12_s N_8_c_194_n N_8_c_188_n N_8_c_182_n
+ N_8_c_189_n N_8_c_197_n N_8_c_184_n N_8_c_199_n N_8_c_200_n N_8_c_201_n
+ N_8_c_202_n N_8_c_235_p N_8_c_185_n N_8_c_220_n N_8_c_186_n N_8_c_221_n
+ N_8_c_224_n N_8_c_208_n VSS PM_DLLX1_ASAP7_75T_SRAM%8
x_PM_DLLX1_ASAP7_75T_SRAM%Q N_Q_M7_d N_Q_M15_d N_Q_c_238_n N_Q_c_236_n Q
+ N_Q_c_240_n N_Q_c_237_n VSS PM_DLLX1_ASAP7_75T_SRAM%Q
x_PM_DLLX1_ASAP7_75T_SRAM%10 N_10_M2_d N_10_M3_s N_10_c_242_n VSS
+ PM_DLLX1_ASAP7_75T_SRAM%10
x_PM_DLLX1_ASAP7_75T_SRAM%11 N_11_M12_d N_11_M13_s N_11_c_250_n VSS
+ PM_DLLX1_ASAP7_75T_SRAM%11
x_PM_DLLX1_ASAP7_75T_SRAM%12 N_12_M5_s N_12_M4_d VSS PM_DLLX1_ASAP7_75T_SRAM%12
x_PM_DLLX1_ASAP7_75T_SRAM%13 N_13_M11_s N_13_M10_d VSS PM_DLLX1_ASAP7_75T_SRAM%13
cc_1 N_CLK_M0_g N_4_M1_g 0.0027643f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_20_n 2.66516e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 N_CLK_c_3_p N_4_c_21_n 2.66516e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.216
cc_4 N_CLK_c_4_p N_4_c_22_n 0.00126555f $X=0.081 $Y=0.1305 $X2=0.018 $Y2=0.144
cc_5 CLK N_4_c_23_n 3.98992e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.081
cc_6 CLK N_4_c_24_n 0.00126555f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.1125
cc_7 N_CLK_c_3_p N_4_c_25_n 0.00127356f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.189
cc_8 CLK N_4_c_26_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_3_p N_4_c_27_n 4.98319e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_4_p N_4_c_28_n 4.17e-19 $X=0.081 $Y=0.1305 $X2=0.152 $Y2=0.135
cc_11 N_CLK_c_11_p N_4_c_29_n 0.00116357f $X=0.081 $Y=0.135 $X2=0.152 $Y2=0.135
cc_12 N_CLK_c_3_p N_4_c_30_n 0.00122788f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.153
cc_13 N_CLK_c_3_p N_4_c_31_n 0.00197837f $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.153
cc_14 CLK N_4_c_32_n 5.08945e-19 $X=0.082 $Y=0.119 $X2=0.229 $Y2=0.153
cc_15 N_CLK_c_3_p N_4_c_32_n 0.00150524f $X=0.081 $Y=0.135 $X2=0.229 $Y2=0.153
cc_16 CLK N_6_c_84_n 6.45949e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.189
cc_17 N_CLK_c_3_p N_6_c_85_n 6.45949e-19 $X=0.081 $Y=0.135 $X2=0.0505 $Y2=0.036
cc_18 CLK N_6_c_86_n 7.98675e-19 $X=0.082 $Y=0.119 $X2=0.152 $Y2=0.135
cc_19 N_4_M3_g N_D_M2_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_20 N_4_c_29_n N_D_c_64_n 2.01856e-19 $X=0.152 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 N_4_c_36_p D 0.00117371f $X=0.317 $Y=0.153 $X2=0.082 $Y2=0.119
cc_22 N_4_M3_g N_6_c_87_n 0.00355599f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_23 N_4_c_38_p N_6_c_87_n 0.00101396f $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.054
cc_24 N_4_M3_g N_6_M4_g 0.00355599f $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_25 N_4_c_40_p N_6_c_90_n 3.2936e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.126
cc_26 N_4_c_31_n N_6_c_91_n 0.00243501f $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_27 N_4_c_36_p N_6_c_92_n 2.3925e-19 $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_28 N_4_c_28_n N_6_c_84_n 9.58415e-19 $X=0.152 $Y=0.135 $X2=0 $Y2=0
cc_29 N_4_c_32_n N_6_c_94_n 2.3925e-19 $X=0.229 $Y=0.153 $X2=0 $Y2=0
cc_30 N_4_c_36_p N_6_c_95_n 2.75285e-19 $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_31 N_4_c_31_n N_6_c_85_n 0.00467935f $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_32 N_4_c_32_n N_6_c_97_n 2.75285e-19 $X=0.229 $Y=0.153 $X2=0 $Y2=0
cc_33 N_4_c_48_p N_6_c_98_n 0.00396181f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_34 N_4_c_36_p N_6_c_98_n 0.00119509f $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_35 N_4_c_31_n N_6_c_100_n 3.89771e-19 $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_36 N_4_c_36_p N_6_c_100_n 0.0160263f $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_37 N_4_c_40_p N_6_c_100_n 8.49272e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_53_p N_6_c_103_n 0.00115166f $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_40_p N_6_c_103_n 0.00433569f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_41 N_4_c_40_p N_8_c_181_n 0.00195725f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_42 N_4_M3_g N_8_c_182_n 2.63086e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_4_c_40_p N_8_c_182_n 0.00122664f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_44 N_4_c_40_p N_8_c_184_n 0.00419136f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_45 N_4_c_40_p N_8_c_185_n 2.60642e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_53_p N_8_c_186_n 9.16428e-19 $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_36_p N_10_c_242_n 8.32437e-19 $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_48 N_D_M2_g N_6_c_87_n 0.00341068f $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_49 N_D_c_64_n N_6_c_87_n 0.00101372f $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_50 D N_6_c_92_n 0.00115278f $X=0.297 $Y=0.1165 $X2=0.018 $Y2=0.144
cc_51 N_D_c_69_p N_6_c_95_n 0.00115278f $X=0.297 $Y=0.135 $X2=0.027 $Y2=0.036
cc_52 N_D_c_69_p N_6_c_109_n 0.00115278f $X=0.297 $Y=0.135 $X2=0.054 $Y2=0.234
cc_53 D N_6_c_98_n 0.00124619f $X=0.297 $Y=0.1165 $X2=0.047 $Y2=0.234
cc_54 D N_6_c_111_n 0.00216863f $X=0.297 $Y=0.1165 $X2=0.152 $Y2=0.135
cc_55 D N_6_c_100_n 8.86605e-19 $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_56 N_D_c_69_p N_6_c_100_n 3.97512e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_57 D N_6_c_103_n 0.00216863f $X=0.297 $Y=0.1165 $X2=0.189 $Y2=0.144
cc_58 D N_6_c_86_n 0.00115278f $X=0.297 $Y=0.1165 $X2=0.152 $Y2=0.135
cc_59 D N_6_c_116_n 0.00115278f $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_60 N_D_c_69_p N_6_c_117_n 0.00115278f $X=0.297 $Y=0.135 $X2=0.405 $Y2=0.135
cc_61 N_D_c_69_p N_8_c_181_n 3.88702e-19 $X=0.297 $Y=0.135 $X2=0.018 $Y2=0.081
cc_62 N_D_c_69_p N_8_c_188_n 8.77202e-19 $X=0.297 $Y=0.135 $X2=0.054 $Y2=0.036
cc_63 D N_8_c_189_n 2.05539e-19 $X=0.297 $Y=0.1165 $X2=0.0505 $Y2=0.036
cc_64 D N_10_c_242_n 0.00428733f $X=0.297 $Y=0.1165 $X2=0.405 $Y2=0.0675
cc_65 N_D_c_69_p N_13_M11_s 3.05674e-19 $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_66 N_6_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_67 N_6_c_119_p N_7_M5_g 0.00199227f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_68 N_6_c_120_p N_7_M5_g 4.91626e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_69 N_6_c_119_p N_7_c_160_n 4.44368e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.135
cc_70 N_6_c_119_p N_7_c_161_n 5.31675e-19 $X=0.513 $Y=0.18 $X2=0.082 $Y2=0.119
cc_71 N_6_c_119_p N_7_c_162_n 0.00169036f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.1305
cc_72 N_6_c_119_p N_7_c_163_n 0.00339185f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_73 N_6_c_120_p N_7_c_163_n 6.11658e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_74 N_6_c_119_p N_7_c_165_n 5.97916e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_75 N_6_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_76 N_6_c_119_p N_8_M6_g 0.00305655f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_77 N_6_c_100_n N_8_c_181_n 2.84357e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_78 N_6_c_103_n N_8_c_181_n 0.00130164f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_79 N_6_c_131_p N_8_c_194_n 7.16323e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_80 N_6_c_100_n N_8_c_188_n 5.53186e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_81 N_6_c_131_p N_8_c_189_n 3.48842e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_82 N_6_c_131_p N_8_c_197_n 2.01793e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_83 N_6_M4_g N_8_c_184_n 2.93184e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_84 N_6_M4_g N_8_c_199_n 3.72919e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_85 N_6_c_119_p N_8_c_200_n 4.41338e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_86 N_6_c_119_p N_8_c_201_n 7.92645e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_87 N_6_c_120_p N_8_c_202_n 0.00100546f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_88 N_6_M4_g N_8_c_185_n 2.27241e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_89 N_6_c_141_p N_8_c_185_n 2.46239e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_90 N_6_c_141_p N_8_c_186_n 0.00694438f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_91 N_6_c_119_p N_8_c_186_n 0.00195448f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_92 N_6_c_120_p N_8_c_186_n 2.84312e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_93 N_6_c_90_n N_8_c_208_n 0.00271026f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_94 N_6_c_141_p N_8_c_208_n 6.73646e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_95 N_6_c_119_p N_8_c_208_n 5.95032e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_96 N_6_c_120_p N_8_c_208_n 0.00182777f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_97 N_6_c_87_n N_10_c_242_n 0.00639848f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_98 N_6_c_103_n N_10_c_242_n 0.00135407f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_99 N_6_c_119_p N_11_M13_s 2.34172e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.216
cc_100 N_6_M4_g N_11_c_250_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_101 N_6_c_90_n N_11_c_250_n 0.0013957f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_102 N_6_c_131_p N_11_c_250_n 7.09553e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_103 N_6_c_119_p N_11_c_250_n 0.00230185f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_104 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_105 N_7_c_167_p N_8_M6_g 4.17397e-19 $X=0.58 $Y=0.036 $X2=0.135 $Y2=0.054
cc_106 N_7_c_168_p N_8_c_189_n 0.00177955f $X=0.522 $Y=0.036 $X2=0.0505
+ $Y2=0.036
cc_107 N_7_c_169_p N_8_c_199_n 0.00177955f $X=0.513 $Y=0.082 $X2=0.0505
+ $Y2=0.234
cc_108 N_7_c_167_p N_8_c_200_n 6.9494e-19 $X=0.58 $Y=0.036 $X2=0.152 $Y2=0.135
cc_109 N_7_c_171_p N_8_c_200_n 9.49516e-19 $X=0.621 $Y=0.14 $X2=0.152 $Y2=0.135
cc_110 N_7_M5_g N_8_c_202_n 4.06683e-19 $X=0.513 $Y=0.0405 $X2=0 $Y2=0
cc_111 N_7_c_169_p N_8_c_202_n 0.00116089f $X=0.513 $Y=0.082 $X2=0 $Y2=0
cc_112 N_7_c_174_p N_8_c_220_n 3.80483e-19 $X=0.621 $Y=0.165 $X2=0.189 $Y2=0.153
cc_113 N_7_c_161_n N_8_c_221_n 2.11538e-19 $X=0.592 $Y=0.0405 $X2=0.405
+ $Y2=0.153
cc_114 N_7_c_174_p N_8_c_221_n 8.70427e-19 $X=0.621 $Y=0.165 $X2=0.405 $Y2=0.153
cc_115 N_7_c_165_n N_8_c_221_n 5.94743e-19 $X=0.612 $Y=0.234 $X2=0.405 $Y2=0.153
cc_116 N_7_c_178_p N_8_c_224_n 0.00117009f $X=0.621 $Y=0.122 $X2=0 $Y2=0
cc_117 N_7_c_179_p N_Q_c_236_n 2.34097e-19 $X=0.612 $Y=0.036 $X2=0.405 $Y2=0.135
cc_118 N_7_c_180_p N_Q_c_237_n 2.15386e-19 $X=0.621 $Y=0.234 $X2=0.018 $Y2=0.081
cc_119 N_8_c_224_n N_Q_c_238_n 0.00114532f $X=0.729 $Y=0.136 $X2=0.405
+ $Y2=0.0675
cc_120 N_8_M7_g N_Q_c_236_n 2.22123e-19 $X=0.729 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_121 N_8_c_220_n N_Q_c_240_n 2.31367e-19 $X=0.729 $Y=0.153 $X2=0.056 $Y2=0.216
cc_122 N_8_c_224_n N_Q_c_240_n 0.00387106f $X=0.729 $Y=0.136 $X2=0.056 $Y2=0.216
cc_123 N_8_c_181_n N_10_c_242_n 0.00119636f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_124 N_8_c_189_n N_10_c_242_n 4.50844e-19 $X=0.45 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_125 N_8_c_197_n N_10_c_242_n 0.00394776f $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_126 N_8_c_181_n N_11_c_250_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_127 N_8_c_194_n N_11_c_250_n 0.00343017f $X=0.45 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_128 N_8_c_197_n N_11_c_250_n 5.72355e-19 $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_129 N_8_c_235_p N_11_c_250_n 0.00116187f $X=0.459 $Y=0.225 $X2=0.405
+ $Y2=0.0675

* END of "./DLLx1_ASAP7_75t_SRAM.pex.sp.DLLX1_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DLLx2_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:28:38 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DLLx2_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DLLx2_ASAP7_75t_SRAM.pex.sp.pex"
* File: DLLx2_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:28:38 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DLLX2_ASAP7_75T_SRAM%CLK 2 5 7 12 14 17 VSS
c18 17 VSS 5.41721e-21 $X=0.081 $Y=0.1305
c19 14 VSS 0.00732563f $X=0.081 $Y=0.135
c20 12 VSS 0.00698013f $X=0.082 $Y=0.119
c21 5 VSS 0.0020626f $X=0.081 $Y=0.135
c22 2 VSS 0.062963f $X=0.081 $Y=0.054
r23 16 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r24 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r25 12 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.126
r26 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DLLX2_ASAP7_75T_SRAM%4 2 7 10 13 15 17 20 22 25 28 29 30 33 37 44 49 51
+ 52 62 66 68 70 71 79 VSS
c44 96 VSS 1.06551e-19 $X=0.03 $Y=0.153
c45 95 VSS 6.89947e-19 $X=0.027 $Y=0.153
c46 79 VSS 0.00117246f $X=0.405 $Y=0.135
c47 71 VSS 0.0029117f $X=0.317 $Y=0.153
c48 70 VSS 0.00767547f $X=0.229 $Y=0.153
c49 68 VSS 0.00297348f $X=0.405 $Y=0.153
c50 66 VSS 0.00148441f $X=0.189 $Y=0.153
c51 62 VSS 9.21052e-19 $X=0.033 $Y=0.153
c52 52 VSS 0.00385436f $X=0.152 $Y=0.135
c53 51 VSS 4.1341e-19 $X=0.152 $Y=0.135
c54 49 VSS 0.00125241f $X=0.18 $Y=0.135
c55 47 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c56 46 VSS 0.00180216f $X=0.047 $Y=0.234
c57 44 VSS 0.00250477f $X=0.054 $Y=0.234
c58 42 VSS 0.00305101f $X=0.027 $Y=0.234
c59 40 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c60 39 VSS 0.00199699f $X=0.047 $Y=0.036
c61 37 VSS 0.00250477f $X=0.054 $Y=0.036
c62 35 VSS 0.00305101f $X=0.027 $Y=0.036
c63 34 VSS 9.44133e-19 $X=0.018 $Y=0.207
c64 33 VSS 0.00134027f $X=0.018 $Y=0.189
c65 32 VSS 8.82937e-19 $X=0.018 $Y=0.225
c66 30 VSS 0.00159315f $X=0.018 $Y=0.1125
c67 29 VSS 0.00142827f $X=0.018 $Y=0.081
c68 28 VSS 0.00144655f $X=0.018 $Y=0.144
c69 25 VSS 0.00453739f $X=0.056 $Y=0.216
c70 22 VSS 2.98509e-19 $X=0.071 $Y=0.216
c71 20 VSS 0.00456252f $X=0.056 $Y=0.054
c72 17 VSS 2.98509e-19 $X=0.071 $Y=0.054
c73 13 VSS 0.0015517f $X=0.405 $Y=0.135
c74 10 VSS 0.059003f $X=0.405 $Y=0.0675
c75 2 VSS 0.0627154f $X=0.135 $Y=0.054
r76 95 96 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r77 92 95 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r78 70 71 5.97531 $w=1.8e-08 $l=8.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.153 $X2=0.317 $Y2=0.153
r79 68 71 5.97531 $w=1.8e-08 $l=8.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.317 $Y2=0.153
r80 68 79 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r81 65 70 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.229 $Y2=0.153
r82 65 66 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.153 $X2=0.189
+ $Y2=0.153
r83 62 96 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r84 61 65 10.5926 $w=1.8e-08 $l=1.56e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.189 $Y2=0.153
r85 61 62 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r86 59 66 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.153
r87 51 52 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.152 $Y=0.135 $X2=0.152
+ $Y2=0.135
r88 49 59 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r89 49 51 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.152 $Y2=0.135
r90 46 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r91 44 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r92 42 46 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r93 39 40 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r94 37 40 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r95 35 39 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r96 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.207
r97 32 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r98 32 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.207
r99 31 92 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r100 31 33 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.189
r101 29 30 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.1125
r102 28 92 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r103 28 30 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1125
r104 27 35 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r105 27 29 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r106 25 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r107 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r108 20 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r109 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r110 13 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r111 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2295
r112 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r113 5 52 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.152 $Y2=0.135
r114 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r115 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DLLX2_ASAP7_75T_SRAM%D 2 5 7 12 16 VSS
c21 16 VSS 0.00596102f $X=0.297 $Y=0.135
c22 12 VSS 0.00848689f $X=0.297 $Y=0.1165
c23 5 VSS 0.0019062f $X=0.297 $Y=0.135
c24 2 VSS 0.061556f $X=0.297 $Y=0.0675
r25 12 16 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1165 $X2=0.297 $Y2=0.135
r26 5 16 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r27 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r28 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DLLX2_ASAP7_75T_SRAM%6 2 5 8 16 18 23 26 28 33 34 35 40 41 43 46 50 52
+ 54 55 59 71 72 75 76 78 VSS
c74 78 VSS 3.82279e-19 $X=0.243 $Y=0.216
c75 76 VSS 4.13588e-19 $X=0.243 $Y=0.126
c76 75 VSS 0.00265408f $X=0.243 $Y=0.117
c77 72 VSS 6.21924e-19 $X=0.513 $Y=0.18
c78 71 VSS 0.0589952f $X=0.513 $Y=0.18
c79 59 VSS 8.58425e-19 $X=0.351 $Y=0.135
c80 55 VSS 0.00132732f $X=0.45 $Y=0.189
c81 54 VSS 0.0053562f $X=0.414 $Y=0.189
c82 52 VSS 0.00304981f $X=0.513 $Y=0.189
c83 50 VSS 6.50668e-19 $X=0.351 $Y=0.189
c84 46 VSS 0.00221329f $X=0.243 $Y=0.189
c85 43 VSS 3.61041e-19 $X=0.243 $Y=0.225
c86 41 VSS 0.0018377f $X=0.216 $Y=0.234
c87 40 VSS 0.0051665f $X=0.198 $Y=0.234
c88 35 VSS 0.00483896f $X=0.234 $Y=0.234
c89 34 VSS 0.00184198f $X=0.216 $Y=0.036
c90 33 VSS 0.00552625f $X=0.198 $Y=0.036
c91 28 VSS 0.00484739f $X=0.234 $Y=0.036
c92 26 VSS 0.00641989f $X=0.16 $Y=0.216
c93 21 VSS 0.00625354f $X=0.16 $Y=0.054
c94 16 VSS 0.00212305f $X=0.464 $Y=0.179
c95 8 VSS 0.059718f $X=0.459 $Y=0.0405
c96 2 VSS 0.060362f $X=0.351 $Y=0.135
r97 77 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.207 $X2=0.243 $Y2=0.216
r98 75 76 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.117 $X2=0.243 $Y2=0.126
r99 71 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18 $X2=0.513
+ $Y2=0.18
r100 54 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.414
+ $Y=0.189 $X2=0.45 $Y2=0.189
r101 52 55 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.45 $Y2=0.189
r102 52 72 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r103 50 59 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.135
r104 49 54 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.414 $Y2=0.189
r105 49 50 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.189 $X2=0.351
+ $Y2=0.189
r106 46 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.207
r107 46 76 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.126
r108 45 49 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.351 $Y2=0.189
r109 45 46 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.189 $X2=0.243
+ $Y2=0.189
r110 43 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.216
r111 42 75 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.117
r112 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.216 $Y2=0.234
r113 37 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.198 $Y2=0.234
r114 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r115 35 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r116 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.216 $Y2=0.036
r117 30 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r118 28 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r119 28 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r120 26 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r121 23 26 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r122 21 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r123 18 21 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r124 16 71 42.2917 $w=2.4e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08 $X=0.464
+ $Y=0.179 $X2=0.513 $Y2=0.179
r125 11 16 3.57143 $w=2.8e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.179 $X2=0.464 $Y2=0.179
r126 8 11 518.891 $w=2e-08 $l=1.385e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.179
r127 2 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r128 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
.ends

.subckt PM_DLLX2_ASAP7_75T_SRAM%7 2 5 7 9 12 14 17 21 24 25 29 33 34 35 36 37 38 39
+ 45 46 VSS
c31 46 VSS 0.00411848f $X=0.612 $Y=0.234
c32 45 VSS 0.00208935f $X=0.621 $Y=0.234
c33 40 VSS 3.32784e-19 $X=0.621 $Y=0.214
c34 39 VSS 4.44772e-19 $X=0.621 $Y=0.203
c35 38 VSS 3.45124e-20 $X=0.621 $Y=0.167
c36 37 VSS 8.18444e-19 $X=0.621 $Y=0.165
c37 36 VSS 5.62221e-19 $X=0.621 $Y=0.14
c38 35 VSS 0.00100849f $X=0.621 $Y=0.122
c39 34 VSS 1.64643e-19 $X=0.621 $Y=0.097
c40 33 VSS 7.03241e-19 $X=0.621 $Y=0.09
c41 32 VSS 5.59839e-19 $X=0.621 $Y=0.225
c42 30 VSS 8.17537e-19 $X=0.587 $Y=0.036
c43 29 VSS 0.00649884f $X=0.58 $Y=0.036
c44 25 VSS 0.0022245f $X=0.522 $Y=0.036
c45 24 VSS 0.00465365f $X=0.612 $Y=0.036
c46 21 VSS 5.81526e-19 $X=0.513 $Y=0.082
c47 17 VSS 0.00441907f $X=0.592 $Y=0.2295
c48 12 VSS 0.00458532f $X=0.592 $Y=0.0405
c49 5 VSS 0.00256679f $X=0.513 $Y=0.082
c50 2 VSS 0.0581876f $X=0.513 $Y=0.0405
r51 46 47 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r52 45 47 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r53 42 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.612 $Y2=0.234
r54 39 40 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.214
r55 38 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.203
r56 37 38 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.167
r57 36 37 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r58 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r59 34 35 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.097 $X2=0.621 $Y2=0.122
r60 33 34 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.621 $Y2=0.097
r61 32 45 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.234
r62 32 40 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.214
r63 31 33 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.09
r64 29 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.58
+ $Y=0.036 $X2=0.587 $Y2=0.036
r65 27 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.587 $Y2=0.036
r66 25 29 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.58 $Y2=0.036
r67 24 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r68 24 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.594 $Y2=0.036
r69 19 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.513 $Y=0.045 $X2=0.522 $Y2=0.036
r70 19 21 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.082
r71 17 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r72 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r73 12 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036 $X2=0.594
+ $Y2=0.036
r74 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.592 $Y2=0.0405
r75 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.082 $X2=0.513
+ $Y2=0.082
r76 5 7 552.609 $w=2e-08 $l=1.475e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.082 $X2=0.513 $Y2=0.2295
r77 2 5 155.48 $w=2e-08 $l=4.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.082
.ends

.subckt PM_DLLX2_ASAP7_75T_SRAM%8 2 5 7 10 15 18 21 23 25 30 33 37 38 41 46 47 48
+ 51 54 55 56 59 61 62 66 69 72 74 75 84 95 VSS
c68 97 VSS 4.52133e-19 $X=0.459 $Y=0.214
c69 96 VSS 5.73001e-20 $X=0.459 $Y=0.203
c70 95 VSS 2.69603e-19 $X=0.459 $Y=0.2
c71 84 VSS 0.00165093f $X=0.783 $Y=0.136
c72 75 VSS 0.00576591f $X=0.655 $Y=0.153
c73 74 VSS 0.00146501f $X=0.527 $Y=0.153
c74 72 VSS 0.00662989f $X=0.783 $Y=0.153
c75 69 VSS 3.75508e-19 $X=0.459 $Y=0.153
c76 66 VSS 3.21606e-19 $X=0.459 $Y=0.225
c77 65 VSS 2.32827e-19 $X=0.459 $Y=0.131
c78 62 VSS 3.60459e-20 $X=0.522 $Y=0.131
c79 61 VSS 0.00173419f $X=0.504 $Y=0.131
c80 59 VSS 0.00147804f $X=0.566 $Y=0.131
c81 56 VSS 3.61032e-19 $X=0.459 $Y=0.106
c82 55 VSS 2.74504e-19 $X=0.459 $Y=0.097
c83 54 VSS 1.75944e-19 $X=0.459 $Y=0.122
c84 51 VSS 0.00271748f $X=0.432 $Y=0.036
c85 48 VSS 0.00636101f $X=0.45 $Y=0.036
c86 47 VSS 0.00146362f $X=0.414 $Y=0.234
c87 46 VSS 0.00368178f $X=0.396 $Y=0.234
c88 41 VSS 0.00571919f $X=0.45 $Y=0.234
c89 40 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c90 37 VSS 0.00348747f $X=0.378 $Y=0.2025
c91 32 VSS 5.36734e-19 $X=0.432 $Y=0.0405
c92 21 VSS 0.0123567f $X=0.783 $Y=0.136
c93 18 VSS 0.0653215f $X=0.783 $Y=0.0675
c94 10 VSS 0.0660363f $X=0.729 $Y=0.0675
c95 5 VSS 0.00310914f $X=0.567 $Y=0.131
c96 2 VSS 0.0627936f $X=0.567 $Y=0.0405
r97 96 97 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.203 $X2=0.459 $Y2=0.214
r98 95 96 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.2 $X2=0.459 $Y2=0.203
r99 94 95 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.2
r100 74 75 8.69136 $w=1.8e-08 $l=1.28e-07 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.655 $Y2=0.153
r101 72 75 8.69136 $w=1.8e-08 $l=1.28e-07 $layer=M2 $thickness=3.6e-08 $X=0.783
+ $Y=0.153 $X2=0.655 $Y2=0.153
r102 72 84 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.783 $Y=0.153 $X2=0.783
+ $Y2=0.153
r103 69 94 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.459 $Y2=0.165
r104 68 74 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.527 $Y2=0.153
r105 68 69 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.459 $Y=0.153 $X2=0.459
+ $Y2=0.153
r106 66 97 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r107 64 69 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.153
r108 64 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r109 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r110 59 62 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.566
+ $Y=0.131 $X2=0.522 $Y2=0.131
r111 57 65 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r112 57 61 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.504 $Y2=0.131
r113 55 56 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.097 $X2=0.459 $Y2=0.106
r114 54 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r115 54 56 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.106
r116 53 55 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.097
r117 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r118 48 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r119 48 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.432 $Y2=0.036
r120 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r121 43 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r122 41 66 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r123 41 47 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.414 $Y2=0.234
r124 38 40 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r125 37 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r126 34 40 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r127 34 37 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r128 33 37 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r129 30 32 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r130 29 51 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r131 26 32 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r132 26 29 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r133 25 29 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r134 21 84 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.136 $X2=0.783
+ $Y2=0.136
r135 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.136 $X2=0.783 $Y2=0.2025
r136 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.136
r137 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.136 $X2=0.783 $Y2=0.136
r138 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.136 $X2=0.729 $Y2=0.2025
r139 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.136
r140 5 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.566 $Y=0.131 $X2=0.566
+ $Y2=0.131
r141 5 7 369.03 $w=2e-08 $l=9.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.131 $X2=0.567 $Y2=0.2295
r142 2 5 339.058 $w=2e-08 $l=9.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.131
.ends

.subckt PM_DLLX2_ASAP7_75T_SRAM%Q 1 6 11 14 16 24 28 29 30 39 40 44 46 VSS
c23 46 VSS 0.00354102f $X=0.838 $Y=0.167
c24 45 VSS 0.00221859f $X=0.838 $Y=0.09
c25 44 VSS 0.00284852f $X=0.84 $Y=0.223
c26 40 VSS 0.00146362f $X=0.792 $Y=0.234
c27 39 VSS 0.0108633f $X=0.774 $Y=0.234
c28 31 VSS 0.00721992f $X=0.829 $Y=0.234
c29 30 VSS 0.00146362f $X=0.792 $Y=0.036
c30 29 VSS 0.010874f $X=0.774 $Y=0.036
c31 28 VSS 0.0064856f $X=0.81 $Y=0.036
c32 24 VSS 0.00562335f $X=0.702 $Y=0.036
c33 21 VSS 0.00719871f $X=0.829 $Y=0.036
c34 19 VSS 0.00691357f $X=0.808 $Y=0.2025
c35 14 VSS 0.00572107f $X=0.704 $Y=0.2025
c36 11 VSS 3.4597e-19 $X=0.719 $Y=0.2025
c37 9 VSS 3.44349e-19 $X=0.808 $Y=0.0675
c38 1 VSS 3.44349e-19 $X=0.719 $Y=0.0675
r39 45 46 5.22839 $w=1.8e-08 $l=7.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.838
+ $Y=0.09 $X2=0.838 $Y2=0.167
r40 44 46 3.80247 $w=1.8e-08 $l=5.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.838
+ $Y=0.223 $X2=0.838 $Y2=0.167
r41 42 44 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.838
+ $Y=0.225 $X2=0.838 $Y2=0.223
r42 41 45 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.838
+ $Y=0.045 $X2=0.838 $Y2=0.09
r43 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.234 $X2=0.792 $Y2=0.234
r44 37 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.234 $X2=0.792 $Y2=0.234
r45 33 39 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.234 $X2=0.774 $Y2=0.234
r46 31 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.829 $Y=0.234 $X2=0.838 $Y2=0.225
r47 31 37 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.829
+ $Y=0.234 $X2=0.81 $Y2=0.234
r48 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.036 $X2=0.792 $Y2=0.036
r49 27 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.036 $X2=0.792 $Y2=0.036
r50 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.036 $X2=0.81
+ $Y2=0.036
r51 23 29 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.036 $X2=0.774 $Y2=0.036
r52 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.036 $X2=0.702
+ $Y2=0.036
r53 21 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.829 $Y=0.036 $X2=0.838 $Y2=0.045
r54 21 27 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.829
+ $Y=0.036 $X2=0.81 $Y2=0.036
r55 19 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.234 $X2=0.81
+ $Y2=0.234
r56 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2025 $X2=0.808 $Y2=0.2025
r57 14 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.234 $X2=0.702
+ $Y2=0.234
r58 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2025 $X2=0.704 $Y2=0.2025
r59 9 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.81
+ $Y=0.0675 $X2=0.81 $Y2=0.036
r60 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.793
+ $Y=0.0675 $X2=0.808 $Y2=0.0675
r61 4 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.702
+ $Y=0.0675 $X2=0.702 $Y2=0.036
r62 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.719
+ $Y=0.0675 $X2=0.704 $Y2=0.0675
.ends

.subckt PM_DLLX2_ASAP7_75T_SRAM%10 1 6 9 VSS
c7 9 VSS 0.0266424f $X=0.38 $Y=0.0675
c8 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c9 4 VSS 3.22674e-19 $X=0.322 $Y=0.0675
r10 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r12 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DLLX2_ASAP7_75T_SRAM%11 1 6 9 VSS
c9 9 VSS 0.0211025f $X=0.488 $Y=0.2295
c10 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c11 4 VSS 2.84146e-19 $X=0.43 $Y=0.2295
r12 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r13 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DLLX2_ASAP7_75T_SRAM%12 1 2 VSS
c0 1 VSS 0.00220425f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DLLX2_ASAP7_75T_SRAM%13 1 2 VSS
c1 1 VSS 0.00201018f $X=0.341 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends


* END of "./DLLx2_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DLLx2_ASAP7_75t_SRAM  VSS VDD CLK D Q
* 
* Q	Q
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_10_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_4_M3_g N_10_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_12_M4_d N_6_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_12_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 VSS N_8_M7_g N_Q_M7_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M8 VSS N_8_M8_g N_Q_M8_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773 $Y=0.027
M9 VDD N_CLK_M9_g N_4_M9_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M10 N_6_M10_d N_4_M10_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M11 N_13_M11_d N_D_M11_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M12 N_8_M12_d N_6_M12_g N_13_M12_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M13 N_11_M13_d N_4_M13_g N_8_M13_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M14 VDD N_7_M14_g N_11_M14_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M15 N_7_M15_d N_8_M15_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M16 VDD N_8_M16_g N_Q_M16_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M17 VDD N_8_M17_g N_Q_M17_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
*
* 
* .include "DLLx2_ASAP7_75t_SRAM.pex.sp.DLLX2_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DLLx2_ASAP7_75t_SRAM.pex.sp.DLLX2_ASAP7_75T_SRAM.pxi"
* File: DLLx2_ASAP7_75t_SRAM.pex.sp.DLLX2_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:28:38 2017
* 
x_PM_DLLX2_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_11_p N_CLK_M9_g CLK N_CLK_c_3_p
+ N_CLK_c_4_p VSS PM_DLLX2_ASAP7_75T_SRAM%CLK
x_PM_DLLX2_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M10_g N_4_M3_g N_4_c_38_p N_4_M13_g
+ N_4_M0_s N_4_c_20_n N_4_M9_s N_4_c_21_n N_4_c_22_n N_4_c_23_n N_4_c_24_n
+ N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_48_p N_4_c_28_n N_4_c_29_n N_4_c_30_n
+ N_4_c_31_n N_4_c_53_p N_4_c_32_n N_4_c_36_p N_4_c_40_p VSS
+ PM_DLLX2_ASAP7_75T_SRAM%4
x_PM_DLLX2_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_64_n N_D_M11_g D N_D_c_69_p VSS
+ PM_DLLX2_ASAP7_75T_SRAM%D
x_PM_DLLX2_ASAP7_75T_SRAM%6 N_6_c_87_n N_6_M12_g N_6_M4_g N_6_c_90_n N_6_M1_d
+ N_6_M10_d N_6_c_91_n N_6_c_92_n N_6_c_84_n N_6_c_94_n N_6_c_95_n N_6_c_85_n
+ N_6_c_97_n N_6_c_109_n N_6_c_98_n N_6_c_111_n N_6_c_142_p N_6_c_100_n
+ N_6_c_132_p N_6_c_103_n N_6_c_119_p N_6_c_120_p N_6_c_86_n N_6_c_116_n
+ N_6_c_117_n VSS PM_DLLX2_ASAP7_75T_SRAM%6
x_PM_DLLX2_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_162_n N_7_M14_g N_7_M6_d N_7_c_163_n
+ N_7_M15_d N_7_c_164_n N_7_c_173_p N_7_c_187_p N_7_c_172_p N_7_c_170_p
+ N_7_c_186_p N_7_c_182_p N_7_c_174_p N_7_c_171_p N_7_c_180_p N_7_c_165_n
+ N_7_c_167_n N_7_c_188_p N_7_c_168_n VSS PM_DLLX2_ASAP7_75T_SRAM%7
x_PM_DLLX2_ASAP7_75T_SRAM%8 N_8_M6_g N_8_c_222_n N_8_M15_g N_8_M7_g N_8_M16_g
+ N_8_M8_g N_8_c_238_p N_8_M17_g N_8_M3_d N_8_M4_s N_8_M12_d N_8_c_189_n
+ N_8_M13_s N_8_c_202_n N_8_c_196_n N_8_c_190_n N_8_c_197_n N_8_c_205_n
+ N_8_c_192_n N_8_c_207_n N_8_c_225_n N_8_c_208_n N_8_c_209_n N_8_c_210_n
+ N_8_c_256_p N_8_c_193_n N_8_c_234_p N_8_c_194_n N_8_c_230_n N_8_c_233_n
+ N_8_c_216_n VSS PM_DLLX2_ASAP7_75T_SRAM%8
x_PM_DLLX2_ASAP7_75T_SRAM%Q N_Q_M7_s N_Q_M8_s N_Q_M16_s N_Q_c_257_n N_Q_M17_s
+ N_Q_c_260_n N_Q_c_266_n N_Q_c_262_n N_Q_c_270_n N_Q_c_263_n N_Q_c_275_n Q
+ N_Q_c_277_n VSS PM_DLLX2_ASAP7_75T_SRAM%Q
x_PM_DLLX2_ASAP7_75T_SRAM%10 N_10_M2_d N_10_M3_s N_10_c_280_n VSS
+ PM_DLLX2_ASAP7_75T_SRAM%10
x_PM_DLLX2_ASAP7_75T_SRAM%11 N_11_M13_d N_11_M14_s N_11_c_288_n VSS
+ PM_DLLX2_ASAP7_75T_SRAM%11
x_PM_DLLX2_ASAP7_75T_SRAM%12 N_12_M5_s N_12_M4_d VSS PM_DLLX2_ASAP7_75T_SRAM%12
x_PM_DLLX2_ASAP7_75T_SRAM%13 N_13_M12_s N_13_M11_d VSS PM_DLLX2_ASAP7_75T_SRAM%13
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_20_n 2.66516e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 N_CLK_c_3_p N_4_c_21_n 2.66516e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.216
cc_4 N_CLK_c_4_p N_4_c_22_n 0.00126555f $X=0.081 $Y=0.1305 $X2=0.018 $Y2=0.144
cc_5 CLK N_4_c_23_n 3.98992e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.081
cc_6 CLK N_4_c_24_n 0.00126555f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.1125
cc_7 N_CLK_c_3_p N_4_c_25_n 0.00127356f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.189
cc_8 CLK N_4_c_26_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_3_p N_4_c_27_n 4.98319e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_4_p N_4_c_28_n 4.17e-19 $X=0.081 $Y=0.1305 $X2=0.152 $Y2=0.135
cc_11 N_CLK_c_11_p N_4_c_29_n 0.00116357f $X=0.081 $Y=0.135 $X2=0.152 $Y2=0.135
cc_12 N_CLK_c_3_p N_4_c_30_n 0.00122788f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.153
cc_13 N_CLK_c_3_p N_4_c_31_n 0.00197837f $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.153
cc_14 CLK N_4_c_32_n 5.08945e-19 $X=0.082 $Y=0.119 $X2=0.229 $Y2=0.153
cc_15 N_CLK_c_3_p N_4_c_32_n 0.00150524f $X=0.081 $Y=0.135 $X2=0.229 $Y2=0.153
cc_16 CLK N_6_c_84_n 6.45949e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.189
cc_17 N_CLK_c_3_p N_6_c_85_n 6.45949e-19 $X=0.081 $Y=0.135 $X2=0.0505 $Y2=0.036
cc_18 CLK N_6_c_86_n 7.98675e-19 $X=0.082 $Y=0.119 $X2=0.152 $Y2=0.135
cc_19 N_4_M3_g N_D_M2_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_20 N_4_c_29_n N_D_c_64_n 2.01856e-19 $X=0.152 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 N_4_c_36_p D 0.00117371f $X=0.317 $Y=0.153 $X2=0.082 $Y2=0.119
cc_22 N_4_M3_g N_6_c_87_n 0.00355599f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_23 N_4_c_38_p N_6_c_87_n 0.00101396f $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.054
cc_24 N_4_M3_g N_6_M4_g 0.00355599f $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_25 N_4_c_40_p N_6_c_90_n 3.2936e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.126
cc_26 N_4_c_31_n N_6_c_91_n 0.00243501f $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_27 N_4_c_36_p N_6_c_92_n 2.3925e-19 $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_28 N_4_c_28_n N_6_c_84_n 9.58415e-19 $X=0.152 $Y=0.135 $X2=0 $Y2=0
cc_29 N_4_c_32_n N_6_c_94_n 2.3925e-19 $X=0.229 $Y=0.153 $X2=0 $Y2=0
cc_30 N_4_c_36_p N_6_c_95_n 2.75285e-19 $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_31 N_4_c_31_n N_6_c_85_n 0.00467935f $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_32 N_4_c_32_n N_6_c_97_n 2.75285e-19 $X=0.229 $Y=0.153 $X2=0 $Y2=0
cc_33 N_4_c_48_p N_6_c_98_n 0.00396181f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_34 N_4_c_36_p N_6_c_98_n 0.00119509f $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_35 N_4_c_31_n N_6_c_100_n 3.89771e-19 $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_36 N_4_c_36_p N_6_c_100_n 0.0160263f $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_37 N_4_c_40_p N_6_c_100_n 8.49272e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_53_p N_6_c_103_n 0.00115166f $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_40_p N_6_c_103_n 0.00433569f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_41 N_4_c_40_p N_8_c_189_n 0.00195725f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_42 N_4_M3_g N_8_c_190_n 2.63086e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_4_c_40_p N_8_c_190_n 0.00122664f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_44 N_4_c_40_p N_8_c_192_n 0.00419136f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_45 N_4_c_40_p N_8_c_193_n 2.60642e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_53_p N_8_c_194_n 9.23088e-19 $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_36_p N_10_c_280_n 8.32437e-19 $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_48 N_D_M2_g N_6_c_87_n 0.00341068f $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_49 N_D_c_64_n N_6_c_87_n 0.00101372f $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_50 D N_6_c_92_n 0.00115278f $X=0.297 $Y=0.1165 $X2=0.018 $Y2=0.144
cc_51 N_D_c_69_p N_6_c_95_n 0.00115278f $X=0.297 $Y=0.135 $X2=0.027 $Y2=0.036
cc_52 N_D_c_69_p N_6_c_109_n 0.00115278f $X=0.297 $Y=0.135 $X2=0.054 $Y2=0.234
cc_53 D N_6_c_98_n 0.00124619f $X=0.297 $Y=0.1165 $X2=0.047 $Y2=0.234
cc_54 D N_6_c_111_n 0.00216863f $X=0.297 $Y=0.1165 $X2=0.152 $Y2=0.135
cc_55 D N_6_c_100_n 8.86605e-19 $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_56 N_D_c_69_p N_6_c_100_n 3.97512e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_57 D N_6_c_103_n 0.00216863f $X=0.297 $Y=0.1165 $X2=0.189 $Y2=0.144
cc_58 D N_6_c_86_n 0.00115278f $X=0.297 $Y=0.1165 $X2=0.152 $Y2=0.135
cc_59 D N_6_c_116_n 0.00115278f $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_60 N_D_c_69_p N_6_c_117_n 0.00115278f $X=0.297 $Y=0.135 $X2=0.405 $Y2=0.135
cc_61 N_D_c_69_p N_8_c_189_n 3.88702e-19 $X=0.297 $Y=0.135 $X2=0.054 $Y2=0.036
cc_62 N_D_c_69_p N_8_c_196_n 8.77202e-19 $X=0.297 $Y=0.135 $X2=0.047 $Y2=0.234
cc_63 D N_8_c_197_n 2.05539e-19 $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_64 D N_10_c_280_n 0.00428733f $X=0.297 $Y=0.1165 $X2=0.405 $Y2=0.0675
cc_65 N_D_c_69_p N_13_M12_s 3.05674e-19 $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_66 N_6_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_67 N_6_c_119_p N_7_M5_g 0.00199227f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_68 N_6_c_120_p N_7_M5_g 4.91626e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_69 N_6_c_119_p N_7_c_162_n 4.44368e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.135
cc_70 N_6_c_119_p N_7_c_163_n 5.31675e-19 $X=0.513 $Y=0.18 $X2=0.082 $Y2=0.119
cc_71 N_6_c_119_p N_7_c_164_n 0.00169036f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.1305
cc_72 N_6_c_119_p N_7_c_165_n 6.34096e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_73 N_6_c_120_p N_7_c_165_n 5.95005e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_74 N_6_c_119_p N_7_c_167_n 0.00267575f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_75 N_6_c_119_p N_7_c_168_n 5.97916e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_76 N_6_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_77 N_6_c_119_p N_8_M6_g 0.00305655f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_78 N_6_c_100_n N_8_c_189_n 2.84357e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_79 N_6_c_103_n N_8_c_189_n 0.00130164f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_80 N_6_c_132_p N_8_c_202_n 7.16323e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_81 N_6_c_100_n N_8_c_196_n 5.53186e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_82 N_6_c_132_p N_8_c_197_n 3.48842e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_83 N_6_c_132_p N_8_c_205_n 2.01793e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_84 N_6_M4_g N_8_c_192_n 2.93184e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_85 N_6_M4_g N_8_c_207_n 3.72919e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_86 N_6_c_119_p N_8_c_208_n 4.41338e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_87 N_6_c_119_p N_8_c_209_n 7.92645e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_88 N_6_c_120_p N_8_c_210_n 0.00100546f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_89 N_6_M4_g N_8_c_193_n 2.27241e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_90 N_6_c_142_p N_8_c_193_n 2.46239e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_91 N_6_c_142_p N_8_c_194_n 0.00694438f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_92 N_6_c_119_p N_8_c_194_n 0.00195448f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_93 N_6_c_120_p N_8_c_194_n 2.84312e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_94 N_6_c_90_n N_8_c_216_n 0.00271026f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_95 N_6_c_142_p N_8_c_216_n 6.73646e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_96 N_6_c_119_p N_8_c_216_n 5.95032e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_97 N_6_c_120_p N_8_c_216_n 0.00182777f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_98 N_6_c_119_p N_Q_c_257_n 0.00114499f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.135
cc_99 N_6_c_87_n N_10_c_280_n 0.00639848f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_100 N_6_c_103_n N_10_c_280_n 0.00135407f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_101 N_6_c_119_p N_11_M14_s 2.34172e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.216
cc_102 N_6_M4_g N_11_c_288_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_103 N_6_c_90_n N_11_c_288_n 0.0013957f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_104 N_6_c_132_p N_11_c_288_n 7.09553e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_105 N_6_c_119_p N_11_c_288_n 0.00230185f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_106 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_107 N_7_c_170_p N_8_M6_g 4.17397e-19 $X=0.58 $Y=0.036 $X2=0.135 $Y2=0.054
cc_108 N_7_c_171_p N_8_c_222_n 3.48572e-19 $X=0.621 $Y=0.14 $X2=0.135 $Y2=0.135
cc_109 N_7_c_172_p N_8_c_197_n 0.00177955f $X=0.522 $Y=0.036 $X2=0 $Y2=0
cc_110 N_7_c_173_p N_8_c_207_n 0.00177955f $X=0.513 $Y=0.082 $X2=0 $Y2=0
cc_111 N_7_c_174_p N_8_c_225_n 2.8599e-19 $X=0.621 $Y=0.122 $X2=0 $Y2=0
cc_112 N_7_c_170_p N_8_c_208_n 6.9494e-19 $X=0.58 $Y=0.036 $X2=0.189 $Y2=0.144
cc_113 N_7_c_171_p N_8_c_208_n 9.49516e-19 $X=0.621 $Y=0.14 $X2=0.189 $Y2=0.144
cc_114 N_7_M5_g N_8_c_210_n 4.06683e-19 $X=0.513 $Y=0.0405 $X2=0.033 $Y2=0.153
cc_115 N_7_c_173_p N_8_c_210_n 0.00116089f $X=0.513 $Y=0.082 $X2=0.033 $Y2=0.153
cc_116 N_7_c_163_n N_8_c_230_n 2.11538e-19 $X=0.592 $Y=0.0405 $X2=0.152
+ $Y2=0.135
cc_117 N_7_c_180_p N_8_c_230_n 0.00133609f $X=0.621 $Y=0.165 $X2=0.152 $Y2=0.135
cc_118 N_7_c_168_n N_8_c_230_n 5.94743e-19 $X=0.612 $Y=0.234 $X2=0.152 $Y2=0.135
cc_119 N_7_c_182_p N_8_c_233_n 4.47522e-19 $X=0.621 $Y=0.097 $X2=0 $Y2=0
cc_120 N_7_c_164_n N_Q_c_257_n 4.7734e-19 $X=0.592 $Y=0.2295 $X2=0.405
+ $Y2=0.2295
cc_121 N_7_c_167_n N_Q_c_257_n 7.18237e-19 $X=0.621 $Y=0.203 $X2=0.405
+ $Y2=0.2295
cc_122 N_7_c_163_n N_Q_c_260_n 4.7734e-19 $X=0.592 $Y=0.0405 $X2=0 $Y2=0
cc_123 N_7_c_186_p N_Q_c_260_n 0.00151703f $X=0.621 $Y=0.09 $X2=0 $Y2=0
cc_124 N_7_c_187_p N_Q_c_262_n 8.34906e-19 $X=0.612 $Y=0.036 $X2=0.018 $Y2=0.081
cc_125 N_7_c_188_p N_Q_c_263_n 7.82687e-19 $X=0.621 $Y=0.234 $X2=0.047 $Y2=0.036
cc_126 N_8_c_234_p N_Q_c_257_n 3.0124e-19 $X=0.783 $Y=0.153 $X2=0.405 $Y2=0.2295
cc_127 N_8_c_234_p N_Q_c_260_n 2.54113e-19 $X=0.783 $Y=0.153 $X2=0 $Y2=0
cc_128 N_8_c_233_n N_Q_c_266_n 5.47049e-19 $X=0.783 $Y=0.136 $X2=0.018 $Y2=0.144
cc_129 N_8_M7_g N_Q_c_262_n 4.61817e-19 $X=0.729 $Y=0.0675 $X2=0.018 $Y2=0.081
cc_130 N_8_c_238_p N_Q_c_262_n 7.47725e-19 $X=0.783 $Y=0.136 $X2=0.018 $Y2=0.081
cc_131 N_8_c_234_p N_Q_c_262_n 8.84447e-19 $X=0.783 $Y=0.153 $X2=0.018 $Y2=0.081
cc_132 N_8_M8_g N_Q_c_270_n 3.24181e-19 $X=0.783 $Y=0.0675 $X2=0.018 $Y2=0.1125
cc_133 N_8_c_233_n N_Q_c_270_n 7.27236e-19 $X=0.783 $Y=0.136 $X2=0.018
+ $Y2=0.1125
cc_134 N_8_M7_g N_Q_c_263_n 4.56556e-19 $X=0.729 $Y=0.0675 $X2=0.047 $Y2=0.036
cc_135 N_8_c_238_p N_Q_c_263_n 4.51177e-19 $X=0.783 $Y=0.136 $X2=0.047 $Y2=0.036
cc_136 N_8_c_234_p N_Q_c_263_n 0.00108469f $X=0.783 $Y=0.153 $X2=0.047 $Y2=0.036
cc_137 N_8_M8_g N_Q_c_275_n 3.50534e-19 $X=0.783 $Y=0.0675 $X2=0.0505 $Y2=0.036
cc_138 N_8_c_233_n N_Q_c_275_n 5.44675e-19 $X=0.783 $Y=0.136 $X2=0.0505
+ $Y2=0.036
cc_139 N_8_c_238_p N_Q_c_277_n 3.48717e-19 $X=0.783 $Y=0.136 $X2=0.047 $Y2=0.234
cc_140 N_8_c_234_p N_Q_c_277_n 2.37083e-19 $X=0.783 $Y=0.153 $X2=0.047 $Y2=0.234
cc_141 N_8_c_233_n N_Q_c_277_n 0.00321733f $X=0.783 $Y=0.136 $X2=0.047 $Y2=0.234
cc_142 N_8_c_189_n N_10_c_280_n 0.00119636f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_143 N_8_c_197_n N_10_c_280_n 4.50844e-19 $X=0.45 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_144 N_8_c_205_n N_10_c_280_n 0.00394776f $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_145 N_8_c_189_n N_11_c_288_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_146 N_8_c_202_n N_11_c_288_n 0.00343017f $X=0.45 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_147 N_8_c_205_n N_11_c_288_n 5.72355e-19 $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_148 N_8_c_256_p N_11_c_288_n 0.00116187f $X=0.459 $Y=0.225 $X2=0.405
+ $Y2=0.0675

* END of "./DLLx2_ASAP7_75t_SRAM.pex.sp.DLLX2_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: DLLx3_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:29:00 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "DLLx3_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./DLLx3_ASAP7_75t_SRAM.pex.sp.pex"
* File: DLLx3_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:29:00 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_DLLX3_ASAP7_75T_SRAM%CLK 2 5 7 12 14 17 VSS
c18 17 VSS 5.41721e-21 $X=0.081 $Y=0.1305
c19 14 VSS 0.00732563f $X=0.081 $Y=0.135
c20 12 VSS 0.00698013f $X=0.082 $Y=0.119
c21 5 VSS 0.0020626f $X=0.081 $Y=0.135
c22 2 VSS 0.062963f $X=0.081 $Y=0.054
r23 16 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r24 14 17 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r25 12 16 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.119 $X2=0.081 $Y2=0.126
r26 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r28 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_DLLX3_ASAP7_75T_SRAM%4 2 7 10 13 15 17 20 22 25 28 29 30 33 37 44 49 51
+ 52 62 66 68 70 71 79 VSS
c44 96 VSS 1.06551e-19 $X=0.03 $Y=0.153
c45 95 VSS 6.89947e-19 $X=0.027 $Y=0.153
c46 79 VSS 0.00117246f $X=0.405 $Y=0.135
c47 71 VSS 0.0029117f $X=0.317 $Y=0.153
c48 70 VSS 0.00767547f $X=0.229 $Y=0.153
c49 68 VSS 0.00297348f $X=0.405 $Y=0.153
c50 66 VSS 0.00148441f $X=0.189 $Y=0.153
c51 62 VSS 9.21052e-19 $X=0.033 $Y=0.153
c52 52 VSS 0.00385436f $X=0.152 $Y=0.135
c53 51 VSS 4.1341e-19 $X=0.152 $Y=0.135
c54 49 VSS 0.00125241f $X=0.18 $Y=0.135
c55 47 VSS 3.02772e-19 $X=0.0505 $Y=0.234
c56 46 VSS 0.00180216f $X=0.047 $Y=0.234
c57 44 VSS 0.00250477f $X=0.054 $Y=0.234
c58 42 VSS 0.00305101f $X=0.027 $Y=0.234
c59 40 VSS 3.02772e-19 $X=0.0505 $Y=0.036
c60 39 VSS 0.00199699f $X=0.047 $Y=0.036
c61 37 VSS 0.00250477f $X=0.054 $Y=0.036
c62 35 VSS 0.00305101f $X=0.027 $Y=0.036
c63 34 VSS 9.44133e-19 $X=0.018 $Y=0.207
c64 33 VSS 0.00134027f $X=0.018 $Y=0.189
c65 32 VSS 8.82937e-19 $X=0.018 $Y=0.225
c66 30 VSS 0.00159315f $X=0.018 $Y=0.1125
c67 29 VSS 0.00142827f $X=0.018 $Y=0.081
c68 28 VSS 0.00144655f $X=0.018 $Y=0.144
c69 25 VSS 0.00453739f $X=0.056 $Y=0.216
c70 22 VSS 2.98509e-19 $X=0.071 $Y=0.216
c71 20 VSS 0.00456252f $X=0.056 $Y=0.054
c72 17 VSS 2.98509e-19 $X=0.071 $Y=0.054
c73 13 VSS 0.0015517f $X=0.405 $Y=0.135
c74 10 VSS 0.059003f $X=0.405 $Y=0.0675
c75 2 VSS 0.0627154f $X=0.135 $Y=0.054
r76 95 96 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.153 $X2=0.03 $Y2=0.153
r77 92 95 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.153 $X2=0.027 $Y2=0.153
r78 70 71 5.97531 $w=1.8e-08 $l=8.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.153 $X2=0.317 $Y2=0.153
r79 68 71 5.97531 $w=1.8e-08 $l=8.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.317 $Y2=0.153
r80 68 79 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.405 $Y=0.153 $X2=0.405
+ $Y2=0.153
r81 65 70 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.189
+ $Y=0.153 $X2=0.229 $Y2=0.153
r82 65 66 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.189 $Y=0.153 $X2=0.189
+ $Y2=0.153
r83 62 96 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.03 $Y2=0.153
r84 61 65 10.5926 $w=1.8e-08 $l=1.56e-07 $layer=M2 $thickness=3.6e-08 $X=0.033
+ $Y=0.153 $X2=0.189 $Y2=0.153
r85 61 62 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.033 $Y=0.153 $X2=0.033
+ $Y2=0.153
r86 59 66 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.153
r87 51 52 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.152 $Y=0.135 $X2=0.152
+ $Y2=0.135
r88 49 59 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r89 49 51 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.152 $Y2=0.135
r90 46 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r91 44 47 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0505 $Y2=0.234
r92 42 46 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.047 $Y2=0.234
r93 39 40 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r94 37 40 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0505 $Y2=0.036
r95 35 39 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.047 $Y2=0.036
r96 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.207
r97 32 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r98 32 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.207
r99 31 92 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.153
r100 31 33 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.162 $X2=0.018 $Y2=0.189
r101 29 30 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.1125
r102 28 92 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.153
r103 28 30 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1125
r104 27 35 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r105 27 29 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.081
r106 25 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r107 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r108 20 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r109 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r110 13 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r111 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2295
r112 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r113 5 52 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.152 $Y2=0.135
r114 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r115 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_DLLX3_ASAP7_75T_SRAM%D 2 5 7 12 16 VSS
c21 16 VSS 0.00596102f $X=0.297 $Y=0.135
c22 12 VSS 0.00848689f $X=0.297 $Y=0.1165
c23 5 VSS 0.0019062f $X=0.297 $Y=0.135
c24 2 VSS 0.061556f $X=0.297 $Y=0.0675
r25 12 16 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1165 $X2=0.297 $Y2=0.135
r26 5 16 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r27 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r28 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_DLLX3_ASAP7_75T_SRAM%6 2 5 8 16 18 23 26 28 33 34 35 40 41 43 46 50 52
+ 54 55 59 71 72 75 76 78 VSS
c72 78 VSS 3.82279e-19 $X=0.243 $Y=0.216
c73 76 VSS 4.13588e-19 $X=0.243 $Y=0.126
c74 75 VSS 0.00265408f $X=0.243 $Y=0.117
c75 72 VSS 6.21924e-19 $X=0.513 $Y=0.18
c76 71 VSS 0.0601566f $X=0.513 $Y=0.18
c77 59 VSS 8.58425e-19 $X=0.351 $Y=0.135
c78 55 VSS 0.00132732f $X=0.45 $Y=0.189
c79 54 VSS 0.0053562f $X=0.414 $Y=0.189
c80 52 VSS 0.00304981f $X=0.513 $Y=0.189
c81 50 VSS 6.50668e-19 $X=0.351 $Y=0.189
c82 46 VSS 0.00221329f $X=0.243 $Y=0.189
c83 43 VSS 3.61041e-19 $X=0.243 $Y=0.225
c84 41 VSS 0.0018377f $X=0.216 $Y=0.234
c85 40 VSS 0.0051665f $X=0.198 $Y=0.234
c86 35 VSS 0.00483896f $X=0.234 $Y=0.234
c87 34 VSS 0.00184198f $X=0.216 $Y=0.036
c88 33 VSS 0.00552625f $X=0.198 $Y=0.036
c89 28 VSS 0.00484739f $X=0.234 $Y=0.036
c90 26 VSS 0.00641989f $X=0.16 $Y=0.216
c91 21 VSS 0.00625354f $X=0.16 $Y=0.054
c92 16 VSS 0.00212305f $X=0.464 $Y=0.179
c93 8 VSS 0.059718f $X=0.459 $Y=0.0405
c94 2 VSS 0.060362f $X=0.351 $Y=0.135
r95 77 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.207 $X2=0.243 $Y2=0.216
r96 75 76 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.117 $X2=0.243 $Y2=0.126
r97 71 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.513 $Y=0.18 $X2=0.513
+ $Y2=0.18
r98 54 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.414
+ $Y=0.189 $X2=0.45 $Y2=0.189
r99 52 55 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.45 $Y2=0.189
r100 52 72 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r101 50 59 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.135
r102 49 54 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.414 $Y2=0.189
r103 49 50 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.351 $Y=0.189 $X2=0.351
+ $Y2=0.189
r104 46 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.207
r105 46 76 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.243 $Y2=0.126
r106 45 49 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.189 $X2=0.351 $Y2=0.189
r107 45 46 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.189 $X2=0.243
+ $Y2=0.189
r108 43 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.216
r109 42 75 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.117
r110 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.216 $Y2=0.234
r111 37 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.198 $Y2=0.234
r112 35 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r113 35 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r114 33 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.216 $Y2=0.036
r115 30 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r116 28 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r117 28 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r118 26 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r119 23 26 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.16 $Y2=0.216
r120 21 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r121 18 21 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.16 $Y2=0.054
r122 16 71 42.2917 $w=2.4e-08 $l=4.9e-08 $layer=LISD $thickness=2.8e-08 $X=0.464
+ $Y=0.179 $X2=0.513 $Y2=0.179
r123 11 16 3.57143 $w=2.8e-08 $l=5e-09 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.179 $X2=0.464 $Y2=0.179
r124 8 11 518.891 $w=2e-08 $l=1.385e-07 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0405 $X2=0.459 $Y2=0.179
r125 2 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r126 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
.ends

.subckt PM_DLLX3_ASAP7_75T_SRAM%7 2 5 7 9 12 14 17 21 25 29 35 36 37 38 39 40 48
+ VSS
c24 48 VSS 0.00411848f $X=0.612 $Y=0.234
c25 47 VSS 0.00242619f $X=0.621 $Y=0.234
c26 42 VSS 3.89262e-19 $X=0.621 $Y=0.2205
c27 41 VSS 6.05812e-19 $X=0.621 $Y=0.216
c28 40 VSS 0.00109986f $X=0.621 $Y=0.203
c29 39 VSS 4.0755e-20 $X=0.621 $Y=0.167
c30 38 VSS 7.68431e-19 $X=0.621 $Y=0.165
c31 37 VSS 5.4967e-19 $X=0.621 $Y=0.14
c32 36 VSS 0.0011376f $X=0.621 $Y=0.122
c33 35 VSS 2.45537e-19 $X=0.621 $Y=0.097
c34 34 VSS 0.00138875f $X=0.621 $Y=0.09
c35 33 VSS 2.06522e-19 $X=0.621 $Y=0.054
c36 32 VSS 4.87917e-19 $X=0.621 $Y=0.225
c37 30 VSS 8.17537e-19 $X=0.587 $Y=0.036
c38 29 VSS 0.00649884f $X=0.58 $Y=0.036
c39 25 VSS 0.0022245f $X=0.522 $Y=0.036
c40 24 VSS 0.00518075f $X=0.612 $Y=0.036
c41 21 VSS 5.81526e-19 $X=0.513 $Y=0.082
c42 17 VSS 0.00494953f $X=0.592 $Y=0.2295
c43 12 VSS 0.00511578f $X=0.592 $Y=0.0405
c44 5 VSS 0.00256679f $X=0.513 $Y=0.082
c45 2 VSS 0.0581876f $X=0.513 $Y=0.0405
r46 48 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r47 47 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.234 $X2=0.6165 $Y2=0.234
r48 44 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.612 $Y2=0.234
r49 41 42 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.216 $X2=0.621 $Y2=0.2205
r50 40 41 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.203 $X2=0.621 $Y2=0.216
r51 39 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.167 $X2=0.621 $Y2=0.203
r52 38 39 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.165 $X2=0.621 $Y2=0.167
r53 37 38 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.14 $X2=0.621 $Y2=0.165
r54 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.122 $X2=0.621 $Y2=0.14
r55 35 36 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.097 $X2=0.621 $Y2=0.122
r56 34 35 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.09 $X2=0.621 $Y2=0.097
r57 33 34 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.054 $X2=0.621 $Y2=0.09
r58 32 47 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.234
r59 32 42 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.2205
r60 31 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.054
r61 29 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.58
+ $Y=0.036 $X2=0.587 $Y2=0.036
r62 27 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.587 $Y2=0.036
r63 25 29 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.58 $Y2=0.036
r64 24 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r65 24 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.594 $Y2=0.036
r66 19 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.513 $Y=0.045 $X2=0.522 $Y2=0.036
r67 19 21 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.082
r68 17 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r69 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2295 $X2=0.592 $Y2=0.2295
r70 12 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036 $X2=0.594
+ $Y2=0.036
r71 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0405 $X2=0.592 $Y2=0.0405
r72 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.082 $X2=0.513
+ $Y2=0.082
r73 5 7 552.609 $w=2e-08 $l=1.475e-07 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.082 $X2=0.513 $Y2=0.2295
r74 2 5 155.48 $w=2e-08 $l=4.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0405 $X2=0.513 $Y2=0.082
.ends

.subckt PM_DLLX3_ASAP7_75T_SRAM%8 2 5 7 10 15 18 23 26 29 31 33 38 41 45 46 49 54
+ 55 56 59 62 63 64 67 69 70 74 77 80 82 83 92 104 VSS
c71 106 VSS 4.52211e-19 $X=0.459 $Y=0.214
c72 105 VSS 5.73001e-20 $X=0.459 $Y=0.203
c73 104 VSS 2.69603e-19 $X=0.459 $Y=0.2
c74 92 VSS 0.00162514f $X=0.783 $Y=0.136
c75 83 VSS 0.00576591f $X=0.655 $Y=0.153
c76 82 VSS 0.00146501f $X=0.527 $Y=0.153
c77 80 VSS 0.00900516f $X=0.783 $Y=0.153
c78 77 VSS 3.75585e-19 $X=0.459 $Y=0.153
c79 74 VSS 3.21683e-19 $X=0.459 $Y=0.225
c80 73 VSS 2.32827e-19 $X=0.459 $Y=0.131
c81 70 VSS 3.60459e-20 $X=0.522 $Y=0.131
c82 69 VSS 0.00173419f $X=0.504 $Y=0.131
c83 67 VSS 0.00147804f $X=0.566 $Y=0.131
c84 64 VSS 3.61032e-19 $X=0.459 $Y=0.106
c85 63 VSS 2.74504e-19 $X=0.459 $Y=0.097
c86 62 VSS 1.75944e-19 $X=0.459 $Y=0.122
c87 59 VSS 0.00271748f $X=0.432 $Y=0.036
c88 56 VSS 0.00636101f $X=0.45 $Y=0.036
c89 55 VSS 0.00146362f $X=0.414 $Y=0.234
c90 54 VSS 0.00368178f $X=0.396 $Y=0.234
c91 49 VSS 0.00571919f $X=0.45 $Y=0.234
c92 48 VSS 5.70081e-19 $X=0.378 $Y=0.2295
c93 45 VSS 0.00348747f $X=0.378 $Y=0.2025
c94 40 VSS 5.36734e-19 $X=0.432 $Y=0.0405
c95 29 VSS 0.0142079f $X=0.837 $Y=0.136
c96 26 VSS 0.0648808f $X=0.837 $Y=0.0675
c97 18 VSS 0.0609677f $X=0.783 $Y=0.0675
c98 10 VSS 0.0625545f $X=0.729 $Y=0.0675
c99 5 VSS 0.0031159f $X=0.567 $Y=0.131
c100 2 VSS 0.0616253f $X=0.567 $Y=0.0405
r101 105 106 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.459 $Y=0.203 $X2=0.459 $Y2=0.214
r102 104 105 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.2 $X2=0.459 $Y2=0.203
r103 103 104 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.165 $X2=0.459 $Y2=0.2
r104 82 83 8.69136 $w=1.8e-08 $l=1.28e-07 $layer=M2 $thickness=3.6e-08 $X=0.527
+ $Y=0.153 $X2=0.655 $Y2=0.153
r105 80 83 8.69136 $w=1.8e-08 $l=1.28e-07 $layer=M2 $thickness=3.6e-08 $X=0.783
+ $Y=0.153 $X2=0.655 $Y2=0.153
r106 80 92 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.783 $Y=0.153 $X2=0.783
+ $Y2=0.153
r107 77 103 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.459 $Y2=0.165
r108 76 82 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.527 $Y2=0.153
r109 76 77 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.459 $Y=0.153 $X2=0.459
+ $Y2=0.153
r110 74 106 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.214
r111 72 77 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.153
r112 72 73 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.14 $X2=0.459 $Y2=0.131
r113 69 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.131 $X2=0.522 $Y2=0.131
r114 67 70 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.566
+ $Y=0.131 $X2=0.522 $Y2=0.131
r115 65 73 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.459 $Y2=0.131
r116 65 69 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.131 $X2=0.504 $Y2=0.131
r117 63 64 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.097 $X2=0.459 $Y2=0.106
r118 62 73 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.131
r119 62 64 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.122 $X2=0.459 $Y2=0.106
r120 61 63 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.097
r121 58 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r122 56 61 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r123 56 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.432 $Y2=0.036
r124 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.414 $Y2=0.234
r125 51 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r126 49 74 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r127 49 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.414 $Y2=0.234
r128 46 48 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2295 $X2=0.378 $Y2=0.2295
r129 45 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r130 42 48 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.378 $Y2=0.2295
r131 42 45 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.3735 $Y=0.216 $X2=0.3735 $Y2=0.189
r132 41 45 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.189 $X2=0.3735 $Y2=0.189
r133 38 40 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0405 $X2=0.432 $Y2=0.0405
r134 37 59 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r135 34 40 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.432 $Y2=0.0405
r136 34 37 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.4275 $Y=0.054 $X2=0.4275 $Y2=0.081
r137 33 37 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.081 $X2=0.4275 $Y2=0.081
r138 29 31 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.136 $X2=0.837 $Y2=0.2025
r139 26 29 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0675 $X2=0.837 $Y2=0.136
r140 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.783
+ $Y=0.136 $X2=0.837 $Y2=0.136
r141 21 92 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.783 $Y=0.136 $X2=0.783
+ $Y2=0.136
r142 21 23 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.136 $X2=0.783 $Y2=0.2025
r143 18 21 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.136
r144 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.136 $X2=0.783 $Y2=0.136
r145 13 15 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.136 $X2=0.729 $Y2=0.2025
r146 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.136
r147 5 67 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.566 $Y=0.131 $X2=0.566
+ $Y2=0.131
r148 5 7 369.03 $w=2e-08 $l=9.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.131 $X2=0.567 $Y2=0.2295
r149 2 5 339.058 $w=2e-08 $l=9.05e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0405 $X2=0.567 $Y2=0.131
.ends

.subckt PM_DLLX3_ASAP7_75T_SRAM%Q 1 2 6 11 12 15 16 21 24 29 30 31 39 40 44 46 VSS
c19 48 VSS 0.00113024f $X=0.8915 $Y=0.1915
c20 46 VSS 5.62354e-19 $X=0.8915 $Y=0.1015
c21 45 VSS 0.00169587f $X=0.8915 $Y=0.09
c22 44 VSS 0.00352425f $X=0.889 $Y=0.113
c23 42 VSS 0.00118619f $X=0.8915 $Y=0.216
c24 40 VSS 9.93081e-19 $X=0.792 $Y=0.225
c25 39 VSS 0.00330792f $X=0.774 $Y=0.225
c26 31 VSS 0.0116023f $X=0.882 $Y=0.225
c27 30 VSS 9.95001e-19 $X=0.792 $Y=0.045
c28 29 VSS 0.00317729f $X=0.774 $Y=0.045
c29 28 VSS 0.00459282f $X=0.864 $Y=0.045
c30 24 VSS 0.00743883f $X=0.756 $Y=0.045
c31 21 VSS 0.0115671f $X=0.882 $Y=0.045
c32 19 VSS 0.00492775f $X=0.862 $Y=0.2025
c33 15 VSS 0.00724558f $X=0.756 $Y=0.2025
c34 11 VSS 6.63935e-19 $X=0.773 $Y=0.2025
c35 9 VSS 3.34937e-19 $X=0.862 $Y=0.0675
c36 1 VSS 6.63935e-19 $X=0.773 $Y=0.0675
r37 47 48 1.55612 $w=1.9e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.8915
+ $Y=0.167 $X2=0.8915 $Y2=0.1915
r38 45 46 0.730426 $w=1.9e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8915
+ $Y=0.09 $X2=0.8915 $Y2=0.1015
r39 44 47 3.42982 $w=1.9e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.8915
+ $Y=0.113 $X2=0.8915 $Y2=0.167
r40 44 46 0.730426 $w=1.9e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.8915
+ $Y=0.113 $X2=0.8915 $Y2=0.1015
r41 42 48 1.55612 $w=1.9e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.8915
+ $Y=0.216 $X2=0.8915 $Y2=0.1915
r42 41 45 2.28655 $w=1.9e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.8915
+ $Y=0.054 $X2=0.8915 $Y2=0.09
r43 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.225 $X2=0.792 $Y2=0.225
r44 37 40 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.225 $X2=0.792 $Y2=0.225
r45 33 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.225 $X2=0.774 $Y2=0.225
r46 31 42 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.225 $X2=0.8915 $Y2=0.216
r47 31 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.225 $X2=0.864 $Y2=0.225
r48 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.045 $X2=0.792 $Y2=0.045
r49 27 30 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.045 $X2=0.792 $Y2=0.045
r50 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.045 $X2=0.864
+ $Y2=0.045
r51 23 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.045 $X2=0.774 $Y2=0.045
r52 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.045 $X2=0.756
+ $Y2=0.045
r53 21 41 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.045 $X2=0.8915 $Y2=0.054
r54 21 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.045 $X2=0.864 $Y2=0.045
r55 19 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.225 $X2=0.864
+ $Y2=0.225
r56 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2025 $X2=0.862 $Y2=0.2025
r57 15 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.225 $X2=0.756
+ $Y2=0.225
r58 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r59 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r60 9 28 19.4196 $w=2.4e-08 $l=2.25e-08 $layer=LISD $thickness=2.8e-08 $X=0.864
+ $Y=0.0675 $X2=0.864 $Y2=0.045
r61 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.847
+ $Y=0.0675 $X2=0.862 $Y2=0.0675
r62 5 24 19.4196 $w=2.4e-08 $l=2.25e-08 $layer=LISD $thickness=2.8e-08 $X=0.756
+ $Y=0.0675 $X2=0.756 $Y2=0.045
r63 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
r64 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
.ends

.subckt PM_DLLX3_ASAP7_75T_SRAM%10 1 6 9 VSS
c7 9 VSS 0.0266424f $X=0.38 $Y=0.0675
c8 6 VSS 3.25039e-19 $X=0.395 $Y=0.0675
c9 4 VSS 3.22674e-19 $X=0.322 $Y=0.0675
r10 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r11 4 9 14.8325 $w=8.1e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.322
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
r12 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_DLLX3_ASAP7_75T_SRAM%11 1 6 9 VSS
c9 9 VSS 0.0211025f $X=0.488 $Y=0.2295
c10 6 VSS 3.14771e-19 $X=0.503 $Y=0.2295
c11 4 VSS 2.84146e-19 $X=0.43 $Y=0.2295
r12 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r13 4 9 44.4974 $w=2.7e-08 $l=5.8e-08 $layer=LISD $thickness=2.8e-08 $X=0.43
+ $Y=0.2295 $X2=0.488 $Y2=0.2295
r14 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2295 $X2=0.43 $Y2=0.2295
.ends

.subckt PM_DLLX3_ASAP7_75T_SRAM%12 1 2 VSS
c0 1 VSS 0.00220425f $X=0.503 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0405 $X2=0.469 $Y2=0.0405
.ends

.subckt PM_DLLX3_ASAP7_75T_SRAM%13 1 2 VSS
c1 1 VSS 0.00201018f $X=0.341 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends


* END of "./DLLx3_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt DLLx3_ASAP7_75t_SRAM  VSS VDD CLK D Q
* 
* Q	Q
* D	D
* CLK	CLK
M0 VSS N_CLK_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.027
M1 N_6_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_10_M2_d N_D_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_8_M3_d N_4_M3_g N_10_M3_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M4 N_12_M4_d N_6_M4_g N_8_M4_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.449
+ $Y=0.027
M5 VSS N_7_M5_g N_12_M5_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.027
M6 N_7_M6_d N_8_M6_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557 $Y=0.027
M7 N_Q_M7_d N_8_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M8 N_Q_M8_d N_8_M8_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773 $Y=0.027
M9 N_Q_M9_d N_8_M9_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827 $Y=0.027
M10 VDD N_CLK_M10_g N_4_M10_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M11 N_6_M11_d N_4_M11_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M12 N_13_M12_d N_D_M12_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M13 N_8_M13_d N_6_M13_g N_13_M13_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M14 N_11_M14_d N_4_M14_g N_8_M14_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1
+ $X=0.395 $Y=0.216
M15 VDD N_7_M15_g N_11_M15_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.503
+ $Y=0.216
M16 N_7_M16_d N_8_M16_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.557
+ $Y=0.216
M17 N_Q_M17_d N_8_M17_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M18 N_Q_M18_d N_8_M18_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
M19 N_Q_M19_d N_8_M19_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.162
*
* 
* .include "DLLx3_ASAP7_75t_SRAM.pex.sp.DLLX3_ASAP7_75T_SRAM.pxi"
* BEGIN of "./DLLx3_ASAP7_75t_SRAM.pex.sp.DLLX3_ASAP7_75T_SRAM.pxi"
* File: DLLx3_ASAP7_75t_SRAM.pex.sp.DLLX3_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:29:00 2017
* 
x_PM_DLLX3_ASAP7_75T_SRAM%CLK N_CLK_M0_g N_CLK_c_11_p N_CLK_M10_g CLK N_CLK_c_3_p
+ N_CLK_c_4_p VSS PM_DLLX3_ASAP7_75T_SRAM%CLK
x_PM_DLLX3_ASAP7_75T_SRAM%4 N_4_M1_g N_4_M11_g N_4_M3_g N_4_c_38_p N_4_M14_g
+ N_4_M0_s N_4_c_20_n N_4_M10_s N_4_c_21_n N_4_c_22_n N_4_c_23_n N_4_c_24_n
+ N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_48_p N_4_c_28_n N_4_c_29_n N_4_c_30_n
+ N_4_c_31_n N_4_c_53_p N_4_c_32_n N_4_c_36_p N_4_c_40_p VSS
+ PM_DLLX3_ASAP7_75T_SRAM%4
x_PM_DLLX3_ASAP7_75T_SRAM%D N_D_M2_g N_D_c_64_n N_D_M12_g D N_D_c_69_p VSS
+ PM_DLLX3_ASAP7_75T_SRAM%D
x_PM_DLLX3_ASAP7_75T_SRAM%6 N_6_c_87_n N_6_M13_g N_6_M4_g N_6_c_90_n N_6_M1_d
+ N_6_M11_d N_6_c_91_n N_6_c_92_n N_6_c_84_n N_6_c_94_n N_6_c_95_n N_6_c_85_n
+ N_6_c_97_n N_6_c_109_n N_6_c_98_n N_6_c_111_n N_6_c_141_p N_6_c_100_n
+ N_6_c_131_p N_6_c_103_n N_6_c_119_p N_6_c_120_p N_6_c_86_n N_6_c_116_n
+ N_6_c_117_n VSS PM_DLLX3_ASAP7_75T_SRAM%6
x_PM_DLLX3_ASAP7_75T_SRAM%7 N_7_M5_g N_7_c_160_n N_7_M15_g N_7_M6_d N_7_c_161_n
+ N_7_M16_d N_7_c_162_n N_7_c_170_p N_7_c_169_p N_7_c_167_p N_7_c_179_p
+ N_7_c_171_p N_7_c_168_p N_7_c_177_p N_7_c_163_n N_7_c_164_n N_7_c_165_n VSS
+ PM_DLLX3_ASAP7_75T_SRAM%7
x_PM_DLLX3_ASAP7_75T_SRAM%8 N_8_M6_g N_8_c_213_n N_8_M16_g N_8_M7_g N_8_M17_g
+ N_8_M8_g N_8_M18_g N_8_M9_g N_8_c_225_p N_8_M19_g N_8_M3_d N_8_M4_s N_8_M13_d
+ N_8_c_180_n N_8_M14_s N_8_c_193_n N_8_c_187_n N_8_c_181_n N_8_c_188_n
+ N_8_c_196_n N_8_c_183_n N_8_c_198_n N_8_c_216_n N_8_c_199_n N_8_c_200_n
+ N_8_c_201_n N_8_c_250_p N_8_c_184_n N_8_c_228_p N_8_c_185_n N_8_c_221_n
+ N_8_c_224_n N_8_c_207_n VSS PM_DLLX3_ASAP7_75T_SRAM%8
x_PM_DLLX3_ASAP7_75T_SRAM%Q N_Q_M8_d N_Q_M7_d N_Q_M9_d N_Q_M18_d N_Q_M17_d
+ N_Q_c_253_n N_Q_M19_d N_Q_c_255_n N_Q_c_257_n N_Q_c_259_n N_Q_c_261_n
+ N_Q_c_263_n N_Q_c_265_n N_Q_c_266_n Q N_Q_c_269_n VSS PM_DLLX3_ASAP7_75T_SRAM%Q
x_PM_DLLX3_ASAP7_75T_SRAM%10 N_10_M2_d N_10_M3_s N_10_c_270_n VSS
+ PM_DLLX3_ASAP7_75T_SRAM%10
x_PM_DLLX3_ASAP7_75T_SRAM%11 N_11_M14_d N_11_M15_s N_11_c_278_n VSS
+ PM_DLLX3_ASAP7_75T_SRAM%11
x_PM_DLLX3_ASAP7_75T_SRAM%12 N_12_M5_s N_12_M4_d VSS PM_DLLX3_ASAP7_75T_SRAM%12
x_PM_DLLX3_ASAP7_75T_SRAM%13 N_13_M13_s N_13_M12_d VSS PM_DLLX3_ASAP7_75T_SRAM%13
cc_1 N_CLK_M0_g N_4_M1_g 0.00268443f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 CLK N_4_c_20_n 2.66516e-19 $X=0.082 $Y=0.119 $X2=0.056 $Y2=0.054
cc_3 N_CLK_c_3_p N_4_c_21_n 2.66516e-19 $X=0.081 $Y=0.135 $X2=0.056 $Y2=0.216
cc_4 N_CLK_c_4_p N_4_c_22_n 0.00126555f $X=0.081 $Y=0.1305 $X2=0.018 $Y2=0.144
cc_5 CLK N_4_c_23_n 3.98992e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.081
cc_6 CLK N_4_c_24_n 0.00126555f $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.1125
cc_7 N_CLK_c_3_p N_4_c_25_n 0.00127356f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.189
cc_8 CLK N_4_c_26_n 4.98319e-19 $X=0.082 $Y=0.119 $X2=0.054 $Y2=0.036
cc_9 N_CLK_c_3_p N_4_c_27_n 4.98319e-19 $X=0.081 $Y=0.135 $X2=0.054 $Y2=0.234
cc_10 N_CLK_c_4_p N_4_c_28_n 4.17e-19 $X=0.081 $Y=0.1305 $X2=0.152 $Y2=0.135
cc_11 N_CLK_c_11_p N_4_c_29_n 0.00116357f $X=0.081 $Y=0.135 $X2=0.152 $Y2=0.135
cc_12 N_CLK_c_3_p N_4_c_30_n 0.00122788f $X=0.081 $Y=0.135 $X2=0.033 $Y2=0.153
cc_13 N_CLK_c_3_p N_4_c_31_n 0.00197837f $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.153
cc_14 CLK N_4_c_32_n 5.08945e-19 $X=0.082 $Y=0.119 $X2=0.229 $Y2=0.153
cc_15 N_CLK_c_3_p N_4_c_32_n 0.00150524f $X=0.081 $Y=0.135 $X2=0.229 $Y2=0.153
cc_16 CLK N_6_c_84_n 6.45949e-19 $X=0.082 $Y=0.119 $X2=0.018 $Y2=0.189
cc_17 N_CLK_c_3_p N_6_c_85_n 6.45949e-19 $X=0.081 $Y=0.135 $X2=0.0505 $Y2=0.036
cc_18 CLK N_6_c_86_n 7.98675e-19 $X=0.082 $Y=0.119 $X2=0.152 $Y2=0.135
cc_19 N_4_M3_g N_D_M2_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_20 N_4_c_29_n N_D_c_64_n 2.01856e-19 $X=0.152 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 N_4_c_36_p D 0.00117371f $X=0.317 $Y=0.153 $X2=0.082 $Y2=0.119
cc_22 N_4_M3_g N_6_c_87_n 0.00355599f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_23 N_4_c_38_p N_6_c_87_n 0.00101396f $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.054
cc_24 N_4_M3_g N_6_M4_g 0.00355599f $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_25 N_4_c_40_p N_6_c_90_n 3.2936e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.126
cc_26 N_4_c_31_n N_6_c_91_n 0.00243501f $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_27 N_4_c_36_p N_6_c_92_n 2.3925e-19 $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_28 N_4_c_28_n N_6_c_84_n 9.58415e-19 $X=0.152 $Y=0.135 $X2=0 $Y2=0
cc_29 N_4_c_32_n N_6_c_94_n 2.3925e-19 $X=0.229 $Y=0.153 $X2=0 $Y2=0
cc_30 N_4_c_36_p N_6_c_95_n 2.75285e-19 $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_31 N_4_c_31_n N_6_c_85_n 0.00467935f $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_32 N_4_c_32_n N_6_c_97_n 2.75285e-19 $X=0.229 $Y=0.153 $X2=0 $Y2=0
cc_33 N_4_c_48_p N_6_c_98_n 0.00396181f $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_34 N_4_c_36_p N_6_c_98_n 0.00119509f $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_35 N_4_c_31_n N_6_c_100_n 3.89771e-19 $X=0.189 $Y=0.153 $X2=0 $Y2=0
cc_36 N_4_c_36_p N_6_c_100_n 0.0160263f $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_37 N_4_c_40_p N_6_c_100_n 8.49272e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_53_p N_6_c_103_n 0.00115166f $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_39 N_4_c_40_p N_6_c_103_n 0.00433569f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_M3_g N_7_M5_g 2.82885e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_41 N_4_c_40_p N_8_c_180_n 0.00195725f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_42 N_4_M3_g N_8_c_181_n 2.63086e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_4_c_40_p N_8_c_181_n 0.00122664f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_44 N_4_c_40_p N_8_c_183_n 0.00419136f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_45 N_4_c_40_p N_8_c_184_n 2.60642e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_53_p N_8_c_185_n 9.23088e-19 $X=0.405 $Y=0.153 $X2=0 $Y2=0
cc_47 N_4_c_36_p N_10_c_270_n 8.32437e-19 $X=0.317 $Y=0.153 $X2=0 $Y2=0
cc_48 N_D_M2_g N_6_c_87_n 0.00341068f $X=0.297 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_49 N_D_c_64_n N_6_c_87_n 0.00101372f $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_50 D N_6_c_92_n 0.00115278f $X=0.297 $Y=0.1165 $X2=0.018 $Y2=0.144
cc_51 N_D_c_69_p N_6_c_95_n 0.00115278f $X=0.297 $Y=0.135 $X2=0.027 $Y2=0.036
cc_52 N_D_c_69_p N_6_c_109_n 0.00115278f $X=0.297 $Y=0.135 $X2=0.054 $Y2=0.234
cc_53 D N_6_c_98_n 0.00124619f $X=0.297 $Y=0.1165 $X2=0.047 $Y2=0.234
cc_54 D N_6_c_111_n 0.00216863f $X=0.297 $Y=0.1165 $X2=0.152 $Y2=0.135
cc_55 D N_6_c_100_n 8.86605e-19 $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_56 N_D_c_69_p N_6_c_100_n 3.97512e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_57 D N_6_c_103_n 0.00216863f $X=0.297 $Y=0.1165 $X2=0.189 $Y2=0.144
cc_58 D N_6_c_86_n 0.00115278f $X=0.297 $Y=0.1165 $X2=0.152 $Y2=0.135
cc_59 D N_6_c_116_n 0.00115278f $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_60 N_D_c_69_p N_6_c_117_n 0.00115278f $X=0.297 $Y=0.135 $X2=0.405 $Y2=0.135
cc_61 N_D_c_69_p N_8_c_180_n 3.88702e-19 $X=0.297 $Y=0.135 $X2=0.054 $Y2=0.234
cc_62 N_D_c_69_p N_8_c_187_n 8.77202e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_63 D N_8_c_188_n 2.05539e-19 $X=0.297 $Y=0.1165 $X2=0 $Y2=0
cc_64 D N_10_c_270_n 0.00428733f $X=0.297 $Y=0.1165 $X2=0.405 $Y2=0.0675
cc_65 N_D_c_69_p N_13_M13_s 3.05674e-19 $X=0.297 $Y=0.135 $X2=0.135 $Y2=0.054
cc_66 N_6_M4_g N_7_M5_g 0.00341068f $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_67 N_6_c_119_p N_7_M5_g 0.00199227f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_68 N_6_c_120_p N_7_M5_g 4.91626e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_69 N_6_c_119_p N_7_c_160_n 4.44368e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.135
cc_70 N_6_c_119_p N_7_c_161_n 5.31675e-19 $X=0.513 $Y=0.18 $X2=0.082 $Y2=0.119
cc_71 N_6_c_119_p N_7_c_162_n 0.00169036f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.1305
cc_72 N_6_c_120_p N_7_c_163_n 5.94045e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_73 N_6_c_119_p N_7_c_164_n 0.00305515f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_74 N_6_c_119_p N_7_c_165_n 5.97916e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_75 N_6_M4_g N_8_M6_g 2.13359e-19 $X=0.459 $Y=0.0405 $X2=0.081 $Y2=0.054
cc_76 N_6_c_119_p N_8_M6_g 0.00305655f $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.054
cc_77 N_6_c_100_n N_8_c_180_n 2.84357e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_78 N_6_c_103_n N_8_c_180_n 0.00130164f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_79 N_6_c_131_p N_8_c_193_n 7.16323e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_80 N_6_c_100_n N_8_c_187_n 5.53186e-19 $X=0.414 $Y=0.189 $X2=0 $Y2=0
cc_81 N_6_c_131_p N_8_c_188_n 3.48842e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_82 N_6_c_131_p N_8_c_196_n 2.01793e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_83 N_6_M4_g N_8_c_183_n 2.93184e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_84 N_6_M4_g N_8_c_198_n 3.72919e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_85 N_6_c_119_p N_8_c_199_n 4.41338e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_86 N_6_c_119_p N_8_c_200_n 7.92645e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_87 N_6_c_120_p N_8_c_201_n 0.00100546f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_88 N_6_M4_g N_8_c_184_n 2.27241e-19 $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_89 N_6_c_141_p N_8_c_184_n 2.46239e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_90 N_6_c_141_p N_8_c_185_n 0.00694438f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_91 N_6_c_119_p N_8_c_185_n 0.00195448f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_92 N_6_c_120_p N_8_c_185_n 2.84312e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_93 N_6_c_90_n N_8_c_207_n 0.00271026f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_94 N_6_c_141_p N_8_c_207_n 6.73646e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_95 N_6_c_119_p N_8_c_207_n 5.95032e-19 $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_96 N_6_c_120_p N_8_c_207_n 0.00182777f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_97 N_6_c_87_n N_10_c_270_n 0.00639848f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_98 N_6_c_103_n N_10_c_270_n 0.00135407f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_99 N_6_c_119_p N_11_M15_s 2.34172e-19 $X=0.513 $Y=0.18 $X2=0.081 $Y2=0.216
cc_100 N_6_M4_g N_11_c_278_n 0.00200065f $X=0.459 $Y=0.0405 $X2=0 $Y2=0
cc_101 N_6_c_90_n N_11_c_278_n 0.0013957f $X=0.464 $Y=0.179 $X2=0 $Y2=0
cc_102 N_6_c_131_p N_11_c_278_n 7.09553e-19 $X=0.45 $Y=0.189 $X2=0 $Y2=0
cc_103 N_6_c_119_p N_11_c_278_n 0.00230185f $X=0.513 $Y=0.18 $X2=0 $Y2=0
cc_104 N_7_M5_g N_8_M6_g 0.00268443f $X=0.513 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_105 N_7_c_167_p N_8_M6_g 4.17397e-19 $X=0.58 $Y=0.036 $X2=0.135 $Y2=0.054
cc_106 N_7_c_168_p N_8_c_213_n 3.44688e-19 $X=0.621 $Y=0.14 $X2=0.135 $Y2=0.135
cc_107 N_7_c_169_p N_8_c_188_n 0.00177955f $X=0.522 $Y=0.036 $X2=0 $Y2=0
cc_108 N_7_c_170_p N_8_c_198_n 0.00177955f $X=0.513 $Y=0.082 $X2=0 $Y2=0
cc_109 N_7_c_171_p N_8_c_216_n 2.88064e-19 $X=0.621 $Y=0.122 $X2=0.189 $Y2=0.153
cc_110 N_7_c_167_p N_8_c_199_n 6.9494e-19 $X=0.58 $Y=0.036 $X2=0.405 $Y2=0.153
cc_111 N_7_c_168_p N_8_c_199_n 9.37002e-19 $X=0.621 $Y=0.14 $X2=0.405 $Y2=0.153
cc_112 N_7_M5_g N_8_c_201_n 4.06683e-19 $X=0.513 $Y=0.0405 $X2=0.229 $Y2=0.153
cc_113 N_7_c_170_p N_8_c_201_n 0.00116089f $X=0.513 $Y=0.082 $X2=0.229 $Y2=0.153
cc_114 N_7_c_161_n N_8_c_221_n 2.11538e-19 $X=0.592 $Y=0.0405 $X2=0 $Y2=0
cc_115 N_7_c_177_p N_8_c_221_n 0.00133609f $X=0.621 $Y=0.165 $X2=0 $Y2=0
cc_116 N_7_c_165_n N_8_c_221_n 5.94743e-19 $X=0.612 $Y=0.234 $X2=0 $Y2=0
cc_117 N_7_c_179_p N_8_c_224_n 4.45934e-19 $X=0.621 $Y=0.097 $X2=0.018 $Y2=0.153
cc_118 N_8_c_225_p N_Q_M8_d 3.7444e-19 $X=0.837 $Y=0.136 $X2=0.135 $Y2=0.054
cc_119 N_8_c_225_p N_Q_M18_d 3.82547e-19 $X=0.837 $Y=0.136 $X2=0 $Y2=0
cc_120 N_8_c_225_p N_Q_c_253_n 8.43851e-19 $X=0.837 $Y=0.136 $X2=0.405
+ $Y2=0.2295
cc_121 N_8_c_228_p N_Q_c_253_n 3.0124e-19 $X=0.783 $Y=0.153 $X2=0.405 $Y2=0.2295
cc_122 N_8_M9_g N_Q_c_255_n 4.75199e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_123 N_8_c_225_p N_Q_c_255_n 8.37011e-19 $X=0.837 $Y=0.136 $X2=0 $Y2=0
cc_124 N_8_c_225_p N_Q_c_257_n 7.60428e-19 $X=0.837 $Y=0.136 $X2=0 $Y2=0
cc_125 N_8_c_224_n N_Q_c_257_n 6.32721e-19 $X=0.783 $Y=0.136 $X2=0 $Y2=0
cc_126 N_8_c_225_p N_Q_c_259_n 3.08094e-19 $X=0.837 $Y=0.136 $X2=0.018 $Y2=0.081
cc_127 N_8_c_228_p N_Q_c_259_n 2.86931e-19 $X=0.783 $Y=0.153 $X2=0.018 $Y2=0.081
cc_128 N_8_M8_g N_Q_c_261_n 3.25912e-19 $X=0.783 $Y=0.0675 $X2=0.018 $Y2=0.1125
cc_129 N_8_c_224_n N_Q_c_261_n 8.86582e-19 $X=0.783 $Y=0.136 $X2=0.018
+ $Y2=0.1125
cc_130 N_8_M9_g N_Q_c_263_n 4.69796e-19 $X=0.837 $Y=0.0675 $X2=0.018 $Y2=0.162
cc_131 N_8_c_225_p N_Q_c_263_n 8.27998e-19 $X=0.837 $Y=0.136 $X2=0.018 $Y2=0.162
cc_132 N_8_c_228_p N_Q_c_265_n 3.66411e-19 $X=0.783 $Y=0.153 $X2=0.047 $Y2=0.036
cc_133 N_8_M8_g N_Q_c_266_n 3.55084e-19 $X=0.783 $Y=0.0675 $X2=0.0505 $Y2=0.036
cc_134 N_8_c_224_n N_Q_c_266_n 6.56888e-19 $X=0.783 $Y=0.136 $X2=0.0505
+ $Y2=0.036
cc_135 N_8_c_225_p Q 3.39128e-19 $X=0.837 $Y=0.136 $X2=0.054 $Y2=0.234
cc_136 N_8_c_224_n N_Q_c_269_n 9.8581e-19 $X=0.783 $Y=0.136 $X2=0.047 $Y2=0.234
cc_137 N_8_c_180_n N_10_c_270_n 0.00119636f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_138 N_8_c_188_n N_10_c_270_n 4.50844e-19 $X=0.45 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_139 N_8_c_196_n N_10_c_270_n 0.00394776f $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_140 N_8_c_180_n N_11_c_278_n 0.00186787f $X=0.378 $Y=0.2025 $X2=0.405
+ $Y2=0.0675
cc_141 N_8_c_193_n N_11_c_278_n 0.00343017f $X=0.45 $Y=0.234 $X2=0.405
+ $Y2=0.0675
cc_142 N_8_c_196_n N_11_c_278_n 5.72355e-19 $X=0.432 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_143 N_8_c_250_p N_11_c_278_n 0.00116187f $X=0.459 $Y=0.225 $X2=0.405
+ $Y2=0.0675

* END of "./DLLx3_ASAP7_75t_SRAM.pex.sp.DLLX3_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

