// This is the LdSelMux datapath block.

module LdSelMux (
	input [31:0] raw_dmem,
	input [2:0] LdSel,

	output [31:0] wb_dmem 
);



endmodule