* File: BUFx10_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:17:47 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx10_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx10_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx10_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:17:47 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX10_ASAP7_75T_SRAM%A 2 7 10 13 15 23 27 VSS
c21 27 VSS 0.00191995f $X=0.081 $Y=0.135
c22 23 VSS 0.0244917f $X=0.0565 $Y=0.1325
c23 13 VSS 0.00510508f $X=0.135 $Y=0.135
c24 10 VSS 0.0605852f $X=0.135 $Y=0.0675
c25 2 VSS 0.0649407f $X=0.081 $Y=0.0675
r26 23 27 1.66358 $w=1.8e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.0565
+ $Y=0.135 $X2=0.081 $Y2=0.135
r27 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r28 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r29 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r30 5 27 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r31 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r32 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX10_ASAP7_75T_SRAM%4 2 5 7 10 15 18 23 26 31 34 39 42 47 50 55 58 63
+ 66 71 74 77 79 81 82 86 87 90 92 94 102 103 126 130 131 135 140 145 149 VSS
c45 146 VSS 0.00214869f $X=0.126 $Y=0.234
c46 145 VSS 0.00263626f $X=0.135 $Y=0.234
c47 140 VSS 0.00188321f $X=0.108 $Y=0.234
c48 136 VSS 0.00214869f $X=0.126 $Y=0.036
c49 135 VSS 0.00263626f $X=0.135 $Y=0.036
c50 131 VSS 0.0106734f $X=0.108 $Y=0.036
c51 130 VSS 0.00188321f $X=0.108 $Y=0.036
c52 126 VSS 0.00781559f $X=0.675 $Y=0.135
c53 103 VSS 7.15556e-19 $X=0.221 $Y=0.135
c54 102 VSS 0.00267522f $X=0.199 $Y=0.135
c55 94 VSS 0.00385172f $X=0.135 $Y=0.225
c56 92 VSS 0.00385172f $X=0.135 $Y=0.126
c57 90 VSS 0.0106734f $X=0.108 $Y=0.2025
c58 86 VSS 5.25448e-19 $X=0.125 $Y=0.2025
c59 81 VSS 5.25448e-19 $X=0.125 $Y=0.0675
c60 77 VSS 0.00293966f $X=0.675 $Y=0.135
c61 74 VSS 0.0639847f $X=0.675 $Y=0.0675
c62 69 VSS 0.00178186f $X=0.621 $Y=0.135
c63 66 VSS 0.0638949f $X=0.621 $Y=0.0675
c64 61 VSS 0.00160407f $X=0.567 $Y=0.135
c65 58 VSS 0.0636879f $X=0.567 $Y=0.0675
c66 53 VSS 0.00166943f $X=0.513 $Y=0.135
c67 50 VSS 0.0636879f $X=0.513 $Y=0.0675
c68 45 VSS 0.00160407f $X=0.459 $Y=0.135
c69 42 VSS 0.0636879f $X=0.459 $Y=0.0675
c70 37 VSS 0.00166943f $X=0.405 $Y=0.135
c71 34 VSS 0.0636879f $X=0.405 $Y=0.0675
c72 29 VSS 0.00160407f $X=0.351 $Y=0.135
c73 26 VSS 0.0636879f $X=0.351 $Y=0.0675
c74 21 VSS 0.00166943f $X=0.297 $Y=0.135
c75 18 VSS 0.0636879f $X=0.297 $Y=0.0675
c76 13 VSS 0.0016373f $X=0.243 $Y=0.135
c77 10 VSS 0.0636879f $X=0.243 $Y=0.0675
c78 5 VSS 0.0017237f $X=0.189 $Y=0.135
c79 2 VSS 0.0615394f $X=0.189 $Y=0.0675
r80 146 147 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r81 145 147 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r82 140 146 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r83 136 137 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r84 135 137 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r85 130 136 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r86 130 131 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r87 123 126 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.135 $X2=0.675 $Y2=0.135
r88 120 123 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.621 $Y2=0.135
r89 117 120 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r90 114 117 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r91 111 114 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r92 108 111 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r93 105 108 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r94 102 103 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.199
+ $Y=0.135 $X2=0.221 $Y2=0.135
r95 100 105 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r96 100 103 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.221 $Y2=0.135
r97 97 102 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.199 $Y2=0.135
r98 95 149 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.135 $Y2=0.135
r99 95 97 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.189 $Y2=0.135
r100 94 145 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.234
r101 93 149 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.135
r102 93 94 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.225
r103 92 149 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.135
r104 91 135 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.036
r105 91 92 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.126
r106 90 140 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r107 87 90 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r108 86 90 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r109 85 131 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.108 $Y=0.0675 $X2=0.108 $Y2=0.036
r110 82 85 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r111 81 85 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r112 77 126 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.135
+ $X2=0.675 $Y2=0.135
r113 77 79 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2025
r114 74 77 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0675 $X2=0.675 $Y2=0.135
r115 69 123 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135
+ $X2=0.621 $Y2=0.135
r116 69 71 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2025
r117 66 69 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r118 61 120 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135
+ $X2=0.567 $Y2=0.135
r119 61 63 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.135 $X2=0.567 $Y2=0.2025
r120 58 61 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.0675 $X2=0.567 $Y2=0.135
r121 53 117 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135
+ $X2=0.513 $Y2=0.135
r122 53 55 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r123 50 53 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r124 45 114 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135
+ $X2=0.459 $Y2=0.135
r125 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r126 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r127 37 111 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135
+ $X2=0.405 $Y2=0.135
r128 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r129 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r130 29 108 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135
+ $X2=0.351 $Y2=0.135
r131 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r132 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r133 21 105 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135
+ $X2=0.297 $Y2=0.135
r134 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.135 $X2=0.297 $Y2=0.2025
r135 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.0675 $X2=0.297 $Y2=0.135
r136 13 100 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135
+ $X2=0.243 $Y2=0.135
r137 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.2025
r138 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.135
r139 5 97 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r140 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r141 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_BUFX10_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 21 22 26 27 31 32 36 37 41
+ 42 46 47 68 87 92 94 VSS
c24 96 VSS 0.00297428f $X=0.729 $Y=0.1845
c25 94 VSS 2.8404e-19 $X=0.729 $Y=0.13275
c26 93 VSS 0.00537436f $X=0.729 $Y=0.126
c27 92 VSS 4.56292e-19 $X=0.7295 $Y=0.1395
c28 90 VSS 0.00239816f $X=0.729 $Y=0.225
c29 88 VSS 0.00294383f $X=0.7045 $Y=0.234
c30 87 VSS 0.0524882f $X=0.689 $Y=0.234
c31 70 VSS 0.00588366f $X=0.72 $Y=0.234
c32 69 VSS 0.00294383f $X=0.7045 $Y=0.036
c33 68 VSS 0.0524882f $X=0.689 $Y=0.036
c34 67 VSS 0.00889316f $X=0.648 $Y=0.036
c35 64 VSS 0.00888519f $X=0.54 $Y=0.036
c36 61 VSS 0.00888519f $X=0.432 $Y=0.036
c37 58 VSS 0.00888519f $X=0.324 $Y=0.036
c38 54 VSS 0.00876044f $X=0.216 $Y=0.036
c39 51 VSS 0.00588366f $X=0.72 $Y=0.036
c40 50 VSS 0.00889316f $X=0.648 $Y=0.2025
c41 46 VSS 7.1893e-19 $X=0.665 $Y=0.2025
c42 45 VSS 0.00888519f $X=0.54 $Y=0.2025
c43 41 VSS 7.1893e-19 $X=0.557 $Y=0.2025
c44 40 VSS 0.00888519f $X=0.432 $Y=0.2025
c45 36 VSS 7.1893e-19 $X=0.449 $Y=0.2025
c46 35 VSS 0.00888519f $X=0.324 $Y=0.2025
c47 31 VSS 7.1893e-19 $X=0.341 $Y=0.2025
c48 30 VSS 0.00876044f $X=0.216 $Y=0.2025
c49 26 VSS 7.1893e-19 $X=0.233 $Y=0.2025
c50 21 VSS 7.1893e-19 $X=0.665 $Y=0.0675
c51 16 VSS 7.1893e-19 $X=0.557 $Y=0.0675
c52 11 VSS 7.1893e-19 $X=0.449 $Y=0.0675
c53 6 VSS 7.1893e-19 $X=0.341 $Y=0.0675
c54 1 VSS 7.1893e-19 $X=0.233 $Y=0.0675
r55 95 96 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.144 $X2=0.729 $Y2=0.1845
r56 93 94 0.458333 $w=1.8e-08 $l=6.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.126 $X2=0.729 $Y2=0.13275
r57 92 95 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.1395 $X2=0.729 $Y2=0.144
r58 92 94 0.458333 $w=1.8e-08 $l=6.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.1395 $X2=0.729 $Y2=0.13275
r59 90 96 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.225 $X2=0.729 $Y2=0.1845
r60 89 93 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.045 $X2=0.729 $Y2=0.126
r61 87 88 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.689
+ $Y=0.234 $X2=0.7045 $Y2=0.234
r62 85 87 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.689 $Y2=0.234
r63 82 85 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.648 $Y2=0.234
r64 79 82 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.54 $Y2=0.234
r65 76 79 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r66 72 76 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.324 $Y2=0.234
r67 70 90 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.234 $X2=0.729 $Y2=0.225
r68 70 88 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.234 $X2=0.7045 $Y2=0.234
r69 68 69 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.689
+ $Y=0.036 $X2=0.7045 $Y2=0.036
r70 66 68 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.689 $Y2=0.036
r71 66 67 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036 $X2=0.648
+ $Y2=0.036
r72 63 66 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.648 $Y2=0.036
r73 63 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r74 60 63 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.54 $Y2=0.036
r75 60 61 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r76 57 60 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r77 57 58 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r78 53 57 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.324 $Y2=0.036
r79 53 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r80 51 89 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.036 $X2=0.729 $Y2=0.045
r81 51 69 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.7045 $Y2=0.036
r82 50 85 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234 $X2=0.648
+ $Y2=0.234
r83 47 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.648 $Y2=0.2025
r84 46 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.648 $Y2=0.2025
r85 45 82 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r86 42 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r87 41 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r88 40 79 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r89 37 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r90 36 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r91 35 76 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r92 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r93 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r94 30 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r95 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r96 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r97 25 67 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.648
+ $Y=0.0675 $X2=0.648 $Y2=0.036
r98 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.648 $Y2=0.0675
r99 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0675 $X2=0.648 $Y2=0.0675
r100 20 64 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r101 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r102 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r103 15 61 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r104 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r105 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r106 10 58 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r107 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r108 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r109 5 54 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r110 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r111 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./BUFx10_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx10_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_4_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_4_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_4_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_4_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_4_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_4_M6_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_4_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_4_M8_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_4_M9_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 N_Y_M10_d N_4_M10_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M11 N_Y_M11_d N_4_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M12 N_4_M12_d N_A_M12_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M13 N_4_M13_d N_A_M13_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M14 N_Y_M14_d N_4_M14_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M15 N_Y_M15_d N_4_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M16 N_Y_M16_d N_4_M16_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M17 N_Y_M17_d N_4_M17_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M18 N_Y_M18_d N_4_M18_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M19 N_Y_M19_d N_4_M19_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M20 N_Y_M20_d N_4_M20_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M21 N_Y_M21_d N_4_M21_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M22 N_Y_M22_d N_4_M22_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M23 N_Y_M23_d N_4_M23_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
*
* 
* .include "BUFx10_ASAP7_75t_SRAM.pex.sp.BUFX10_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx10_ASAP7_75t_SRAM.pex.sp.BUFX10_ASAP7_75T_SRAM.pxi"
* File: BUFx10_ASAP7_75t_SRAM.pex.sp.BUFX10_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:17:47 2017
* 
x_PM_BUFX10_ASAP7_75T_SRAM%A N_A_M0_g N_A_M12_g N_A_M1_g N_A_c_3_p N_A_M13_g A
+ N_A_c_21_p VSS PM_BUFX10_ASAP7_75T_SRAM%A
x_PM_BUFX10_ASAP7_75T_SRAM%4 N_4_M2_g N_4_c_24_n N_4_M14_g N_4_M3_g N_4_M15_g
+ N_4_M4_g N_4_M16_g N_4_M5_g N_4_M17_g N_4_M6_g N_4_M18_g N_4_M7_g N_4_M19_g
+ N_4_M8_g N_4_M20_g N_4_M9_g N_4_M21_g N_4_M10_g N_4_M22_g N_4_M11_g N_4_c_65_p
+ N_4_M23_g N_4_M1_d N_4_M0_d N_4_M13_d N_4_M12_d N_4_c_28_n N_4_c_29_n
+ N_4_c_32_n N_4_c_35_n N_4_c_52_p N_4_c_66_p N_4_c_36_n N_4_c_38_n N_4_c_53_p
+ N_4_c_39_n N_4_c_64_p N_4_c_41_n VSS PM_BUFX10_ASAP7_75T_SRAM%4
x_PM_BUFX10_ASAP7_75T_SRAM%Y N_Y_M3_d N_Y_M2_d N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M6_d
+ N_Y_M9_d N_Y_M8_d N_Y_M11_d N_Y_M10_d N_Y_M15_d N_Y_M14_d N_Y_M17_d N_Y_M16_d
+ N_Y_M19_d N_Y_M18_d N_Y_M21_d N_Y_M20_d N_Y_M23_d N_Y_M22_d N_Y_c_67_n
+ N_Y_c_78_n Y N_Y_c_89_n VSS PM_BUFX10_ASAP7_75T_SRAM%Y
cc_1 N_A_M0_g N_4_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_A_M1_g N_4_M2_g 0.00284417f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A_c_3_p N_4_c_24_n 0.00153702f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_4 N_A_M1_g N_4_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_5 N_A_c_3_p N_4_M1_d 3.80485e-19 $X=0.135 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_6 N_A_c_3_p N_4_M13_d 3.80485e-19 $X=0.135 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_7 N_A_c_3_p N_4_c_28_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_8 N_A_M1_g N_4_c_29_n 6.45702e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.126
cc_9 N_A_c_3_p N_4_c_29_n 4.76064e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.126
cc_10 A N_4_c_29_n 6.96001e-19 $X=0.0565 $Y=0.1325 $X2=0.135 $Y2=0.126
cc_11 N_A_M1_g N_4_c_32_n 6.45702e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.225
cc_12 N_A_c_3_p N_4_c_32_n 4.76064e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.225
cc_13 A N_4_c_32_n 6.96001e-19 $X=0.0565 $Y=0.1325 $X2=0.135 $Y2=0.225
cc_14 N_A_c_3_p N_4_c_35_n 5.83755e-19 $X=0.135 $Y=0.135 $X2=0.199 $Y2=0.135
cc_15 N_A_c_3_p N_4_c_36_n 3.46853e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.036
cc_16 A N_4_c_36_n 5.37037e-19 $X=0.0565 $Y=0.1325 $X2=0.108 $Y2=0.036
cc_17 N_A_c_3_p N_4_c_38_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.036
cc_18 N_A_c_3_p N_4_c_39_n 3.46853e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.234
cc_19 A N_4_c_39_n 5.37037e-19 $X=0.0565 $Y=0.1325 $X2=0.108 $Y2=0.234
cc_20 N_A_c_3_p N_4_c_41_n 0.00105301f $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.135
cc_21 N_A_c_21_p N_4_c_41_n 9.54523e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_22 N_4_M3_g N_Y_c_67_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_23 N_4_M4_g N_Y_c_67_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_24 N_4_M5_g N_Y_c_67_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_25 N_4_M6_g N_Y_c_67_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_4_M7_g N_Y_c_67_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_4_M8_g N_Y_c_67_n 4.28653e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_28 N_4_M9_g N_Y_c_67_n 4.28653e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_29 N_4_M10_g N_Y_c_67_n 4.28653e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_4_M11_g N_Y_c_67_n 4.28653e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_4_c_52_p N_Y_c_67_n 0.00875941f $X=0.221 $Y=0.135 $X2=0 $Y2=0
cc_32 N_4_c_53_p N_Y_c_67_n 3.93194e-19 $X=0.135 $Y=0.036 $X2=0 $Y2=0
cc_33 N_4_M3_g N_Y_c_78_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_34 N_4_M4_g N_Y_c_78_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_4_M5_g N_Y_c_78_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_4_M6_g N_Y_c_78_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_4_M7_g N_Y_c_78_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_38 N_4_M8_g N_Y_c_78_n 4.28653e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_4_M9_g N_Y_c_78_n 4.28653e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_40 N_4_M10_g N_Y_c_78_n 4.28653e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_41 N_4_M11_g N_Y_c_78_n 4.28653e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_42 N_4_c_52_p N_Y_c_78_n 0.00875941f $X=0.221 $Y=0.135 $X2=0 $Y2=0
cc_43 N_4_c_64_p N_Y_c_78_n 3.93194e-19 $X=0.135 $Y=0.234 $X2=0 $Y2=0
cc_44 N_4_c_65_p N_Y_c_89_n 3.22307e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_45 N_4_c_66_p N_Y_c_89_n 0.00102787f $X=0.675 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx10_ASAP7_75t_SRAM.pex.sp.BUFX10_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx12_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:18:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx12_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx12_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx12_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:18:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX12_ASAP7_75T_SRAM%A 2 7 10 13 15 23 VSS
c21 23 VSS 0.0250318f $X=0.061 $Y=0.1325
c22 13 VSS 0.00838749f $X=0.135 $Y=0.135
c23 10 VSS 0.0611086f $X=0.135 $Y=0.0675
c24 2 VSS 0.0655089f $X=0.081 $Y=0.0675
r25 23 27 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r26 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r27 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r28 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r29 5 27 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r30 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r31 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX12_ASAP7_75T_SRAM%4 2 7 10 15 18 23 26 31 34 39 42 47 50 55 58 63 66
+ 71 74 79 82 87 90 93 95 97 98 102 103 106 108 110 115 116 124 129 131 132 139
+ 140 143 VSS
c63 140 VSS 0.00367046f $X=0.126 $Y=0.234
c64 139 VSS 0.00263512f $X=0.135 $Y=0.234
c65 132 VSS 0.00367046f $X=0.126 $Y=0.036
c66 131 VSS 0.00263512f $X=0.135 $Y=0.036
c67 129 VSS 0.0106727f $X=0.108 $Y=0.036
c68 124 VSS 2.42544e-19 $X=0.729 $Y=0.135
c69 115 VSS 0.00271998f $X=0.199 $Y=0.135
c70 110 VSS 0.00385172f $X=0.135 $Y=0.225
c71 108 VSS 0.00385172f $X=0.135 $Y=0.126
c72 106 VSS 0.0106727f $X=0.108 $Y=0.2025
c73 102 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c74 97 VSS 5.72268e-19 $X=0.125 $Y=0.0675
c75 93 VSS 0.0407297f $X=0.783 $Y=0.135
c76 90 VSS 0.0645347f $X=0.783 $Y=0.0675
c77 82 VSS 0.0644226f $X=0.729 $Y=0.0675
c78 74 VSS 0.0642127f $X=0.675 $Y=0.0675
c79 66 VSS 0.0642127f $X=0.621 $Y=0.0675
c80 58 VSS 0.0642127f $X=0.567 $Y=0.0675
c81 50 VSS 0.0642127f $X=0.513 $Y=0.0675
c82 42 VSS 0.0642127f $X=0.459 $Y=0.0675
c83 34 VSS 0.0642127f $X=0.405 $Y=0.0675
c84 26 VSS 0.0642127f $X=0.351 $Y=0.0675
c85 18 VSS 0.0642127f $X=0.297 $Y=0.0675
c86 10 VSS 0.0642127f $X=0.243 $Y=0.0675
c87 2 VSS 0.0620627f $X=0.189 $Y=0.0675
r88 140 141 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r89 139 141 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r90 136 140 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r91 132 133 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r92 131 133 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r93 128 132 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r94 128 129 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r95 121 124 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.729 $Y2=0.135
r96 118 121 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.567 $Y2=0.135
r97 115 116 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.199
+ $Y=0.135 $X2=0.221 $Y2=0.135
r98 113 118 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.405 $Y2=0.135
r99 113 116 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.221 $Y2=0.135
r100 111 143 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.135 $Y2=0.135
r101 111 115 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.199 $Y2=0.135
r102 110 139 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.234
r103 109 143 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.135
r104 109 110 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.225
r105 108 143 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.135
r106 107 131 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.036
r107 107 108 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.126
r108 106 136 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r109 103 106 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r110 102 106 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r111 101 129 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.108 $Y=0.0675 $X2=0.108 $Y2=0.036
r112 98 101 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r113 97 101 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r114 93 95 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.135 $X2=0.783 $Y2=0.2025
r115 90 93 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.135
r116 85 93 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.135 $X2=0.783 $Y2=0.135
r117 85 124 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.729 $Y=0.135
+ $X2=0.729 $Y2=0.135
r118 85 87 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.135 $X2=0.729 $Y2=0.2025
r119 82 85 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.135
r120 77 85 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.729 $Y2=0.135
r121 77 79 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2025
r122 74 77 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0675 $X2=0.675 $Y2=0.135
r123 69 77 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621
+ $Y=0.135 $X2=0.675 $Y2=0.135
r124 69 71 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2025
r125 66 69 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r126 61 69 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.567
+ $Y=0.135 $X2=0.621 $Y2=0.135
r127 61 121 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.567 $Y=0.135
+ $X2=0.567 $Y2=0.135
r128 61 63 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.135 $X2=0.567 $Y2=0.2025
r129 58 61 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.0675 $X2=0.567 $Y2=0.135
r130 53 61 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r131 53 55 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r132 50 53 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r133 45 53 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r134 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r135 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r136 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r137 37 118 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.405 $Y=0.135
+ $X2=0.405 $Y2=0.135
r138 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r139 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r140 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r141 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r142 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r143 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r144 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.135 $X2=0.297 $Y2=0.2025
r145 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.0675 $X2=0.297 $Y2=0.135
r146 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r147 13 113 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.243 $Y=0.135
+ $X2=0.243 $Y2=0.135
r148 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.2025
r149 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.135
r150 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r151 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r152 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_BUFX12_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 21 22 26 27 31 32 36 37 41
+ 42 46 47 51 52 56 57 81 103 108 110 VSS
c42 110 VSS 7.43984e-19 $X=0.837 $Y=0.144
c43 109 VSS 0.00538621f $X=0.837 $Y=0.126
c44 108 VSS 0.00538621f $X=0.839 $Y=0.1495
c45 104 VSS 0.00237022f $X=0.814 $Y=0.234
c46 103 VSS 0.064037f $X=0.8 $Y=0.234
c47 83 VSS 0.00564375f $X=0.828 $Y=0.234
c48 82 VSS 0.00237022f $X=0.814 $Y=0.036
c49 81 VSS 0.064037f $X=0.8 $Y=0.036
c50 80 VSS 0.00929752f $X=0.756 $Y=0.036
c51 77 VSS 0.00928955f $X=0.648 $Y=0.036
c52 74 VSS 0.00928955f $X=0.54 $Y=0.036
c53 71 VSS 0.00928955f $X=0.432 $Y=0.036
c54 68 VSS 0.00928955f $X=0.324 $Y=0.036
c55 64 VSS 0.00916652f $X=0.216 $Y=0.036
c56 61 VSS 0.00564375f $X=0.828 $Y=0.036
c57 60 VSS 0.00929752f $X=0.756 $Y=0.2025
c58 56 VSS 5.38922e-19 $X=0.773 $Y=0.2025
c59 55 VSS 0.00928955f $X=0.648 $Y=0.2025
c60 51 VSS 5.38922e-19 $X=0.665 $Y=0.2025
c61 50 VSS 0.00928955f $X=0.54 $Y=0.2025
c62 46 VSS 5.38922e-19 $X=0.557 $Y=0.2025
c63 45 VSS 0.00928955f $X=0.432 $Y=0.2025
c64 41 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c65 40 VSS 0.00928955f $X=0.324 $Y=0.2025
c66 36 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c67 35 VSS 0.00916652f $X=0.216 $Y=0.2025
c68 31 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c69 26 VSS 5.38922e-19 $X=0.773 $Y=0.0675
c70 21 VSS 5.38922e-19 $X=0.665 $Y=0.0675
c71 16 VSS 5.38922e-19 $X=0.557 $Y=0.0675
c72 11 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c73 6 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c74 1 VSS 5.38922e-19 $X=0.233 $Y=0.0675
r75 109 110 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.126 $X2=0.837 $Y2=0.144
r76 108 110 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.1495 $X2=0.837 $Y2=0.144
r77 106 108 5.12654 $w=1.8e-08 $l=7.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.1495
r78 105 109 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.045 $X2=0.837 $Y2=0.126
r79 103 104 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.8
+ $Y=0.234 $X2=0.814 $Y2=0.234
r80 101 103 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.8 $Y2=0.234
r81 98 101 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.756 $Y2=0.234
r82 95 98 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.648 $Y2=0.234
r83 92 95 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.54 $Y2=0.234
r84 89 92 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r85 85 89 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.324 $Y2=0.234
r86 83 106 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r87 83 104 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.814 $Y2=0.234
r88 81 82 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.8
+ $Y=0.036 $X2=0.814 $Y2=0.036
r89 79 81 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.8 $Y2=0.036
r90 79 80 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r91 76 79 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.756 $Y2=0.036
r92 76 77 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036 $X2=0.648
+ $Y2=0.036
r93 73 76 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.648 $Y2=0.036
r94 73 74 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r95 70 73 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.54 $Y2=0.036
r96 70 71 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r97 67 70 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r98 67 68 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r99 63 67 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.324 $Y2=0.036
r100 63 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r101 61 105 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.036 $X2=0.837 $Y2=0.045
r102 61 82 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.814 $Y2=0.036
r103 60 101 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234
+ $X2=0.756 $Y2=0.234
r104 57 60 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r105 56 60 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r106 55 98 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234
+ $X2=0.648 $Y2=0.234
r107 52 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.648 $Y2=0.2025
r108 51 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.648 $Y2=0.2025
r109 50 95 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r110 47 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r111 46 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r112 45 92 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r113 42 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r114 41 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r115 40 89 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r116 37 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r117 36 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r118 35 85 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r119 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r120 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r121 30 80 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.756 $Y=0.0675 $X2=0.756 $Y2=0.036
r122 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.756 $Y2=0.0675
r123 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.756 $Y2=0.0675
r124 25 77 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r125 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.648 $Y2=0.0675
r126 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0675 $X2=0.648 $Y2=0.0675
r127 20 74 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r128 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r129 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r130 15 71 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r131 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r132 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r133 10 68 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r134 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r135 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r136 5 64 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r137 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r138 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./BUFx12_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx12_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_4_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_4_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_4_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_4_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_4_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_4_M6_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_4_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_4_M8_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_4_M9_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 N_Y_M10_d N_4_M10_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M11 N_Y_M11_d N_4_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M12 N_Y_M12_d N_4_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M13 N_Y_M13_d N_4_M13_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.027
M14 N_4_M14_d N_A_M14_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M15 N_4_M15_d N_A_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M16 N_Y_M16_d N_4_M16_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M17 N_Y_M17_d N_4_M17_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M18 N_Y_M18_d N_4_M18_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M19 N_Y_M19_d N_4_M19_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M20 N_Y_M20_d N_4_M20_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M21 N_Y_M21_d N_4_M21_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M22 N_Y_M22_d N_4_M22_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M23 N_Y_M23_d N_4_M23_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M24 N_Y_M24_d N_4_M24_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M25 N_Y_M25_d N_4_M25_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
M26 N_Y_M26_d N_4_M26_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M27 N_Y_M27_d N_4_M27_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
*
* 
* .include "BUFx12_ASAP7_75t_SRAM.pex.sp.BUFX12_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx12_ASAP7_75t_SRAM.pex.sp.BUFX12_ASAP7_75T_SRAM.pxi"
* File: BUFx12_ASAP7_75t_SRAM.pex.sp.BUFX12_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:18:10 2017
* 
x_PM_BUFX12_ASAP7_75T_SRAM%A N_A_M0_g N_A_M14_g N_A_M1_g N_A_c_4_p N_A_M15_g A VSS
+ PM_BUFX12_ASAP7_75T_SRAM%A
x_PM_BUFX12_ASAP7_75T_SRAM%4 N_4_M2_g N_4_M16_g N_4_M3_g N_4_M17_g N_4_M4_g
+ N_4_M18_g N_4_M5_g N_4_M19_g N_4_M6_g N_4_M20_g N_4_M7_g N_4_M21_g N_4_M8_g
+ N_4_M22_g N_4_M9_g N_4_M23_g N_4_M10_g N_4_M24_g N_4_M11_g N_4_M25_g N_4_M12_g
+ N_4_M26_g N_4_M13_g N_4_c_25_n N_4_M27_g N_4_M1_d N_4_M0_d N_4_M15_d N_4_M14_d
+ N_4_c_28_n N_4_c_29_n N_4_c_32_n N_4_c_35_n N_4_c_67_p N_4_c_84_p N_4_c_36_n
+ N_4_c_68_p N_4_c_37_n N_4_c_82_p N_4_c_39_n N_4_c_41_n VSS
+ PM_BUFX12_ASAP7_75T_SRAM%4
x_PM_BUFX12_ASAP7_75T_SRAM%Y N_Y_M3_d N_Y_M2_d N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M6_d
+ N_Y_M9_d N_Y_M8_d N_Y_M11_d N_Y_M10_d N_Y_M13_d N_Y_M12_d N_Y_M17_d N_Y_M16_d
+ N_Y_M19_d N_Y_M18_d N_Y_M21_d N_Y_M20_d N_Y_M23_d N_Y_M22_d N_Y_M25_d
+ N_Y_M24_d N_Y_M27_d N_Y_M26_d N_Y_c_97_n N_Y_c_111_n Y N_Y_c_125_n VSS
+ PM_BUFX12_ASAP7_75T_SRAM%Y
cc_1 N_A_M0_g N_4_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_A_M1_g N_4_M2_g 0.00287079f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A_M1_g N_4_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_4 N_A_c_4_p N_4_c_25_n 0.00154931f $X=0.135 $Y=0.135 $X2=0.783 $Y2=0.135
cc_5 N_A_c_4_p N_4_M1_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_6 N_A_c_4_p N_4_M15_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_7 N_A_c_4_p N_4_c_28_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_8 N_A_M1_g N_4_c_29_n 6.45702e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.126
cc_9 N_A_c_4_p N_4_c_29_n 4.76064e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.126
cc_10 A N_4_c_29_n 6.94026e-19 $X=0.061 $Y=0.1325 $X2=0.135 $Y2=0.126
cc_11 N_A_M1_g N_4_c_32_n 6.45702e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.225
cc_12 N_A_c_4_p N_4_c_32_n 4.76064e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.225
cc_13 A N_4_c_32_n 6.94026e-19 $X=0.061 $Y=0.1325 $X2=0.135 $Y2=0.225
cc_14 N_A_c_4_p N_4_c_35_n 4.61514e-19 $X=0.135 $Y=0.135 $X2=0.199 $Y2=0.135
cc_15 N_A_c_4_p N_4_c_36_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.036
cc_16 N_A_c_4_p N_4_c_37_n 3.38382e-19 $X=0.135 $Y=0.135 $X2=0.126 $Y2=0.036
cc_17 A N_4_c_37_n 5.11982e-19 $X=0.061 $Y=0.1325 $X2=0.126 $Y2=0.036
cc_18 N_A_c_4_p N_4_c_39_n 3.38382e-19 $X=0.135 $Y=0.135 $X2=0.126 $Y2=0.234
cc_19 A N_4_c_39_n 5.11982e-19 $X=0.061 $Y=0.1325 $X2=0.126 $Y2=0.234
cc_20 N_A_c_4_p N_4_c_41_n 0.00117248f $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.135
cc_21 A N_4_c_41_n 5.86795e-19 $X=0.061 $Y=0.1325 $X2=0.135 $Y2=0.135
cc_22 N_4_c_25_n N_Y_M3_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_23 N_4_c_25_n N_Y_M5_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_24 N_4_c_25_n N_Y_M7_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_25 N_4_c_25_n N_Y_M9_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_26 N_4_c_25_n N_Y_M11_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_27 N_4_c_25_n N_Y_M13_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0.064 $Y2=0.135
cc_28 N_4_c_25_n N_Y_M17_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_29 N_4_c_25_n N_Y_M19_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0.081 $Y2=0.135
cc_30 N_4_c_25_n N_Y_M21_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_31 N_4_c_25_n N_Y_M23_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_32 N_4_c_25_n N_Y_M25_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_33 N_4_c_25_n N_Y_M27_d 3.80218e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_34 N_4_M3_g N_Y_c_97_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_4_M4_g N_Y_c_97_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_4_M5_g N_Y_c_97_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_4_M6_g N_Y_c_97_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_38 N_4_M7_g N_Y_c_97_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_4_M8_g N_Y_c_97_n 4.28653e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_40 N_4_M9_g N_Y_c_97_n 4.28653e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_41 N_4_M10_g N_Y_c_97_n 4.28653e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_42 N_4_M11_g N_Y_c_97_n 4.28653e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_4_M12_g N_Y_c_97_n 4.28653e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_4_M13_g N_Y_c_97_n 4.28653e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_45 N_4_c_25_n N_Y_c_97_n 0.00222875f $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_67_p N_Y_c_97_n 0.00813322f $X=0.221 $Y=0.135 $X2=0 $Y2=0
cc_47 N_4_c_68_p N_Y_c_97_n 3.91654e-19 $X=0.135 $Y=0.036 $X2=0 $Y2=0
cc_48 N_4_M3_g N_Y_c_111_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_49 N_4_M4_g N_Y_c_111_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_50 N_4_M5_g N_Y_c_111_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_51 N_4_M6_g N_Y_c_111_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_52 N_4_M7_g N_Y_c_111_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_53 N_4_M8_g N_Y_c_111_n 4.28653e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_54 N_4_M9_g N_Y_c_111_n 4.28653e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_55 N_4_M10_g N_Y_c_111_n 4.28653e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_56 N_4_M11_g N_Y_c_111_n 4.28653e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_57 N_4_M12_g N_Y_c_111_n 4.28653e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_4_M13_g N_Y_c_111_n 4.28653e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_59 N_4_c_25_n N_Y_c_111_n 0.00222875f $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_60 N_4_c_67_p N_Y_c_111_n 0.00813322f $X=0.221 $Y=0.135 $X2=0 $Y2=0
cc_61 N_4_c_82_p N_Y_c_111_n 3.91654e-19 $X=0.135 $Y=0.234 $X2=0 $Y2=0
cc_62 N_4_c_25_n N_Y_c_125_n 5.11403e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_63 N_4_c_84_p N_Y_c_125_n 0.00113063f $X=0.729 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx12_ASAP7_75t_SRAM.pex.sp.BUFX12_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx12f_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:18:32 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx12f_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx12f_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx12f_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:18:32 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX12F_ASAP7_75T_SRAM%A 2 7 10 15 18 23 26 29 31 34 VSS
c24 34 VSS 0.00762485f $X=0.064 $Y=0.135
c25 29 VSS 0.0195581f $X=0.243 $Y=0.135
c26 26 VSS 0.061051f $X=0.243 $Y=0.0675
c27 18 VSS 0.0642127f $X=0.189 $Y=0.0675
c28 10 VSS 0.0644226f $X=0.135 $Y=0.0675
c29 2 VSS 0.0656042f $X=0.081 $Y=0.0675
r30 34 37 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r31 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r32 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r33 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r34 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r35 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r36 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r37 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r38 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r39 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r40 5 37 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r41 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r42 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX12F_ASAP7_75T_SRAM%4 2 7 10 15 18 23 26 31 34 39 42 47 50 55 58 63
+ 66 71 74 79 82 87 90 93 95 97 98 102 103 107 108 111 112 113 116 117 120 124
+ 125 134 136 VSS
c75 147 VSS 4.77902e-19 $X=0.288 $Y=0.135
c76 146 VSS 5.7781e-20 $X=0.279 $Y=0.135
c77 144 VSS 6.48584e-19 $X=0.297 $Y=0.135
c78 140 VSS 3.90656e-19 $X=0.27 $Y=0.214
c79 139 VSS 0.00327153f $X=0.27 $Y=0.203
c80 138 VSS 3.65892e-19 $X=0.27 $Y=0.225
c81 136 VSS 0.00133736f $X=0.27 $Y=0.0965
c82 135 VSS 7.56089e-19 $X=0.27 $Y=0.067
c83 134 VSS 0.00193417f $X=0.27 $Y=0.126
c84 125 VSS 0.0222181f $X=0.261 $Y=0.234
c85 124 VSS 0.00939167f $X=0.216 $Y=0.036
c86 120 VSS 0.00947391f $X=0.108 $Y=0.036
c87 117 VSS 0.0222181f $X=0.261 $Y=0.036
c88 116 VSS 0.00939167f $X=0.216 $Y=0.2025
c89 112 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c90 111 VSS 0.00947391f $X=0.108 $Y=0.2025
c91 107 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c92 102 VSS 5.38922e-19 $X=0.233 $Y=0.0675
c93 97 VSS 5.72268e-19 $X=0.125 $Y=0.0675
c94 93 VSS 0.0553909f $X=0.891 $Y=0.135
c95 90 VSS 0.0645347f $X=0.891 $Y=0.0675
c96 82 VSS 0.0644226f $X=0.837 $Y=0.0675
c97 74 VSS 0.0642127f $X=0.783 $Y=0.0675
c98 66 VSS 0.0642127f $X=0.729 $Y=0.0675
c99 58 VSS 0.0642127f $X=0.675 $Y=0.0675
c100 50 VSS 0.0642127f $X=0.621 $Y=0.0675
c101 42 VSS 0.0642127f $X=0.567 $Y=0.0675
c102 34 VSS 0.0642127f $X=0.513 $Y=0.0675
c103 26 VSS 0.0642127f $X=0.459 $Y=0.0675
c104 18 VSS 0.0642127f $X=0.405 $Y=0.0675
c105 10 VSS 0.0642127f $X=0.351 $Y=0.0675
c106 2 VSS 0.0616955f $X=0.297 $Y=0.0675
r107 146 147 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.135 $X2=0.288 $Y2=0.135
r108 144 147 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.288 $Y2=0.135
r109 141 146 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.135 $X2=0.279 $Y2=0.135
r110 139 140 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.203 $X2=0.27 $Y2=0.214
r111 138 140 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.225 $X2=0.27 $Y2=0.214
r112 137 141 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.144 $X2=0.27 $Y2=0.135
r113 137 139 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.144 $X2=0.27 $Y2=0.203
r114 135 136 2.00309 $w=1.8e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.067 $X2=0.27 $Y2=0.0965
r115 134 141 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.126 $X2=0.27 $Y2=0.135
r116 134 136 2.00309 $w=1.8e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.126 $X2=0.27 $Y2=0.0965
r117 133 135 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.045 $X2=0.27 $Y2=0.067
r118 127 131 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.108 $Y=0.234 $X2=0.216 $Y2=0.234
r119 125 138 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.261 $Y=0.234 $X2=0.27 $Y2=0.225
r120 125 131 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.234 $X2=0.216 $Y2=0.234
r121 123 124 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r122 119 123 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.108 $Y=0.036 $X2=0.216 $Y2=0.036
r123 119 120 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r124 117 133 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.261 $Y=0.036 $X2=0.27 $Y2=0.045
r125 117 123 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.036 $X2=0.216 $Y2=0.036
r126 116 131 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r127 113 116 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r128 112 116 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r129 111 127 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r130 108 111 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r131 107 111 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r132 106 124 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.216 $Y=0.0675 $X2=0.216 $Y2=0.036
r133 103 106 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r134 102 106 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r135 101 120 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.108 $Y=0.0675 $X2=0.108 $Y2=0.036
r136 98 101 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r137 97 101 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r138 93 95 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.135 $X2=0.891 $Y2=0.2025
r139 90 93 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.0675 $X2=0.891 $Y2=0.135
r140 85 93 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.837
+ $Y=0.135 $X2=0.891 $Y2=0.135
r141 85 87 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.135 $X2=0.837 $Y2=0.2025
r142 82 85 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0675 $X2=0.837 $Y2=0.135
r143 77 85 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.783
+ $Y=0.135 $X2=0.837 $Y2=0.135
r144 77 79 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.135 $X2=0.783 $Y2=0.2025
r145 74 77 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.135
r146 69 77 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.135 $X2=0.783 $Y2=0.135
r147 69 71 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.135 $X2=0.729 $Y2=0.2025
r148 66 69 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.135
r149 61 69 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.729 $Y2=0.135
r150 61 63 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2025
r151 58 61 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0675 $X2=0.675 $Y2=0.135
r152 53 61 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621
+ $Y=0.135 $X2=0.675 $Y2=0.135
r153 53 55 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2025
r154 50 53 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r155 45 53 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.567
+ $Y=0.135 $X2=0.621 $Y2=0.135
r156 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.135 $X2=0.567 $Y2=0.2025
r157 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.0675 $X2=0.567 $Y2=0.135
r158 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r159 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r160 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r161 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r162 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r163 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r164 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r165 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r166 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r167 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r168 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r169 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r170 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r171 5 144 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r172 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r173 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_BUFX12F_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 21 22 26 27 31 32 35 36 37
+ 40 41 42 45 46 47 50 51 52 55 56 57 60 61 63 64 70 73 76 79 82 83 85 108 VSS
c51 108 VSS 0.0113708f $X=0.945 $Y=0.132
c52 85 VSS 0.00124235f $X=0.324 $Y=0.234
c53 83 VSS 0.0736356f $X=0.936 $Y=0.234
c54 82 VSS 0.00929752f $X=0.864 $Y=0.036
c55 79 VSS 0.00928953f $X=0.756 $Y=0.036
c56 76 VSS 0.00928955f $X=0.648 $Y=0.036
c57 73 VSS 0.00928955f $X=0.54 $Y=0.036
c58 70 VSS 0.00928943f $X=0.432 $Y=0.036
c59 64 VSS 0.00908821f $X=0.324 $Y=0.036
c60 63 VSS 0.00124235f $X=0.324 $Y=0.036
c61 61 VSS 0.0736356f $X=0.936 $Y=0.036
c62 60 VSS 0.00929752f $X=0.864 $Y=0.2025
c63 56 VSS 5.38922e-19 $X=0.881 $Y=0.2025
c64 55 VSS 0.00928953f $X=0.756 $Y=0.2025
c65 51 VSS 5.38922e-19 $X=0.773 $Y=0.2025
c66 50 VSS 0.00928955f $X=0.648 $Y=0.2025
c67 46 VSS 5.38922e-19 $X=0.665 $Y=0.2025
c68 45 VSS 0.00928955f $X=0.54 $Y=0.2025
c69 41 VSS 5.38922e-19 $X=0.557 $Y=0.2025
c70 40 VSS 0.00928943f $X=0.432 $Y=0.2025
c71 36 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c72 35 VSS 0.00908821f $X=0.324 $Y=0.2025
c73 31 VSS 5.58795e-19 $X=0.341 $Y=0.2025
c74 26 VSS 5.38922e-19 $X=0.881 $Y=0.0675
c75 21 VSS 5.38922e-19 $X=0.773 $Y=0.0675
c76 16 VSS 5.38922e-19 $X=0.665 $Y=0.0675
c77 11 VSS 5.38922e-19 $X=0.557 $Y=0.0675
c78 6 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c79 1 VSS 5.58795e-19 $X=0.341 $Y=0.0675
r80 106 108 6.31482 $w=1.8e-08 $l=9.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.225 $X2=0.945 $Y2=0.132
r81 105 108 5.90741 $w=1.8e-08 $l=8.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.945
+ $Y=0.045 $X2=0.945 $Y2=0.132
r82 100 103 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.864 $Y2=0.234
r83 97 100 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.756 $Y2=0.234
r84 94 97 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.648 $Y2=0.234
r85 91 94 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.54 $Y2=0.234
r86 85 91 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r87 83 106 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.234 $X2=0.945 $Y2=0.225
r88 83 103 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.234 $X2=0.864 $Y2=0.234
r89 81 82 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036 $X2=0.864
+ $Y2=0.036
r90 78 81 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.864 $Y2=0.036
r91 78 79 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r92 75 78 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.756 $Y2=0.036
r93 75 76 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036 $X2=0.648
+ $Y2=0.036
r94 72 75 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.648 $Y2=0.036
r95 72 73 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r96 69 72 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.54 $Y2=0.036
r97 69 70 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r98 63 69 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r99 63 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r100 61 105 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.936 $Y=0.036 $X2=0.945 $Y2=0.045
r101 61 81 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.936
+ $Y=0.036 $X2=0.864 $Y2=0.036
r102 60 103 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234
+ $X2=0.864 $Y2=0.234
r103 57 60 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2025 $X2=0.864 $Y2=0.2025
r104 56 60 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2025 $X2=0.864 $Y2=0.2025
r105 55 100 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234
+ $X2=0.756 $Y2=0.234
r106 52 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r107 51 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r108 50 97 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234
+ $X2=0.648 $Y2=0.234
r109 47 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.648 $Y2=0.2025
r110 46 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.648 $Y2=0.2025
r111 45 94 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r112 42 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r113 41 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r114 40 91 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r115 37 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r116 36 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r117 35 85 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r118 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r119 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r120 30 82 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.864 $Y=0.0675 $X2=0.864 $Y2=0.036
r121 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0675 $X2=0.864 $Y2=0.0675
r122 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0675 $X2=0.864 $Y2=0.0675
r123 25 79 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.756 $Y=0.0675 $X2=0.756 $Y2=0.036
r124 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.756 $Y2=0.0675
r125 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.756 $Y2=0.0675
r126 20 76 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r127 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.648 $Y2=0.0675
r128 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0675 $X2=0.648 $Y2=0.0675
r129 15 73 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r130 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r131 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r132 10 70 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r133 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r134 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r135 5 64 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r136 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r137 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
.ends


* END of "./BUFx12f_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx12f_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_4_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_4_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_4_M2_d N_A_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_4_M3_d N_A_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_4_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_4_M6_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_4_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_4_M8_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_4_M9_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 N_Y_M10_d N_4_M10_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M11 N_Y_M11_d N_4_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M12 N_Y_M12_d N_4_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M13 N_Y_M13_d N_4_M13_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.027
M14 N_Y_M14_d N_4_M14_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.027
M15 N_Y_M15_d N_4_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.027
M16 N_4_M16_d N_A_M16_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M17 N_4_M17_d N_A_M17_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M18 N_4_M18_d N_A_M18_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M19 N_4_M19_d N_A_M19_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M20 N_Y_M20_d N_4_M20_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M21 N_Y_M21_d N_4_M21_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M22 N_Y_M22_d N_4_M22_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M23 N_Y_M23_d N_4_M23_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M24 N_Y_M24_d N_4_M24_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M25 N_Y_M25_d N_4_M25_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M26 N_Y_M26_d N_4_M26_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M27 N_Y_M27_d N_4_M27_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
M28 N_Y_M28_d N_4_M28_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M29 N_Y_M29_d N_4_M29_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
M30 N_Y_M30_d N_4_M30_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.162
M31 N_Y_M31_d N_4_M31_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.162
*
* 
* .include "BUFx12f_ASAP7_75t_SRAM.pex.sp.BUFX12F_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx12f_ASAP7_75t_SRAM.pex.sp.BUFX12F_ASAP7_75T_SRAM.pxi"
* File: BUFx12f_ASAP7_75t_SRAM.pex.sp.BUFX12F_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:18:32 2017
* 
x_PM_BUFX12F_ASAP7_75T_SRAM%A N_A_M0_g N_A_M16_g N_A_M1_g N_A_M17_g N_A_M2_g
+ N_A_M18_g N_A_M3_g N_A_c_4_p N_A_M19_g A VSS PM_BUFX12F_ASAP7_75T_SRAM%A
x_PM_BUFX12F_ASAP7_75T_SRAM%4 N_4_M4_g N_4_M20_g N_4_M5_g N_4_M21_g N_4_M6_g
+ N_4_M22_g N_4_M7_g N_4_M23_g N_4_M8_g N_4_M24_g N_4_M9_g N_4_M25_g N_4_M10_g
+ N_4_M26_g N_4_M11_g N_4_M27_g N_4_M12_g N_4_M28_g N_4_M13_g N_4_M29_g
+ N_4_M14_g N_4_M30_g N_4_M15_g N_4_c_28_n N_4_M31_g N_4_M1_d N_4_M0_d N_4_M3_d
+ N_4_M2_d N_4_M17_d N_4_M16_d N_4_c_32_n N_4_M19_d N_4_M18_d N_4_c_35_n
+ N_4_c_36_n N_4_c_40_n N_4_c_42_n N_4_c_43_n N_4_c_47_n N_4_c_48_n VSS
+ PM_BUFX12F_ASAP7_75T_SRAM%4
x_PM_BUFX12F_ASAP7_75T_SRAM%Y N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M6_d N_Y_M9_d N_Y_M8_d
+ N_Y_M11_d N_Y_M10_d N_Y_M13_d N_Y_M12_d N_Y_M15_d N_Y_M14_d N_Y_M21_d
+ N_Y_M20_d N_Y_c_107_n N_Y_M23_d N_Y_M22_d N_Y_c_109_n N_Y_M25_d N_Y_M24_d
+ N_Y_c_111_n N_Y_M27_d N_Y_M26_d N_Y_c_113_n N_Y_M29_d N_Y_M28_d N_Y_c_115_n
+ N_Y_M31_d N_Y_M30_d N_Y_c_117_n N_Y_c_118_n N_Y_c_129_n N_Y_c_131_n
+ N_Y_c_132_n N_Y_c_133_n N_Y_c_134_n N_Y_c_135_n N_Y_c_136_n N_Y_c_137_n
+ N_Y_c_148_n Y VSS PM_BUFX12F_ASAP7_75T_SRAM%Y
cc_1 N_A_M2_g N_4_M4_g 2.34385e-19 $X=0.189 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_2 N_A_M3_g N_4_M4_g 0.00287079f $X=0.243 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_3 N_A_M3_g N_4_M5_g 2.34385e-19 $X=0.243 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_4 N_A_c_4_p N_4_c_28_n 0.00109521f $X=0.243 $Y=0.135 $X2=0.891 $Y2=0.135
cc_5 N_A_c_4_p N_4_M1_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_6 N_A_c_4_p N_4_M3_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.233 $Y2=0.0675
cc_7 N_A_c_4_p N_4_M17_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_8 N_A_c_4_p N_4_c_32_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_9 A N_4_c_32_n 0.00116725f $X=0.064 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_10 N_A_c_4_p N_4_M19_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.233 $Y2=0.2025
cc_11 N_A_c_4_p N_4_c_35_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.216 $Y2=0.2025
cc_12 N_A_M1_g N_4_c_36_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.261 $Y2=0.036
cc_13 N_A_M2_g N_4_c_36_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.261 $Y2=0.036
cc_14 N_A_M3_g N_4_c_36_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.261 $Y2=0.036
cc_15 N_A_c_4_p N_4_c_36_n 0.00189731f $X=0.243 $Y=0.135 $X2=0.261 $Y2=0.036
cc_16 N_A_c_4_p N_4_c_40_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.108 $Y2=0.036
cc_17 A N_4_c_40_n 0.00116725f $X=0.064 $Y=0.135 $X2=0.108 $Y2=0.036
cc_18 N_A_c_4_p N_4_c_42_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.216 $Y2=0.036
cc_19 N_A_M1_g N_4_c_43_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.261 $Y2=0.234
cc_20 N_A_M2_g N_4_c_43_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.261 $Y2=0.234
cc_21 N_A_M3_g N_4_c_43_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.261 $Y2=0.234
cc_22 N_A_c_4_p N_4_c_43_n 0.00189731f $X=0.243 $Y=0.135 $X2=0.261 $Y2=0.234
cc_23 N_A_c_4_p N_4_c_47_n 3.90981e-19 $X=0.243 $Y=0.135 $X2=0.27 $Y2=0.126
cc_24 A N_4_c_48_n 6.51825e-19 $X=0.064 $Y=0.135 $X2=0.27 $Y2=0.0965
cc_25 N_4_c_28_n N_Y_M5_d 3.80485e-19 $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_26 N_4_c_28_n N_Y_M7_d 3.80663e-19 $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_27 N_4_c_28_n N_Y_M9_d 3.80663e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_28 N_4_c_28_n N_Y_M11_d 3.80663e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_29 N_4_c_28_n N_Y_M13_d 3.80663e-19 $X=0.891 $Y=0.135 $X2=0.189 $Y2=0.135
cc_30 N_4_c_28_n N_Y_M15_d 3.80663e-19 $X=0.891 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_31 N_4_c_28_n N_Y_M21_d 3.80485e-19 $X=0.891 $Y=0.135 $X2=0.243 $Y2=0.2025
cc_32 N_4_c_28_n N_Y_c_107_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_33 N_4_c_28_n N_Y_M23_d 3.80663e-19 $X=0.891 $Y=0.135 $X2=0.064 $Y2=0.135
cc_34 N_4_c_28_n N_Y_c_109_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_35 N_4_c_28_n N_Y_M25_d 3.80663e-19 $X=0.891 $Y=0.135 $X2=0.081 $Y2=0.135
cc_36 N_4_c_28_n N_Y_c_111_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_28_n N_Y_M27_d 3.80663e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_28_n N_Y_c_113_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_39 N_4_c_28_n N_Y_M29_d 3.80663e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_28_n N_Y_c_115_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_41 N_4_c_28_n N_Y_M31_d 3.80663e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_42 N_4_c_28_n N_Y_c_117_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_43 N_4_M5_g N_Y_c_118_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_4_M6_g N_Y_c_118_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_45 N_4_M7_g N_Y_c_118_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_46 N_4_M8_g N_Y_c_118_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_4_M9_g N_Y_c_118_n 4.59284e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_48 N_4_M10_g N_Y_c_118_n 4.59284e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_49 N_4_M11_g N_Y_c_118_n 4.59284e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_50 N_4_M12_g N_Y_c_118_n 4.59284e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_51 N_4_M13_g N_Y_c_118_n 4.59284e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_52 N_4_M14_g N_Y_c_118_n 4.59284e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_53 N_4_M15_g N_Y_c_118_n 4.59284e-19 $X=0.891 $Y=0.0675 $X2=0 $Y2=0
cc_54 N_4_c_28_n N_Y_c_129_n 0.00738027f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_55 N_4_c_36_n N_Y_c_129_n 0.00106268f $X=0.261 $Y=0.036 $X2=0 $Y2=0
cc_56 N_4_c_28_n N_Y_c_131_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_57 N_4_c_28_n N_Y_c_132_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_58 N_4_c_28_n N_Y_c_133_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_59 N_4_c_28_n N_Y_c_134_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_60 N_4_c_28_n N_Y_c_135_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_61 N_4_c_28_n N_Y_c_136_n 8.00061e-19 $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_62 N_4_M5_g N_Y_c_137_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_63 N_4_M6_g N_Y_c_137_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_4_M7_g N_Y_c_137_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_65 N_4_M8_g N_Y_c_137_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_66 N_4_M9_g N_Y_c_137_n 4.59284e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_67 N_4_M10_g N_Y_c_137_n 4.59284e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_68 N_4_M11_g N_Y_c_137_n 4.59284e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_69 N_4_M12_g N_Y_c_137_n 4.59284e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_70 N_4_M13_g N_Y_c_137_n 4.59284e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_71 N_4_M14_g N_Y_c_137_n 4.59284e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_72 N_4_M15_g N_Y_c_137_n 4.59284e-19 $X=0.891 $Y=0.0675 $X2=0 $Y2=0
cc_73 N_4_c_28_n N_Y_c_148_n 0.00738027f $X=0.891 $Y=0.135 $X2=0 $Y2=0
cc_74 N_4_c_43_n N_Y_c_148_n 0.00106268f $X=0.261 $Y=0.234 $X2=0 $Y2=0
cc_75 N_4_c_28_n Y 0.00104674f $X=0.891 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx12f_ASAP7_75t_SRAM.pex.sp.BUFX12F_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx16f_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:18:54 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx16f_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx16f_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx16f_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:18:54 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX16F_ASAP7_75T_SRAM%A 2 7 10 15 18 23 26 29 31 34 38 VSS
c28 34 VSS 0.00760081f $X=0.064 $Y=0.135
c29 29 VSS 0.0198635f $X=0.243 $Y=0.135
c30 26 VSS 0.0609945f $X=0.243 $Y=0.0675
c31 18 VSS 0.0642127f $X=0.189 $Y=0.0675
c32 10 VSS 0.0644226f $X=0.135 $Y=0.0675
c33 2 VSS 0.0656042f $X=0.081 $Y=0.0675
r34 34 38 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.135 $X2=0.064 $Y2=0.1495
r35 34 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r36 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r37 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r38 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r39 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r40 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r41 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r42 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r43 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r44 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r45 5 35 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r46 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r47 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX16F_ASAP7_75T_SRAM%4 2 7 10 15 18 23 26 31 34 39 42 47 50 55 58 63
+ 66 71 74 79 82 87 90 95 98 103 106 111 114 119 122 125 127 129 130 134 135 139
+ 140 143 144 145 148 149 152 156 157 166 168 171 177 178 192 195 VSS
c82 195 VSS 2.15872e-20 $X=0.243 $Y=0.135
c83 192 VSS 3.38107e-19 $X=1.107 $Y=0.135
c84 177 VSS 0.00280817f $X=0.31 $Y=0.135
c85 172 VSS 5.69453e-19 $X=0.243 $Y=0.214
c86 171 VSS 0.00250569f $X=0.243 $Y=0.203
c87 170 VSS 5.5755e-19 $X=0.243 $Y=0.225
c88 168 VSS 0.00142491f $X=0.243 $Y=0.0965
c89 167 VSS 0.00112792f $X=0.243 $Y=0.067
c90 166 VSS 0.00108079f $X=0.243 $Y=0.126
c91 157 VSS 0.0190647f $X=0.234 $Y=0.234
c92 156 VSS 0.0104726f $X=0.216 $Y=0.036
c93 152 VSS 0.0094735f $X=0.108 $Y=0.036
c94 149 VSS 0.0190647f $X=0.234 $Y=0.036
c95 148 VSS 0.0104726f $X=0.216 $Y=0.2025
c96 144 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c97 143 VSS 0.0094735f $X=0.108 $Y=0.2025
c98 139 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c99 134 VSS 5.38922e-19 $X=0.233 $Y=0.0675
c100 129 VSS 5.72268e-19 $X=0.125 $Y=0.0675
c101 125 VSS 0.0544265f $X=1.107 $Y=0.135
c102 122 VSS 0.0645347f $X=1.107 $Y=0.0675
c103 114 VSS 0.0644226f $X=1.053 $Y=0.0675
c104 106 VSS 0.0642127f $X=0.999 $Y=0.0675
c105 98 VSS 0.0642127f $X=0.945 $Y=0.0675
c106 90 VSS 0.0642127f $X=0.891 $Y=0.0675
c107 82 VSS 0.0642127f $X=0.837 $Y=0.0675
c108 74 VSS 0.0642127f $X=0.783 $Y=0.0675
c109 66 VSS 0.0642127f $X=0.729 $Y=0.0675
c110 58 VSS 0.0642127f $X=0.675 $Y=0.0675
c111 50 VSS 0.0642127f $X=0.621 $Y=0.0675
c112 42 VSS 0.0642127f $X=0.567 $Y=0.0675
c113 34 VSS 0.0642127f $X=0.513 $Y=0.0675
c114 26 VSS 0.0642127f $X=0.459 $Y=0.0675
c115 18 VSS 0.0642127f $X=0.405 $Y=0.0675
c116 10 VSS 0.0642127f $X=0.351 $Y=0.0675
c117 2 VSS 0.0616955f $X=0.297 $Y=0.0675
r118 189 192 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.999 $Y=0.135 $X2=1.107 $Y2=0.135
r119 186 189 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.135 $X2=0.999 $Y2=0.135
r120 183 186 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.135 $X2=0.837 $Y2=0.135
r121 180 183 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.675 $Y2=0.135
r122 177 178 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.31
+ $Y=0.135 $X2=0.3305 $Y2=0.135
r123 175 180 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.513 $Y2=0.135
r124 175 178 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.351 $Y=0.135 $X2=0.3305 $Y2=0.135
r125 173 195 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.243 $Y2=0.135
r126 173 177 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.31 $Y2=0.135
r127 171 172 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.243 $Y=0.203 $X2=0.243 $Y2=0.214
r128 170 172 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.243 $Y=0.225 $X2=0.243 $Y2=0.214
r129 169 195 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.144 $X2=0.243 $Y2=0.135
r130 169 171 4.00617 $w=1.8e-08 $l=5.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.144 $X2=0.243 $Y2=0.203
r131 167 168 2.00309 $w=1.8e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.243 $Y=0.067 $X2=0.243 $Y2=0.0965
r132 166 195 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.135
r133 166 168 2.00309 $w=1.8e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.243 $Y=0.126 $X2=0.243 $Y2=0.0965
r134 165 167 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.067
r135 159 163 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.108 $Y=0.234 $X2=0.216 $Y2=0.234
r136 157 170 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r137 157 163 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r138 155 156 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r139 151 155 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.108 $Y=0.036 $X2=0.216 $Y2=0.036
r140 151 152 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r141 149 165 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r142 149 155 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r143 148 163 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r144 145 148 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r145 144 148 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r146 143 159 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r147 140 143 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r148 139 143 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r149 138 156 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.216 $Y=0.0675 $X2=0.216 $Y2=0.036
r150 135 138 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r151 134 138 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r152 133 152 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.108 $Y=0.0675 $X2=0.108 $Y2=0.036
r153 130 133 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r154 129 133 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r155 125 192 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=1.107 $Y=0.135
+ $X2=1.107 $Y2=0.135
r156 125 127 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.135 $X2=1.107 $Y2=0.2025
r157 122 125 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.0675 $X2=1.107 $Y2=0.135
r158 117 125 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.053
+ $Y=0.135 $X2=1.107 $Y2=0.135
r159 117 119 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.135 $X2=1.053 $Y2=0.2025
r160 114 117 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.0675 $X2=1.053 $Y2=0.135
r161 109 117 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.999
+ $Y=0.135 $X2=1.053 $Y2=0.135
r162 109 189 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.999 $Y=0.135
+ $X2=0.999 $Y2=0.135
r163 109 111 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.135 $X2=0.999 $Y2=0.2025
r164 106 109 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.135
r165 101 109 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.945
+ $Y=0.135 $X2=0.999 $Y2=0.135
r166 101 103 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.135 $X2=0.945 $Y2=0.2025
r167 98 101 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.0675 $X2=0.945 $Y2=0.135
r168 93 101 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.891
+ $Y=0.135 $X2=0.945 $Y2=0.135
r169 93 95 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.135 $X2=0.891 $Y2=0.2025
r170 90 93 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.0675 $X2=0.891 $Y2=0.135
r171 85 93 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.837
+ $Y=0.135 $X2=0.891 $Y2=0.135
r172 85 186 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.837 $Y=0.135
+ $X2=0.837 $Y2=0.135
r173 85 87 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.135 $X2=0.837 $Y2=0.2025
r174 82 85 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0675 $X2=0.837 $Y2=0.135
r175 77 85 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.783
+ $Y=0.135 $X2=0.837 $Y2=0.135
r176 77 79 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.135 $X2=0.783 $Y2=0.2025
r177 74 77 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.135
r178 69 77 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.135 $X2=0.783 $Y2=0.135
r179 69 71 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.135 $X2=0.729 $Y2=0.2025
r180 66 69 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.135
r181 61 69 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.729 $Y2=0.135
r182 61 183 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.675 $Y=0.135
+ $X2=0.675 $Y2=0.135
r183 61 63 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2025
r184 58 61 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0675 $X2=0.675 $Y2=0.135
r185 53 61 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621
+ $Y=0.135 $X2=0.675 $Y2=0.135
r186 53 55 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2025
r187 50 53 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r188 45 53 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.567
+ $Y=0.135 $X2=0.621 $Y2=0.135
r189 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.135 $X2=0.567 $Y2=0.2025
r190 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.0675 $X2=0.567 $Y2=0.135
r191 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r192 37 180 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.513 $Y=0.135
+ $X2=0.513 $Y2=0.135
r193 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r194 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r195 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r196 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r197 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r198 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r199 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r200 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r201 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r202 13 175 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.351 $Y=0.135
+ $X2=0.351 $Y2=0.135
r203 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r204 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r205 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r206 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r207 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_BUFX16F_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 21 22 26 27 31 32 36 37 41
+ 42 46 47 51 52 56 57 61 62 66 67 71 72 76 77 107 135 140 142 VSS
c54 142 VSS 7.43984e-19 $X=1.161 $Y=0.144
c55 141 VSS 0.00538269f $X=1.161 $Y=0.126
c56 140 VSS 0.00538269f $X=1.16 $Y=0.1495
c57 136 VSS 0.00237022f $X=1.138 $Y=0.234
c58 135 VSS 0.0867056f $X=1.124 $Y=0.234
c59 109 VSS 0.00566127f $X=1.152 $Y=0.234
c60 108 VSS 0.00237022f $X=1.138 $Y=0.036
c61 107 VSS 0.0867056f $X=1.124 $Y=0.036
c62 106 VSS 0.00929752f $X=1.08 $Y=0.036
c63 103 VSS 0.00928953f $X=0.972 $Y=0.036
c64 100 VSS 0.00928955f $X=0.864 $Y=0.036
c65 97 VSS 0.00928955f $X=0.756 $Y=0.036
c66 94 VSS 0.00928955f $X=0.648 $Y=0.036
c67 91 VSS 0.00928955f $X=0.54 $Y=0.036
c68 88 VSS 0.00928953f $X=0.432 $Y=0.036
c69 84 VSS 0.00917567f $X=0.324 $Y=0.036
c70 81 VSS 0.00566127f $X=1.152 $Y=0.036
c71 80 VSS 0.00929752f $X=1.08 $Y=0.2025
c72 76 VSS 5.38922e-19 $X=1.097 $Y=0.2025
c73 75 VSS 0.00928953f $X=0.972 $Y=0.2025
c74 71 VSS 5.38922e-19 $X=0.989 $Y=0.2025
c75 70 VSS 0.00928955f $X=0.864 $Y=0.2025
c76 66 VSS 5.38922e-19 $X=0.881 $Y=0.2025
c77 65 VSS 0.00928955f $X=0.756 $Y=0.2025
c78 61 VSS 5.38922e-19 $X=0.773 $Y=0.2025
c79 60 VSS 0.00928955f $X=0.648 $Y=0.2025
c80 56 VSS 5.38922e-19 $X=0.665 $Y=0.2025
c81 55 VSS 0.00928955f $X=0.54 $Y=0.2025
c82 51 VSS 5.38922e-19 $X=0.557 $Y=0.2025
c83 50 VSS 0.00928953f $X=0.432 $Y=0.2025
c84 46 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c85 45 VSS 0.00917567f $X=0.324 $Y=0.2025
c86 41 VSS 5.72268e-19 $X=0.341 $Y=0.2025
c87 36 VSS 5.38922e-19 $X=1.097 $Y=0.0675
c88 31 VSS 5.38922e-19 $X=0.989 $Y=0.0675
c89 26 VSS 5.38922e-19 $X=0.881 $Y=0.0675
c90 21 VSS 5.38922e-19 $X=0.773 $Y=0.0675
c91 16 VSS 5.38922e-19 $X=0.665 $Y=0.0675
c92 11 VSS 5.38922e-19 $X=0.557 $Y=0.0675
c93 6 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c94 1 VSS 5.72268e-19 $X=0.341 $Y=0.0675
r95 141 142 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.126 $X2=1.161 $Y2=0.144
r96 140 142 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.1495 $X2=1.161 $Y2=0.144
r97 138 140 5.12654 $w=1.8e-08 $l=7.55e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.225 $X2=1.161 $Y2=0.1495
r98 137 141 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.045 $X2=1.161 $Y2=0.126
r99 135 136 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.124
+ $Y=0.234 $X2=1.138 $Y2=0.234
r100 133 135 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.124 $Y2=0.234
r101 130 133 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.972 $Y=0.234 $X2=1.08 $Y2=0.234
r102 127 130 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.864 $Y=0.234 $X2=0.972 $Y2=0.234
r103 124 127 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.756 $Y=0.234 $X2=0.864 $Y2=0.234
r104 121 124 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.648 $Y=0.234 $X2=0.756 $Y2=0.234
r105 118 121 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.648 $Y2=0.234
r106 115 118 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.432 $Y=0.234 $X2=0.54 $Y2=0.234
r107 111 115 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.324 $Y=0.234 $X2=0.432 $Y2=0.234
r108 109 138 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.152 $Y=0.234 $X2=1.161 $Y2=0.225
r109 109 136 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.152 $Y=0.234 $X2=1.138 $Y2=0.234
r110 107 108 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.124 $Y=0.036 $X2=1.138 $Y2=0.036
r111 105 107 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.036 $X2=1.124 $Y2=0.036
r112 105 106 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.036
+ $X2=1.08 $Y2=0.036
r113 102 105 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.972 $Y=0.036 $X2=1.08 $Y2=0.036
r114 102 103 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.036
+ $X2=0.972 $Y2=0.036
r115 99 102 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.972 $Y2=0.036
r116 99 100 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036
+ $X2=0.864 $Y2=0.036
r117 96 99 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.864 $Y2=0.036
r118 96 97 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036
+ $X2=0.756 $Y2=0.036
r119 93 96 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.756 $Y2=0.036
r120 93 94 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r121 90 93 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.648 $Y2=0.036
r122 90 91 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r123 87 90 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.54 $Y2=0.036
r124 87 88 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r125 83 87 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r126 83 84 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r127 81 137 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.152 $Y=0.036 $X2=1.161 $Y2=0.045
r128 81 108 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.152
+ $Y=0.036 $X2=1.138 $Y2=0.036
r129 80 133 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234 $X2=1.08
+ $Y2=0.234
r130 77 80 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2025 $X2=1.08 $Y2=0.2025
r131 76 80 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.097 $Y=0.2025 $X2=1.08 $Y2=0.2025
r132 75 130 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.234
+ $X2=0.972 $Y2=0.234
r133 72 75 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.2025 $X2=0.972 $Y2=0.2025
r134 71 75 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.989 $Y=0.2025 $X2=0.972 $Y2=0.2025
r135 70 127 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234
+ $X2=0.864 $Y2=0.234
r136 67 70 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2025 $X2=0.864 $Y2=0.2025
r137 66 70 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2025 $X2=0.864 $Y2=0.2025
r138 65 124 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234
+ $X2=0.756 $Y2=0.234
r139 62 65 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r140 61 65 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r141 60 121 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234
+ $X2=0.648 $Y2=0.234
r142 57 60 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.648 $Y2=0.2025
r143 56 60 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.648 $Y2=0.2025
r144 55 118 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r145 52 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r146 51 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r147 50 115 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r148 47 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r149 46 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r150 45 111 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r151 42 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r152 41 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r153 40 106 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=1.08 $Y=0.0675 $X2=1.08 $Y2=0.036
r154 37 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.0675 $X2=1.08 $Y2=0.0675
r155 36 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.097 $Y=0.0675 $X2=1.08 $Y2=0.0675
r156 35 103 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.972 $Y=0.0675 $X2=0.972 $Y2=0.036
r157 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.0675 $X2=0.972 $Y2=0.0675
r158 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.989 $Y=0.0675 $X2=0.972 $Y2=0.0675
r159 30 100 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.864 $Y=0.0675 $X2=0.864 $Y2=0.036
r160 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0675 $X2=0.864 $Y2=0.0675
r161 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0675 $X2=0.864 $Y2=0.0675
r162 25 97 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.756 $Y=0.0675 $X2=0.756 $Y2=0.036
r163 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.756 $Y2=0.0675
r164 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.756 $Y2=0.0675
r165 20 94 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r166 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.648 $Y2=0.0675
r167 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0675 $X2=0.648 $Y2=0.0675
r168 15 91 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r169 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r170 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r171 10 88 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r172 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r173 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r174 5 84 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r175 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r176 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
.ends


* END of "./BUFx16f_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx16f_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_4_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_4_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_4_M2_d N_A_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_4_M3_d N_A_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_4_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_4_M6_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_4_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_4_M8_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_4_M9_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 N_Y_M10_d N_4_M10_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M11 N_Y_M11_d N_4_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M12 N_Y_M12_d N_4_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M13 N_Y_M13_d N_4_M13_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.027
M14 N_Y_M14_d N_4_M14_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.027
M15 N_Y_M15_d N_4_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.027
M16 N_Y_M16_d N_4_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.027
M17 N_Y_M17_d N_4_M17_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M18 N_Y_M18_d N_4_M18_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.027
M19 N_Y_M19_d N_4_M19_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.027
M20 N_4_M20_d N_A_M20_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M21 N_4_M21_d N_A_M21_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M22 N_4_M22_d N_A_M22_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M23 N_4_M23_d N_A_M23_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M24 N_Y_M24_d N_4_M24_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M25 N_Y_M25_d N_4_M25_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M26 N_Y_M26_d N_4_M26_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M27 N_Y_M27_d N_4_M27_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M28 N_Y_M28_d N_4_M28_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M29 N_Y_M29_d N_4_M29_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M30 N_Y_M30_d N_4_M30_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M31 N_Y_M31_d N_4_M31_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
M32 N_Y_M32_d N_4_M32_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M33 N_Y_M33_d N_4_M33_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
M34 N_Y_M34_d N_4_M34_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.162
M35 N_Y_M35_d N_4_M35_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.162
M36 N_Y_M36_d N_4_M36_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.162
M37 N_Y_M37_d N_4_M37_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
M38 N_Y_M38_d N_4_M38_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.162
M39 N_Y_M39_d N_4_M39_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.162
*
* 
* .include "BUFx16f_ASAP7_75t_SRAM.pex.sp.BUFX16F_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx16f_ASAP7_75t_SRAM.pex.sp.BUFX16F_ASAP7_75T_SRAM.pxi"
* File: BUFx16f_ASAP7_75t_SRAM.pex.sp.BUFX16F_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:18:54 2017
* 
x_PM_BUFX16F_ASAP7_75T_SRAM%A N_A_M0_g N_A_M20_g N_A_M1_g N_A_M21_g N_A_M2_g
+ N_A_M22_g N_A_M3_g N_A_c_4_p N_A_M23_g N_A_c_9_p A VSS
+ PM_BUFX16F_ASAP7_75T_SRAM%A
x_PM_BUFX16F_ASAP7_75T_SRAM%4 N_4_M4_g N_4_M24_g N_4_M5_g N_4_M25_g N_4_M6_g
+ N_4_M26_g N_4_M7_g N_4_M27_g N_4_M8_g N_4_M28_g N_4_M9_g N_4_M29_g N_4_M10_g
+ N_4_M30_g N_4_M11_g N_4_M31_g N_4_M12_g N_4_M32_g N_4_M13_g N_4_M33_g
+ N_4_M14_g N_4_M34_g N_4_M15_g N_4_M35_g N_4_M16_g N_4_M36_g N_4_M17_g
+ N_4_M37_g N_4_M18_g N_4_M38_g N_4_M19_g N_4_c_32_n N_4_M39_g N_4_M1_d N_4_M0_d
+ N_4_M3_d N_4_M2_d N_4_M21_d N_4_M20_d N_4_c_36_n N_4_M23_d N_4_M22_d
+ N_4_c_39_n N_4_c_40_n N_4_c_43_n N_4_c_45_n N_4_c_46_n N_4_c_49_n N_4_c_51_n
+ N_4_c_53_n N_4_c_55_n N_4_c_90_p N_4_c_110_p N_4_c_56_n VSS
+ PM_BUFX16F_ASAP7_75T_SRAM%4
x_PM_BUFX16F_ASAP7_75T_SRAM%Y N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M6_d N_Y_M9_d N_Y_M8_d
+ N_Y_M11_d N_Y_M10_d N_Y_M13_d N_Y_M12_d N_Y_M15_d N_Y_M14_d N_Y_M17_d
+ N_Y_M16_d N_Y_M19_d N_Y_M18_d N_Y_M25_d N_Y_M24_d N_Y_M27_d N_Y_M26_d
+ N_Y_M29_d N_Y_M28_d N_Y_M31_d N_Y_M30_d N_Y_M33_d N_Y_M32_d N_Y_M35_d
+ N_Y_M34_d N_Y_M37_d N_Y_M36_d N_Y_M39_d N_Y_M38_d N_Y_c_127_n N_Y_c_145_n Y
+ N_Y_c_163_n VSS PM_BUFX16F_ASAP7_75T_SRAM%Y
cc_1 N_A_M2_g N_4_M4_g 2.34385e-19 $X=0.189 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_2 N_A_M3_g N_4_M4_g 0.00287079f $X=0.243 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_3 N_A_M3_g N_4_M5_g 2.34385e-19 $X=0.243 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_4 N_A_c_4_p N_4_c_32_n 0.00159669f $X=0.243 $Y=0.135 $X2=1.107 $Y2=0.135
cc_5 N_A_c_4_p N_4_M1_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_6 N_A_c_4_p N_4_M3_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.233 $Y2=0.0675
cc_7 N_A_c_4_p N_4_M21_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_8 N_A_c_4_p N_4_c_36_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_9 N_A_c_9_p N_4_c_36_n 0.00115917f $X=0.064 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_10 N_A_c_4_p N_4_M23_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.233 $Y2=0.2025
cc_11 N_A_c_4_p N_4_c_39_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.216 $Y2=0.2025
cc_12 N_A_M1_g N_4_c_40_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.234 $Y2=0.036
cc_13 N_A_M2_g N_4_c_40_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.234 $Y2=0.036
cc_14 N_A_c_4_p N_4_c_40_n 0.00169924f $X=0.243 $Y=0.135 $X2=0.234 $Y2=0.036
cc_15 N_A_c_4_p N_4_c_43_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.108 $Y2=0.036
cc_16 N_A_c_9_p N_4_c_43_n 0.00115917f $X=0.064 $Y=0.135 $X2=0.108 $Y2=0.036
cc_17 N_A_c_4_p N_4_c_45_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.216 $Y2=0.036
cc_18 N_A_M1_g N_4_c_46_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.234 $Y2=0.234
cc_19 N_A_M2_g N_4_c_46_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.234 $Y2=0.234
cc_20 N_A_c_4_p N_4_c_46_n 0.00169924f $X=0.243 $Y=0.135 $X2=0.234 $Y2=0.234
cc_21 N_A_M3_g N_4_c_49_n 3.38818e-19 $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.126
cc_22 N_A_c_4_p N_4_c_49_n 4.8779e-19 $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.126
cc_23 N_A_M3_g N_4_c_51_n 2.9712e-19 $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.0965
cc_24 N_A_c_9_p N_4_c_51_n 6.83571e-19 $X=0.064 $Y=0.135 $X2=0.243 $Y2=0.0965
cc_25 N_A_M3_g N_4_c_53_n 6.35938e-19 $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.203
cc_26 N_A_c_4_p N_4_c_53_n 4.8779e-19 $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.203
cc_27 N_A_c_4_p N_4_c_55_n 4.66834e-19 $X=0.243 $Y=0.135 $X2=0.31 $Y2=0.135
cc_28 N_A_c_4_p N_4_c_56_n 0.00152364f $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.135
cc_29 N_4_c_32_n N_Y_M5_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_30 N_4_c_32_n N_Y_M7_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_31 N_4_c_32_n N_Y_M9_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_32 N_4_c_32_n N_Y_M11_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_33 N_4_c_32_n N_Y_M13_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0.189 $Y2=0.135
cc_34 N_4_c_32_n N_Y_M15_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_35 N_4_c_32_n N_Y_M17_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0.243 $Y2=0.2025
cc_36 N_4_c_32_n N_Y_M19_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_32_n N_Y_M25_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_32_n N_Y_M27_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_39 N_4_c_32_n N_Y_M29_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_32_n N_Y_M31_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_41 N_4_c_32_n N_Y_M33_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_42 N_4_c_32_n N_Y_M35_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_43 N_4_c_32_n N_Y_M37_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_44 N_4_c_32_n N_Y_M39_d 3.80218e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_45 N_4_M5_g N_Y_c_127_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_46 N_4_M6_g N_Y_c_127_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_4_M7_g N_Y_c_127_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_48 N_4_M8_g N_Y_c_127_n 4.28653e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_49 N_4_M9_g N_Y_c_127_n 4.28653e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_50 N_4_M10_g N_Y_c_127_n 4.28653e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_51 N_4_M11_g N_Y_c_127_n 4.28653e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_52 N_4_M12_g N_Y_c_127_n 4.28653e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_53 N_4_M13_g N_Y_c_127_n 4.28653e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_54 N_4_M14_g N_Y_c_127_n 4.28653e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_55 N_4_M15_g N_Y_c_127_n 4.28653e-19 $X=0.891 $Y=0.0675 $X2=0 $Y2=0
cc_56 N_4_M16_g N_Y_c_127_n 4.28653e-19 $X=0.945 $Y=0.0675 $X2=0 $Y2=0
cc_57 N_4_M17_g N_Y_c_127_n 4.28653e-19 $X=0.999 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_4_M18_g N_Y_c_127_n 4.28653e-19 $X=1.053 $Y=0.0675 $X2=0 $Y2=0
cc_59 N_4_M19_g N_Y_c_127_n 4.28653e-19 $X=1.107 $Y=0.0675 $X2=0 $Y2=0
cc_60 N_4_c_32_n N_Y_c_127_n 0.00298598f $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_61 N_4_c_40_n N_Y_c_127_n 4.53942e-19 $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_62 N_4_c_90_p N_Y_c_127_n 0.011021f $X=0.3305 $Y=0.135 $X2=0 $Y2=0
cc_63 N_4_M5_g N_Y_c_145_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_4_M6_g N_Y_c_145_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_65 N_4_M7_g N_Y_c_145_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_66 N_4_M8_g N_Y_c_145_n 4.28653e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_67 N_4_M9_g N_Y_c_145_n 4.28653e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_68 N_4_M10_g N_Y_c_145_n 4.28653e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_69 N_4_M11_g N_Y_c_145_n 4.28653e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_70 N_4_M12_g N_Y_c_145_n 4.28653e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_71 N_4_M13_g N_Y_c_145_n 4.28653e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_72 N_4_M14_g N_Y_c_145_n 4.28653e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_73 N_4_M15_g N_Y_c_145_n 4.28653e-19 $X=0.891 $Y=0.0675 $X2=0 $Y2=0
cc_74 N_4_M16_g N_Y_c_145_n 4.28653e-19 $X=0.945 $Y=0.0675 $X2=0 $Y2=0
cc_75 N_4_M17_g N_Y_c_145_n 4.28653e-19 $X=0.999 $Y=0.0675 $X2=0 $Y2=0
cc_76 N_4_M18_g N_Y_c_145_n 4.28653e-19 $X=1.053 $Y=0.0675 $X2=0 $Y2=0
cc_77 N_4_M19_g N_Y_c_145_n 4.28653e-19 $X=1.107 $Y=0.0675 $X2=0 $Y2=0
cc_78 N_4_c_32_n N_Y_c_145_n 0.00298598f $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_79 N_4_c_46_n N_Y_c_145_n 4.53942e-19 $X=0.234 $Y=0.234 $X2=0 $Y2=0
cc_80 N_4_c_90_p N_Y_c_145_n 0.011021f $X=0.3305 $Y=0.135 $X2=0 $Y2=0
cc_81 N_4_c_32_n N_Y_c_163_n 4.69552e-19 $X=1.107 $Y=0.135 $X2=0 $Y2=0
cc_82 N_4_c_110_p N_Y_c_163_n 0.00114058f $X=1.107 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx16f_ASAP7_75t_SRAM.pex.sp.BUFX16F_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx24_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:19:17 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx24_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx24_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx24_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:19:17 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX24_ASAP7_75T_SRAM%A 2 7 10 15 18 23 26 29 31 39 VSS
c26 39 VSS 0.027631f $X=0.061 $Y=0.1335
c27 29 VSS 0.0184912f $X=0.243 $Y=0.135
c28 26 VSS 0.0609562f $X=0.243 $Y=0.0675
c29 18 VSS 0.0642127f $X=0.189 $Y=0.0675
c30 10 VSS 0.0644226f $X=0.135 $Y=0.0675
c31 2 VSS 0.0655089f $X=0.081 $Y=0.0675
r32 39 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r33 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r34 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r35 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r36 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r37 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r38 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r39 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r40 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r41 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r42 5 43 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r43 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r44 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX24_ASAP7_75T_SRAM%4 2 7 10 15 18 23 26 31 34 39 42 47 50 55 58 63 66
+ 71 74 79 82 87 90 95 98 103 106 111 114 119 122 127 130 135 138 143 146 151
+ 154 159 162 167 170 175 178 183 186 189 191 193 194 198 199 203 204 207 208
+ 209 212 213 216 220 221 230 232 237 238 258 261 VSS
c104 261 VSS 1.38647e-19 $X=0.243 $Y=0.135
c105 258 VSS 3.05218e-19 $X=1.485 $Y=0.135
c106 237 VSS 0.00280817f $X=0.31 $Y=0.135
c107 232 VSS 0.00386854f $X=0.243 $Y=0.225
c108 230 VSS 0.00386854f $X=0.243 $Y=0.126
c109 221 VSS 0.0187138f $X=0.234 $Y=0.234
c110 220 VSS 0.0104726f $X=0.216 $Y=0.036
c111 216 VSS 0.00904032f $X=0.108 $Y=0.036
c112 213 VSS 0.0187138f $X=0.234 $Y=0.036
c113 212 VSS 0.0104726f $X=0.216 $Y=0.2025
c114 208 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c115 207 VSS 0.00904032f $X=0.108 $Y=0.2025
c116 203 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c117 198 VSS 5.38922e-19 $X=0.233 $Y=0.0675
c118 193 VSS 5.72268e-19 $X=0.125 $Y=0.0675
c119 189 VSS 0.0823945f $X=1.539 $Y=0.135
c120 186 VSS 0.0645347f $X=1.539 $Y=0.0675
c121 178 VSS 0.0644226f $X=1.485 $Y=0.0675
c122 170 VSS 0.0642127f $X=1.431 $Y=0.0675
c123 162 VSS 0.0642127f $X=1.377 $Y=0.0675
c124 154 VSS 0.0642127f $X=1.323 $Y=0.0675
c125 146 VSS 0.0642127f $X=1.269 $Y=0.0675
c126 138 VSS 0.0642127f $X=1.215 $Y=0.0675
c127 130 VSS 0.0642127f $X=1.161 $Y=0.0675
c128 122 VSS 0.0642127f $X=1.107 $Y=0.0675
c129 114 VSS 0.0642127f $X=1.053 $Y=0.0675
c130 106 VSS 0.0642127f $X=0.999 $Y=0.0675
c131 98 VSS 0.0642127f $X=0.945 $Y=0.0675
c132 90 VSS 0.0642127f $X=0.891 $Y=0.0675
c133 82 VSS 0.0642127f $X=0.837 $Y=0.0675
c134 74 VSS 0.0642127f $X=0.783 $Y=0.0675
c135 66 VSS 0.0642127f $X=0.729 $Y=0.0675
c136 58 VSS 0.0642127f $X=0.675 $Y=0.0675
c137 50 VSS 0.0642127f $X=0.621 $Y=0.0675
c138 42 VSS 0.0642127f $X=0.567 $Y=0.0675
c139 34 VSS 0.0642127f $X=0.513 $Y=0.0675
c140 26 VSS 0.0642127f $X=0.459 $Y=0.0675
c141 18 VSS 0.0642127f $X=0.405 $Y=0.0675
c142 10 VSS 0.0642127f $X=0.351 $Y=0.0675
c143 2 VSS 0.0616955f $X=0.297 $Y=0.0675
r144 255 258 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=1.323
+ $Y=0.135 $X2=1.485 $Y2=0.135
r145 252 255 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=1.161
+ $Y=0.135 $X2=1.323 $Y2=0.135
r146 249 252 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.999
+ $Y=0.135 $X2=1.161 $Y2=0.135
r147 246 249 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.135 $X2=0.999 $Y2=0.135
r148 243 246 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.135 $X2=0.837 $Y2=0.135
r149 240 243 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.675 $Y2=0.135
r150 237 238 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.31
+ $Y=0.135 $X2=0.3305 $Y2=0.135
r151 235 240 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.513 $Y2=0.135
r152 235 238 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.351 $Y=0.135 $X2=0.3305 $Y2=0.135
r153 233 261 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.243 $Y2=0.135
r154 233 237 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.135 $X2=0.31 $Y2=0.135
r155 231 261 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.144 $X2=0.243 $Y2=0.135
r156 231 232 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.144 $X2=0.243 $Y2=0.225
r157 230 261 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.135
r158 229 230 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.126
r159 223 227 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.108 $Y=0.234 $X2=0.216 $Y2=0.234
r160 221 232 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r161 221 227 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r162 219 220 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r163 215 219 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.108 $Y=0.036 $X2=0.216 $Y2=0.036
r164 215 216 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r165 213 229 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r166 213 219 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r167 212 227 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r168 209 212 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r169 208 212 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r170 207 223 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r171 204 207 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r172 203 207 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r173 202 220 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.216 $Y=0.0675 $X2=0.216 $Y2=0.036
r174 199 202 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r175 198 202 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r176 197 216 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.108 $Y=0.0675 $X2=0.108 $Y2=0.036
r177 194 197 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r178 193 197 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r179 189 191 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.539 $Y=0.135 $X2=1.539 $Y2=0.2025
r180 186 189 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.539 $Y=0.0675 $X2=1.539 $Y2=0.135
r181 181 189 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.485
+ $Y=0.135 $X2=1.539 $Y2=0.135
r182 181 258 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=1.485 $Y=0.135
+ $X2=1.485 $Y2=0.135
r183 181 183 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.485 $Y=0.135 $X2=1.485 $Y2=0.2025
r184 178 181 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.485 $Y=0.0675 $X2=1.485 $Y2=0.135
r185 173 181 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.431
+ $Y=0.135 $X2=1.485 $Y2=0.135
r186 173 175 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.431 $Y=0.135 $X2=1.431 $Y2=0.2025
r187 170 173 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.431 $Y=0.0675 $X2=1.431 $Y2=0.135
r188 165 173 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.377
+ $Y=0.135 $X2=1.431 $Y2=0.135
r189 165 167 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.377 $Y=0.135 $X2=1.377 $Y2=0.2025
r190 162 165 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.377 $Y=0.0675 $X2=1.377 $Y2=0.135
r191 157 165 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.323
+ $Y=0.135 $X2=1.377 $Y2=0.135
r192 157 255 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=1.323 $Y=0.135
+ $X2=1.323 $Y2=0.135
r193 157 159 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.135 $X2=1.323 $Y2=0.2025
r194 154 157 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.323 $Y=0.0675 $X2=1.323 $Y2=0.135
r195 149 157 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.269
+ $Y=0.135 $X2=1.323 $Y2=0.135
r196 149 151 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.135 $X2=1.269 $Y2=0.2025
r197 146 149 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.269 $Y=0.0675 $X2=1.269 $Y2=0.135
r198 141 149 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.215
+ $Y=0.135 $X2=1.269 $Y2=0.135
r199 141 143 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.135 $X2=1.215 $Y2=0.2025
r200 138 141 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.215 $Y=0.0675 $X2=1.215 $Y2=0.135
r201 133 141 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.161
+ $Y=0.135 $X2=1.215 $Y2=0.135
r202 133 252 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=1.161 $Y=0.135
+ $X2=1.161 $Y2=0.135
r203 133 135 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.161 $Y=0.135 $X2=1.161 $Y2=0.2025
r204 130 133 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.161 $Y=0.0675 $X2=1.161 $Y2=0.135
r205 125 133 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.107
+ $Y=0.135 $X2=1.161 $Y2=0.135
r206 125 127 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.135 $X2=1.107 $Y2=0.2025
r207 122 125 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.107 $Y=0.0675 $X2=1.107 $Y2=0.135
r208 117 125 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=1.053
+ $Y=0.135 $X2=1.107 $Y2=0.135
r209 117 119 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.135 $X2=1.053 $Y2=0.2025
r210 114 117 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=1.053 $Y=0.0675 $X2=1.053 $Y2=0.135
r211 109 117 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.999
+ $Y=0.135 $X2=1.053 $Y2=0.135
r212 109 249 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.999 $Y=0.135
+ $X2=0.999 $Y2=0.135
r213 109 111 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.135 $X2=0.999 $Y2=0.2025
r214 106 109 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.135
r215 101 109 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.945
+ $Y=0.135 $X2=0.999 $Y2=0.135
r216 101 103 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.135 $X2=0.945 $Y2=0.2025
r217 98 101 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.945 $Y=0.0675 $X2=0.945 $Y2=0.135
r218 93 101 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.891
+ $Y=0.135 $X2=0.945 $Y2=0.135
r219 93 95 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.135 $X2=0.891 $Y2=0.2025
r220 90 93 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.891 $Y=0.0675 $X2=0.891 $Y2=0.135
r221 85 93 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.837
+ $Y=0.135 $X2=0.891 $Y2=0.135
r222 85 246 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.837 $Y=0.135
+ $X2=0.837 $Y2=0.135
r223 85 87 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.135 $X2=0.837 $Y2=0.2025
r224 82 85 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0675 $X2=0.837 $Y2=0.135
r225 77 85 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.783
+ $Y=0.135 $X2=0.837 $Y2=0.135
r226 77 79 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.135 $X2=0.783 $Y2=0.2025
r227 74 77 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.135
r228 69 77 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.135 $X2=0.783 $Y2=0.135
r229 69 71 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.135 $X2=0.729 $Y2=0.2025
r230 66 69 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.135
r231 61 69 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.729 $Y2=0.135
r232 61 243 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.675 $Y=0.135
+ $X2=0.675 $Y2=0.135
r233 61 63 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2025
r234 58 61 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0675 $X2=0.675 $Y2=0.135
r235 53 61 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621
+ $Y=0.135 $X2=0.675 $Y2=0.135
r236 53 55 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2025
r237 50 53 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r238 45 53 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.567
+ $Y=0.135 $X2=0.621 $Y2=0.135
r239 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.135 $X2=0.567 $Y2=0.2025
r240 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.0675 $X2=0.567 $Y2=0.135
r241 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r242 37 240 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.513 $Y=0.135
+ $X2=0.513 $Y2=0.135
r243 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r244 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r245 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r246 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r247 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r248 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r249 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r250 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r251 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r252 13 235 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.351 $Y=0.135
+ $X2=0.351 $Y2=0.135
r253 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r254 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r255 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r256 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r257 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_BUFX24_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 21 22 26 27 31 32 36 37 41
+ 42 46 47 51 52 56 57 61 62 66 67 71 72 76 77 81 82 86 87 91 92 96 97 101 102
+ 106 107 111 112 116 117 159 199 204 206 VSS
c78 206 VSS 7.46953e-19 $X=1.593 $Y=0.144
c79 205 VSS 0.00538047f $X=1.593 $Y=0.126
c80 204 VSS 0.00538047f $X=1.595 $Y=0.1495
c81 200 VSS 0.00294383f $X=1.5685 $Y=0.234
c82 199 VSS 0.131925f $X=1.553 $Y=0.234
c83 161 VSS 0.00593798f $X=1.584 $Y=0.234
c84 160 VSS 0.00294383f $X=1.5685 $Y=0.036
c85 159 VSS 0.131925f $X=1.553 $Y=0.036
c86 158 VSS 0.00929752f $X=1.512 $Y=0.036
c87 155 VSS 0.00928953f $X=1.404 $Y=0.036
c88 152 VSS 0.00928955f $X=1.296 $Y=0.036
c89 149 VSS 0.00928955f $X=1.188 $Y=0.036
c90 146 VSS 0.00928955f $X=1.08 $Y=0.036
c91 143 VSS 0.00928955f $X=0.972 $Y=0.036
c92 140 VSS 0.00928955f $X=0.864 $Y=0.036
c93 137 VSS 0.00928955f $X=0.756 $Y=0.036
c94 134 VSS 0.00928955f $X=0.648 $Y=0.036
c95 131 VSS 0.00928955f $X=0.54 $Y=0.036
c96 128 VSS 0.00928953f $X=0.432 $Y=0.036
c97 124 VSS 0.00917567f $X=0.324 $Y=0.036
c98 121 VSS 0.00593798f $X=1.584 $Y=0.036
c99 120 VSS 0.00929752f $X=1.512 $Y=0.2025
c100 116 VSS 5.38922e-19 $X=1.529 $Y=0.2025
c101 115 VSS 0.00928953f $X=1.404 $Y=0.2025
c102 111 VSS 5.38922e-19 $X=1.421 $Y=0.2025
c103 110 VSS 0.00928955f $X=1.296 $Y=0.2025
c104 106 VSS 5.38922e-19 $X=1.313 $Y=0.2025
c105 105 VSS 0.00928955f $X=1.188 $Y=0.2025
c106 101 VSS 5.38922e-19 $X=1.205 $Y=0.2025
c107 100 VSS 0.00928955f $X=1.08 $Y=0.2025
c108 96 VSS 5.38922e-19 $X=1.097 $Y=0.2025
c109 95 VSS 0.00928955f $X=0.972 $Y=0.2025
c110 91 VSS 5.38922e-19 $X=0.989 $Y=0.2025
c111 90 VSS 0.00928955f $X=0.864 $Y=0.2025
c112 86 VSS 5.38922e-19 $X=0.881 $Y=0.2025
c113 85 VSS 0.00928955f $X=0.756 $Y=0.2025
c114 81 VSS 5.38922e-19 $X=0.773 $Y=0.2025
c115 80 VSS 0.00928955f $X=0.648 $Y=0.2025
c116 76 VSS 5.38922e-19 $X=0.665 $Y=0.2025
c117 75 VSS 0.00928955f $X=0.54 $Y=0.2025
c118 71 VSS 5.38922e-19 $X=0.557 $Y=0.2025
c119 70 VSS 0.00928953f $X=0.432 $Y=0.2025
c120 66 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c121 65 VSS 0.00917567f $X=0.324 $Y=0.2025
c122 61 VSS 5.72268e-19 $X=0.341 $Y=0.2025
c123 56 VSS 5.38922e-19 $X=1.529 $Y=0.0675
c124 51 VSS 5.38922e-19 $X=1.421 $Y=0.0675
c125 46 VSS 5.38922e-19 $X=1.313 $Y=0.0675
c126 41 VSS 5.38922e-19 $X=1.205 $Y=0.0675
c127 36 VSS 5.38922e-19 $X=1.097 $Y=0.0675
c128 31 VSS 5.38922e-19 $X=0.989 $Y=0.0675
c129 26 VSS 5.38922e-19 $X=0.881 $Y=0.0675
c130 21 VSS 5.38922e-19 $X=0.773 $Y=0.0675
c131 16 VSS 5.38922e-19 $X=0.665 $Y=0.0675
c132 11 VSS 5.38922e-19 $X=0.557 $Y=0.0675
c133 6 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c134 1 VSS 5.72268e-19 $X=0.341 $Y=0.0675
r135 205 206 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.593
+ $Y=0.126 $X2=1.593 $Y2=0.144
r136 204 206 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08
+ $X=1.593 $Y=0.1495 $X2=1.593 $Y2=0.144
r137 202 204 5.12654 $w=1.8e-08 $l=7.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.593 $Y=0.225 $X2=1.593 $Y2=0.1495
r138 201 205 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.593
+ $Y=0.045 $X2=1.593 $Y2=0.126
r139 199 200 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.553 $Y=0.234 $X2=1.5685 $Y2=0.234
r140 197 199 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.512
+ $Y=0.234 $X2=1.553 $Y2=0.234
r141 194 197 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=1.404 $Y=0.234 $X2=1.512 $Y2=0.234
r142 191 194 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=1.296 $Y=0.234 $X2=1.404 $Y2=0.234
r143 188 191 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=1.188 $Y=0.234 $X2=1.296 $Y2=0.234
r144 185 188 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.234 $X2=1.188 $Y2=0.234
r145 182 185 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.972 $Y=0.234 $X2=1.08 $Y2=0.234
r146 179 182 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.864 $Y=0.234 $X2=0.972 $Y2=0.234
r147 176 179 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.756 $Y=0.234 $X2=0.864 $Y2=0.234
r148 173 176 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.648 $Y=0.234 $X2=0.756 $Y2=0.234
r149 170 173 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.648 $Y2=0.234
r150 167 170 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.432 $Y=0.234 $X2=0.54 $Y2=0.234
r151 163 167 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.324 $Y=0.234 $X2=0.432 $Y2=0.234
r152 161 202 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.584 $Y=0.234 $X2=1.593 $Y2=0.225
r153 161 200 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.584 $Y=0.234 $X2=1.5685 $Y2=0.234
r154 159 160 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.553 $Y=0.036 $X2=1.5685 $Y2=0.036
r155 157 159 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.512
+ $Y=0.036 $X2=1.553 $Y2=0.036
r156 157 158 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.512 $Y=0.036
+ $X2=1.512 $Y2=0.036
r157 154 157 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=1.404 $Y=0.036 $X2=1.512 $Y2=0.036
r158 154 155 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.404 $Y=0.036
+ $X2=1.404 $Y2=0.036
r159 151 154 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=1.296 $Y=0.036 $X2=1.404 $Y2=0.036
r160 151 152 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.036
+ $X2=1.296 $Y2=0.036
r161 148 151 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=1.188 $Y=0.036 $X2=1.296 $Y2=0.036
r162 148 149 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.188 $Y=0.036
+ $X2=1.188 $Y2=0.036
r163 145 148 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=1.08
+ $Y=0.036 $X2=1.188 $Y2=0.036
r164 145 146 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.036
+ $X2=1.08 $Y2=0.036
r165 142 145 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.972 $Y=0.036 $X2=1.08 $Y2=0.036
r166 142 143 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.036
+ $X2=0.972 $Y2=0.036
r167 139 142 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.864 $Y=0.036 $X2=0.972 $Y2=0.036
r168 139 140 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036
+ $X2=0.864 $Y2=0.036
r169 136 139 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.756 $Y=0.036 $X2=0.864 $Y2=0.036
r170 136 137 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036
+ $X2=0.756 $Y2=0.036
r171 133 136 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.648 $Y=0.036 $X2=0.756 $Y2=0.036
r172 133 134 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r173 130 133 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.648 $Y2=0.036
r174 130 131 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036
+ $X2=0.54 $Y2=0.036
r175 127 130 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.432 $Y=0.036 $X2=0.54 $Y2=0.036
r176 127 128 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r177 123 127 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.324 $Y=0.036 $X2=0.432 $Y2=0.036
r178 123 124 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r179 121 201 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.584 $Y=0.036 $X2=1.593 $Y2=0.045
r180 121 160 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.584 $Y=0.036 $X2=1.5685 $Y2=0.036
r181 120 197 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.512 $Y=0.234
+ $X2=1.512 $Y2=0.234
r182 117 120 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.495 $Y=0.2025 $X2=1.512 $Y2=0.2025
r183 116 120 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.529 $Y=0.2025 $X2=1.512 $Y2=0.2025
r184 115 194 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.404 $Y=0.234
+ $X2=1.404 $Y2=0.234
r185 112 115 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.387 $Y=0.2025 $X2=1.404 $Y2=0.2025
r186 111 115 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.421 $Y=0.2025 $X2=1.404 $Y2=0.2025
r187 110 191 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.296 $Y=0.234
+ $X2=1.296 $Y2=0.234
r188 107 110 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.279 $Y=0.2025 $X2=1.296 $Y2=0.2025
r189 106 110 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.313 $Y=0.2025 $X2=1.296 $Y2=0.2025
r190 105 188 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.188 $Y=0.234
+ $X2=1.188 $Y2=0.234
r191 102 105 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.171 $Y=0.2025 $X2=1.188 $Y2=0.2025
r192 101 105 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.2025 $X2=1.188 $Y2=0.2025
r193 100 185 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.08 $Y=0.234
+ $X2=1.08 $Y2=0.234
r194 97 100 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.2025 $X2=1.08 $Y2=0.2025
r195 96 100 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.097 $Y=0.2025 $X2=1.08 $Y2=0.2025
r196 95 182 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.234
+ $X2=0.972 $Y2=0.234
r197 92 95 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.2025 $X2=0.972 $Y2=0.2025
r198 91 95 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.989 $Y=0.2025 $X2=0.972 $Y2=0.2025
r199 90 179 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234
+ $X2=0.864 $Y2=0.234
r200 87 90 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2025 $X2=0.864 $Y2=0.2025
r201 86 90 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2025 $X2=0.864 $Y2=0.2025
r202 85 176 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234
+ $X2=0.756 $Y2=0.234
r203 82 85 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r204 81 85 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r205 80 173 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234
+ $X2=0.648 $Y2=0.234
r206 77 80 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.648 $Y2=0.2025
r207 76 80 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.648 $Y2=0.2025
r208 75 170 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r209 72 75 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r210 71 75 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r211 70 167 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r212 67 70 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r213 66 70 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r214 65 163 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r215 62 65 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r216 61 65 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r217 60 158 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=1.512 $Y=0.0675 $X2=1.512 $Y2=0.036
r218 57 60 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.495 $Y=0.0675 $X2=1.512 $Y2=0.0675
r219 56 60 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.529 $Y=0.0675 $X2=1.512 $Y2=0.0675
r220 55 155 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=1.404 $Y=0.0675 $X2=1.404 $Y2=0.036
r221 52 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.387 $Y=0.0675 $X2=1.404 $Y2=0.0675
r222 51 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.421 $Y=0.0675 $X2=1.404 $Y2=0.0675
r223 50 152 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=1.296 $Y=0.0675 $X2=1.296 $Y2=0.036
r224 47 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.279 $Y=0.0675 $X2=1.296 $Y2=0.0675
r225 46 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.313 $Y=0.0675 $X2=1.296 $Y2=0.0675
r226 45 149 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=1.188 $Y=0.0675 $X2=1.188 $Y2=0.036
r227 42 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.171 $Y=0.0675 $X2=1.188 $Y2=0.0675
r228 41 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.205 $Y=0.0675 $X2=1.188 $Y2=0.0675
r229 40 146 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=1.08 $Y=0.0675 $X2=1.08 $Y2=0.036
r230 37 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.063 $Y=0.0675 $X2=1.08 $Y2=0.0675
r231 36 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.097 $Y=0.0675 $X2=1.08 $Y2=0.0675
r232 35 143 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.972 $Y=0.0675 $X2=0.972 $Y2=0.036
r233 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.0675 $X2=0.972 $Y2=0.0675
r234 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.989 $Y=0.0675 $X2=0.972 $Y2=0.0675
r235 30 140 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.864 $Y=0.0675 $X2=0.864 $Y2=0.036
r236 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0675 $X2=0.864 $Y2=0.0675
r237 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0675 $X2=0.864 $Y2=0.0675
r238 25 137 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.756 $Y=0.0675 $X2=0.756 $Y2=0.036
r239 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.756 $Y2=0.0675
r240 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.756 $Y2=0.0675
r241 20 134 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r242 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.648 $Y2=0.0675
r243 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0675 $X2=0.648 $Y2=0.0675
r244 15 131 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.54 $Y=0.0675 $X2=0.54 $Y2=0.036
r245 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r246 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r247 10 128 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r248 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r249 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r250 5 124 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r251 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r252 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
.ends


* END of "./BUFx24_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx24_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_4_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_4_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_4_M2_d N_A_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_4_M3_d N_A_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_4_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_4_M6_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_4_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_4_M8_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_4_M9_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 N_Y_M10_d N_4_M10_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M11 N_Y_M11_d N_4_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M12 N_Y_M12_d N_4_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M13 N_Y_M13_d N_4_M13_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.027
M14 N_Y_M14_d N_4_M14_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.027
M15 N_Y_M15_d N_4_M15_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.027
M16 N_Y_M16_d N_4_M16_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.027
M17 N_Y_M17_d N_4_M17_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M18 N_Y_M18_d N_4_M18_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.027
M19 N_Y_M19_d N_4_M19_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.027
M20 N_Y_M20_d N_4_M20_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.151
+ $Y=0.027
M21 N_Y_M21_d N_4_M21_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.027
M22 N_Y_M22_d N_4_M22_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.027
M23 N_Y_M23_d N_4_M23_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.027
M24 N_Y_M24_d N_4_M24_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.367
+ $Y=0.027
M25 N_Y_M25_d N_4_M25_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.421
+ $Y=0.027
M26 N_Y_M26_d N_4_M26_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.475
+ $Y=0.027
M27 N_Y_M27_d N_4_M27_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.529
+ $Y=0.027
M28 N_4_M28_d N_A_M28_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M29 N_4_M29_d N_A_M29_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M30 N_4_M30_d N_A_M30_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M31 N_4_M31_d N_A_M31_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M32 N_Y_M32_d N_4_M32_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M33 N_Y_M33_d N_4_M33_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M34 N_Y_M34_d N_4_M34_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M35 N_Y_M35_d N_4_M35_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M36 N_Y_M36_d N_4_M36_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M37 N_Y_M37_d N_4_M37_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M38 N_Y_M38_d N_4_M38_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M39 N_Y_M39_d N_4_M39_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
M40 N_Y_M40_d N_4_M40_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M41 N_Y_M41_d N_4_M41_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
M42 N_Y_M42_d N_4_M42_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.162
M43 N_Y_M43_d N_4_M43_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.162
M44 N_Y_M44_d N_4_M44_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.162
M45 N_Y_M45_d N_4_M45_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
M46 N_Y_M46_d N_4_M46_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.043
+ $Y=0.162
M47 N_Y_M47_d N_4_M47_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.097
+ $Y=0.162
M48 N_Y_M48_d N_4_M48_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.151
+ $Y=0.162
M49 N_Y_M49_d N_4_M49_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.205
+ $Y=0.162
M50 N_Y_M50_d N_4_M50_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.259
+ $Y=0.162
M51 N_Y_M51_d N_4_M51_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.313
+ $Y=0.162
M52 N_Y_M52_d N_4_M52_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.367
+ $Y=0.162
M53 N_Y_M53_d N_4_M53_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.421
+ $Y=0.162
M54 N_Y_M54_d N_4_M54_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.475
+ $Y=0.162
M55 N_Y_M55_d N_4_M55_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=1.529
+ $Y=0.162
*
* 
* .include "BUFx24_ASAP7_75t_SRAM.pex.sp.BUFX24_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx24_ASAP7_75t_SRAM.pex.sp.BUFX24_ASAP7_75T_SRAM.pxi"
* File: BUFx24_ASAP7_75t_SRAM.pex.sp.BUFX24_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:19:17 2017
* 
x_PM_BUFX24_ASAP7_75T_SRAM%A N_A_M0_g N_A_M28_g N_A_M1_g N_A_M29_g N_A_M2_g
+ N_A_M30_g N_A_M3_g N_A_c_4_p N_A_M31_g A VSS PM_BUFX24_ASAP7_75T_SRAM%A
x_PM_BUFX24_ASAP7_75T_SRAM%4 N_4_M4_g N_4_M32_g N_4_M5_g N_4_M33_g N_4_M6_g
+ N_4_M34_g N_4_M7_g N_4_M35_g N_4_M8_g N_4_M36_g N_4_M9_g N_4_M37_g N_4_M10_g
+ N_4_M38_g N_4_M11_g N_4_M39_g N_4_M12_g N_4_M40_g N_4_M13_g N_4_M41_g
+ N_4_M14_g N_4_M42_g N_4_M15_g N_4_M43_g N_4_M16_g N_4_M44_g N_4_M17_g
+ N_4_M45_g N_4_M18_g N_4_M46_g N_4_M19_g N_4_M47_g N_4_M20_g N_4_M48_g
+ N_4_M21_g N_4_M49_g N_4_M22_g N_4_M50_g N_4_M23_g N_4_M51_g N_4_M24_g
+ N_4_M52_g N_4_M25_g N_4_M53_g N_4_M26_g N_4_M54_g N_4_M27_g N_4_c_30_n
+ N_4_M55_g N_4_M1_d N_4_M0_d N_4_M3_d N_4_M2_d N_4_M29_d N_4_M28_d N_4_c_34_n
+ N_4_M31_d N_4_M30_d N_4_c_36_n N_4_c_37_n N_4_c_41_n N_4_c_42_n N_4_c_43_n
+ N_4_c_47_n N_4_c_49_n N_4_c_51_n N_4_c_102_p N_4_c_130_p N_4_c_52_n VSS
+ PM_BUFX24_ASAP7_75T_SRAM%4
x_PM_BUFX24_ASAP7_75T_SRAM%Y N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M6_d N_Y_M9_d N_Y_M8_d
+ N_Y_M11_d N_Y_M10_d N_Y_M13_d N_Y_M12_d N_Y_M15_d N_Y_M14_d N_Y_M17_d
+ N_Y_M16_d N_Y_M19_d N_Y_M18_d N_Y_M21_d N_Y_M20_d N_Y_M23_d N_Y_M22_d
+ N_Y_M25_d N_Y_M24_d N_Y_M27_d N_Y_M26_d N_Y_M33_d N_Y_M32_d N_Y_M35_d
+ N_Y_M34_d N_Y_M37_d N_Y_M36_d N_Y_M39_d N_Y_M38_d N_Y_M41_d N_Y_M40_d
+ N_Y_M43_d N_Y_M42_d N_Y_M45_d N_Y_M44_d N_Y_M47_d N_Y_M46_d N_Y_M49_d
+ N_Y_M48_d N_Y_M51_d N_Y_M50_d N_Y_M53_d N_Y_M52_d N_Y_M55_d N_Y_M54_d
+ N_Y_c_155_n N_Y_c_181_n Y N_Y_c_207_n VSS PM_BUFX24_ASAP7_75T_SRAM%Y
cc_1 N_A_M2_g N_4_M4_g 2.34385e-19 $X=0.189 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_2 N_A_M3_g N_4_M4_g 0.00287079f $X=0.243 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_3 N_A_M3_g N_4_M5_g 2.34385e-19 $X=0.243 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_4 N_A_c_4_p N_4_c_30_n 0.00160439f $X=0.243 $Y=0.135 $X2=1.539 $Y2=0.135
cc_5 N_A_c_4_p N_4_M1_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_6 N_A_c_4_p N_4_M3_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.233 $Y2=0.0675
cc_7 N_A_c_4_p N_4_M29_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_8 N_A_c_4_p N_4_c_34_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_9 N_A_c_4_p N_4_M31_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.233 $Y2=0.2025
cc_10 N_A_c_4_p N_4_c_36_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.216 $Y2=0.2025
cc_11 N_A_M1_g N_4_c_37_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.234 $Y2=0.036
cc_12 N_A_M2_g N_4_c_37_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.234 $Y2=0.036
cc_13 N_A_c_4_p N_4_c_37_n 0.00169924f $X=0.243 $Y=0.135 $X2=0.234 $Y2=0.036
cc_14 A N_4_c_37_n 5.28865e-19 $X=0.061 $Y=0.1335 $X2=0.234 $Y2=0.036
cc_15 N_A_c_4_p N_4_c_41_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.108 $Y2=0.036
cc_16 N_A_c_4_p N_4_c_42_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.216 $Y2=0.036
cc_17 N_A_M1_g N_4_c_43_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.234 $Y2=0.234
cc_18 N_A_M2_g N_4_c_43_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.234 $Y2=0.234
cc_19 N_A_c_4_p N_4_c_43_n 0.00169924f $X=0.243 $Y=0.135 $X2=0.234 $Y2=0.234
cc_20 A N_4_c_43_n 5.28865e-19 $X=0.061 $Y=0.1335 $X2=0.234 $Y2=0.234
cc_21 N_A_M3_g N_4_c_47_n 5.85531e-19 $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.126
cc_22 N_A_c_4_p N_4_c_47_n 4.78945e-19 $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.126
cc_23 N_A_M3_g N_4_c_49_n 5.85531e-19 $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.225
cc_24 N_A_c_4_p N_4_c_49_n 4.78945e-19 $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.225
cc_25 N_A_c_4_p N_4_c_51_n 4.66834e-19 $X=0.243 $Y=0.135 $X2=0.31 $Y2=0.135
cc_26 N_A_c_4_p N_4_c_52_n 0.00153171f $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.135
cc_27 N_4_c_30_n N_Y_M5_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_28 N_4_c_30_n N_Y_M7_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_29 N_4_c_30_n N_Y_M9_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_30 N_4_c_30_n N_Y_M11_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_31 N_4_c_30_n N_Y_M13_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0.189 $Y2=0.135
cc_32 N_4_c_30_n N_Y_M15_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_33 N_4_c_30_n N_Y_M17_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0.243 $Y2=0.2025
cc_34 N_4_c_30_n N_Y_M19_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_35 N_4_c_30_n N_Y_M21_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_36 N_4_c_30_n N_Y_M23_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_30_n N_Y_M25_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_30_n N_Y_M27_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_39 N_4_c_30_n N_Y_M33_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_30_n N_Y_M35_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_41 N_4_c_30_n N_Y_M37_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_42 N_4_c_30_n N_Y_M39_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_43 N_4_c_30_n N_Y_M41_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_44 N_4_c_30_n N_Y_M43_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_45 N_4_c_30_n N_Y_M45_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_30_n N_Y_M47_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_47 N_4_c_30_n N_Y_M49_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_48 N_4_c_30_n N_Y_M51_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_49 N_4_c_30_n N_Y_M53_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_50 N_4_c_30_n N_Y_M55_d 3.80218e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_51 N_4_M5_g N_Y_c_155_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_52 N_4_M6_g N_Y_c_155_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_53 N_4_M7_g N_Y_c_155_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_54 N_4_M8_g N_Y_c_155_n 4.28653e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_55 N_4_M9_g N_Y_c_155_n 4.28653e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_56 N_4_M10_g N_Y_c_155_n 4.28653e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_57 N_4_M11_g N_Y_c_155_n 4.28653e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_4_M12_g N_Y_c_155_n 4.28653e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_59 N_4_M13_g N_Y_c_155_n 4.28653e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_60 N_4_M14_g N_Y_c_155_n 4.28653e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_61 N_4_M15_g N_Y_c_155_n 4.28653e-19 $X=0.891 $Y=0.0675 $X2=0 $Y2=0
cc_62 N_4_M16_g N_Y_c_155_n 4.28653e-19 $X=0.945 $Y=0.0675 $X2=0 $Y2=0
cc_63 N_4_M17_g N_Y_c_155_n 4.28653e-19 $X=0.999 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_4_M18_g N_Y_c_155_n 4.28653e-19 $X=1.053 $Y=0.0675 $X2=0 $Y2=0
cc_65 N_4_M19_g N_Y_c_155_n 4.28653e-19 $X=1.107 $Y=0.0675 $X2=0 $Y2=0
cc_66 N_4_M20_g N_Y_c_155_n 4.28653e-19 $X=1.161 $Y=0.0675 $X2=0 $Y2=0
cc_67 N_4_M21_g N_Y_c_155_n 4.28653e-19 $X=1.215 $Y=0.0675 $X2=0 $Y2=0
cc_68 N_4_M22_g N_Y_c_155_n 4.28653e-19 $X=1.269 $Y=0.0675 $X2=0 $Y2=0
cc_69 N_4_M23_g N_Y_c_155_n 4.28653e-19 $X=1.323 $Y=0.0675 $X2=0 $Y2=0
cc_70 N_4_M24_g N_Y_c_155_n 4.28653e-19 $X=1.377 $Y=0.0675 $X2=0 $Y2=0
cc_71 N_4_M25_g N_Y_c_155_n 4.28653e-19 $X=1.431 $Y=0.0675 $X2=0 $Y2=0
cc_72 N_4_M26_g N_Y_c_155_n 4.28653e-19 $X=1.485 $Y=0.0675 $X2=0 $Y2=0
cc_73 N_4_M27_g N_Y_c_155_n 4.28653e-19 $X=1.539 $Y=0.0675 $X2=0 $Y2=0
cc_74 N_4_c_30_n N_Y_c_155_n 0.00456243f $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_75 N_4_c_37_n N_Y_c_155_n 4.66342e-19 $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_76 N_4_c_102_p N_Y_c_155_n 0.0168187f $X=0.3305 $Y=0.135 $X2=0 $Y2=0
cc_77 N_4_M5_g N_Y_c_181_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_78 N_4_M6_g N_Y_c_181_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_79 N_4_M7_g N_Y_c_181_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_80 N_4_M8_g N_Y_c_181_n 4.28653e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_81 N_4_M9_g N_Y_c_181_n 4.28653e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_82 N_4_M10_g N_Y_c_181_n 4.28653e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_83 N_4_M11_g N_Y_c_181_n 4.28653e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_84 N_4_M12_g N_Y_c_181_n 4.28653e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_85 N_4_M13_g N_Y_c_181_n 4.28653e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_86 N_4_M14_g N_Y_c_181_n 4.28653e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_87 N_4_M15_g N_Y_c_181_n 4.28653e-19 $X=0.891 $Y=0.0675 $X2=0 $Y2=0
cc_88 N_4_M16_g N_Y_c_181_n 4.28653e-19 $X=0.945 $Y=0.0675 $X2=0 $Y2=0
cc_89 N_4_M17_g N_Y_c_181_n 4.28653e-19 $X=0.999 $Y=0.0675 $X2=0 $Y2=0
cc_90 N_4_M18_g N_Y_c_181_n 4.28653e-19 $X=1.053 $Y=0.0675 $X2=0 $Y2=0
cc_91 N_4_M19_g N_Y_c_181_n 4.28653e-19 $X=1.107 $Y=0.0675 $X2=0 $Y2=0
cc_92 N_4_M20_g N_Y_c_181_n 4.28653e-19 $X=1.161 $Y=0.0675 $X2=0 $Y2=0
cc_93 N_4_M21_g N_Y_c_181_n 4.28653e-19 $X=1.215 $Y=0.0675 $X2=0 $Y2=0
cc_94 N_4_M22_g N_Y_c_181_n 4.28653e-19 $X=1.269 $Y=0.0675 $X2=0 $Y2=0
cc_95 N_4_M23_g N_Y_c_181_n 4.28653e-19 $X=1.323 $Y=0.0675 $X2=0 $Y2=0
cc_96 N_4_M24_g N_Y_c_181_n 4.28653e-19 $X=1.377 $Y=0.0675 $X2=0 $Y2=0
cc_97 N_4_M25_g N_Y_c_181_n 4.28653e-19 $X=1.431 $Y=0.0675 $X2=0 $Y2=0
cc_98 N_4_M26_g N_Y_c_181_n 4.28653e-19 $X=1.485 $Y=0.0675 $X2=0 $Y2=0
cc_99 N_4_M27_g N_Y_c_181_n 4.28653e-19 $X=1.539 $Y=0.0675 $X2=0 $Y2=0
cc_100 N_4_c_30_n N_Y_c_181_n 0.00456243f $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_101 N_4_c_43_n N_Y_c_181_n 4.66342e-19 $X=0.234 $Y=0.234 $X2=0 $Y2=0
cc_102 N_4_c_102_p N_Y_c_181_n 0.0168187f $X=0.3305 $Y=0.135 $X2=0 $Y2=0
cc_103 N_4_c_30_n N_Y_c_207_n 4.48746e-19 $X=1.539 $Y=0.135 $X2=0 $Y2=0
cc_104 N_4_c_130_p N_Y_c_207_n 0.00104492f $X=1.485 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx24_ASAP7_75t_SRAM.pex.sp.BUFX24_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx2_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:19:39 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx2_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx2_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx2_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:19:39 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX2_ASAP7_75T_SRAM%A 2 5 7 15 VSS
c16 15 VSS 0.0121486f $X=0.061 $Y=0.1335
c17 5 VSS 0.00434551f $X=0.081 $Y=0.135
c18 2 VSS 0.0647198f $X=0.081 $Y=0.054
r19 15 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r20 5 19 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r21 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r22 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX2_ASAP7_75T_SRAM%4 2 5 7 10 13 15 17 20 22 25 27 29 34 35 36 38 43
+ 44 46 47 48 51 52 58 61 63 VSS
c29 63 VSS 4.59783e-20 $X=0.111 $Y=0.135
c30 61 VSS 7.83125e-19 $X=0.167 $Y=0.135
c31 60 VSS 8.67243e-19 $X=0.145 $Y=0.135
c32 58 VSS 4.18403e-19 $X=0.189 $Y=0.135
c33 52 VSS 0.00145678f $X=0.111 $Y=0.207
c34 51 VSS 0.00321212f $X=0.111 $Y=0.189
c35 50 VSS 0.00120585f $X=0.111 $Y=0.225
c36 48 VSS 0.00145678f $X=0.111 $Y=0.081
c37 47 VSS 0.00120585f $X=0.111 $Y=0.063
c38 46 VSS 0.00331711f $X=0.111 $Y=0.126
c39 44 VSS 0.00126761f $X=0.0875 $Y=0.234
c40 43 VSS 0.00194817f $X=0.073 $Y=0.234
c41 38 VSS 0.00208886f $X=0.054 $Y=0.234
c42 36 VSS 0.0057867f $X=0.102 $Y=0.234
c43 35 VSS 0.00126761f $X=0.0875 $Y=0.036
c44 34 VSS 0.00194817f $X=0.073 $Y=0.036
c45 29 VSS 0.00208886f $X=0.054 $Y=0.036
c46 27 VSS 0.0057867f $X=0.102 $Y=0.036
c47 25 VSS 0.00694652f $X=0.056 $Y=0.216
c48 22 VSS 2.6657e-19 $X=0.071 $Y=0.216
c49 20 VSS 0.00660761f $X=0.056 $Y=0.054
c50 17 VSS 2.6657e-19 $X=0.071 $Y=0.054
c51 13 VSS 0.00264127f $X=0.189 $Y=0.135
c52 10 VSS 0.0645347f $X=0.189 $Y=0.0675
c53 5 VSS 0.00135968f $X=0.135 $Y=0.135
c54 2 VSS 0.0623485f $X=0.135 $Y=0.0675
r55 60 61 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.145
+ $Y=0.135 $X2=0.167 $Y2=0.135
r56 58 61 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.167 $Y2=0.135
r57 55 60 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.145 $Y2=0.135
r58 53 63 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.12
+ $Y=0.135 $X2=0.111 $Y2=0.135
r59 53 55 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.12
+ $Y=0.135 $X2=0.135 $Y2=0.135
r60 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.189 $X2=0.111 $Y2=0.207
r61 50 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.225 $X2=0.111 $Y2=0.207
r62 49 63 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.144 $X2=0.111 $Y2=0.135
r63 49 51 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.144 $X2=0.111 $Y2=0.189
r64 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.063 $X2=0.111 $Y2=0.081
r65 46 63 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.126 $X2=0.111 $Y2=0.135
r66 46 48 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.126 $X2=0.111 $Y2=0.081
r67 45 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.045 $X2=0.111 $Y2=0.063
r68 43 44 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.073
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r69 38 43 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.073 $Y2=0.234
r70 36 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.102 $Y=0.234 $X2=0.111 $Y2=0.225
r71 36 44 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.102
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r72 34 35 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.073
+ $Y=0.036 $X2=0.0875 $Y2=0.036
r73 29 34 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.073 $Y2=0.036
r74 27 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.102 $Y=0.036 $X2=0.111 $Y2=0.045
r75 27 35 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.102
+ $Y=0.036 $X2=0.0875 $Y2=0.036
r76 25 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r77 22 25 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r78 20 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r79 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r80 13 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r81 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r82 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r83 5 55 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r84 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r85 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_BUFX2_ASAP7_75T_SRAM%Y 1 2 6 7 10 14 16 23 28 29 30 VSS
c13 30 VSS 7.46953e-19 $X=0.243 $Y=0.144
c14 29 VSS 0.00454153f $X=0.243 $Y=0.126
c15 28 VSS 0.00454153f $X=0.244 $Y=0.1495
c16 24 VSS 0.00294383f $X=0.2185 $Y=0.234
c17 23 VSS 0.00543563f $X=0.203 $Y=0.234
c18 18 VSS 0.00579255f $X=0.234 $Y=0.234
c19 17 VSS 0.00294383f $X=0.2185 $Y=0.036
c20 16 VSS 0.00543563f $X=0.203 $Y=0.036
c21 14 VSS 0.0099843f $X=0.162 $Y=0.036
c22 11 VSS 0.00579255f $X=0.234 $Y=0.036
c23 10 VSS 0.00978811f $X=0.162 $Y=0.2025
c24 6 VSS 6.67211e-19 $X=0.179 $Y=0.2025
c25 1 VSS 6.67211e-19 $X=0.179 $Y=0.0675
r26 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.144
r27 28 30 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.1495 $X2=0.243 $Y2=0.144
r28 26 28 5.12654 $w=1.8e-08 $l=7.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.1495
r29 25 29 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.126
r30 23 24 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.203
+ $Y=0.234 $X2=0.2185 $Y2=0.234
r31 20 23 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.203 $Y2=0.234
r32 18 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r33 18 24 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.2185 $Y2=0.234
r34 16 17 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.203
+ $Y=0.036 $X2=0.2185 $Y2=0.036
r35 13 16 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.203 $Y2=0.036
r36 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r37 11 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r38 11 17 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.2185 $Y2=0.036
r39 10 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r40 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r41 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r42 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r43 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.0675 $X2=0.162 $Y2=0.0675
r44 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.162 $Y2=0.0675
.ends


* END of "./BUFx2_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx2_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 VSS N_A_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_4_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 VDD N_A_M3_g N_4_M3_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M4 N_Y_M4_d N_4_M4_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M5 N_Y_M5_d N_4_M5_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
*
* 
* .include "BUFx2_ASAP7_75t_SRAM.pex.sp.BUFX2_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx2_ASAP7_75t_SRAM.pex.sp.BUFX2_ASAP7_75T_SRAM.pxi"
* File: BUFx2_ASAP7_75t_SRAM.pex.sp.BUFX2_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:19:39 2017
* 
x_PM_BUFX2_ASAP7_75T_SRAM%A N_A_M0_g N_A_c_2_p N_A_M3_g A VSS
+ PM_BUFX2_ASAP7_75T_SRAM%A
x_PM_BUFX2_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_18_n N_4_M4_g N_4_M2_g N_4_c_44_p
+ N_4_M5_g N_4_M0_s N_4_c_20_n N_4_M3_s N_4_c_21_n N_4_c_37_p N_4_c_22_n
+ N_4_c_23_n N_4_c_24_n N_4_c_40_p N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_28_n
+ N_4_c_35_p N_4_c_29_n N_4_c_30_n N_4_c_31_n N_4_c_45_p N_4_c_38_p N_4_c_32_n
+ VSS PM_BUFX2_ASAP7_75T_SRAM%4
x_PM_BUFX2_ASAP7_75T_SRAM%Y N_Y_M2_d N_Y_M1_d N_Y_M5_d N_Y_M4_d N_Y_c_46_n
+ N_Y_c_48_n N_Y_c_49_n N_Y_c_52_n Y N_Y_c_56_n N_Y_c_57_n VSS
+ PM_BUFX2_ASAP7_75T_SRAM%Y
cc_1 N_A_M0_g N_4_M1_g 0.00287079f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_4_c_18_n 9.64278e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A_M0_g N_4_M2_g 2.34385e-19 $X=0.081 $Y=0.054 $X2=0.189 $Y2=0.0675
cc_4 A N_4_c_20_n 0.00198071f $X=0.061 $Y=0.1335 $X2=0.056 $Y2=0.054
cc_5 A N_4_c_21_n 0.00198071f $X=0.061 $Y=0.1335 $X2=0.056 $Y2=0.216
cc_6 A N_4_c_22_n 6.00641e-19 $X=0.061 $Y=0.1335 $X2=0.054 $Y2=0.036
cc_7 N_A_c_2_p N_4_c_23_n 2.61546e-19 $X=0.081 $Y=0.135 $X2=0.073 $Y2=0.036
cc_8 N_A_M0_g N_4_c_24_n 3.10016e-19 $X=0.081 $Y=0.054 $X2=0.0875 $Y2=0.036
cc_9 A N_4_c_25_n 6.00641e-19 $X=0.061 $Y=0.1335 $X2=0.054 $Y2=0.234
cc_10 N_A_c_2_p N_4_c_26_n 2.61546e-19 $X=0.081 $Y=0.135 $X2=0.073 $Y2=0.234
cc_11 N_A_M0_g N_4_c_27_n 3.10016e-19 $X=0.081 $Y=0.054 $X2=0.0875 $Y2=0.234
cc_12 A N_4_c_28_n 7.49723e-19 $X=0.061 $Y=0.1335 $X2=0.111 $Y2=0.126
cc_13 A N_4_c_29_n 3.37664e-19 $X=0.061 $Y=0.1335 $X2=0.111 $Y2=0.081
cc_14 A N_4_c_30_n 7.49723e-19 $X=0.061 $Y=0.1335 $X2=0.111 $Y2=0.189
cc_15 A N_4_c_31_n 3.37664e-19 $X=0.061 $Y=0.1335 $X2=0.111 $Y2=0.207
cc_16 A N_4_c_32_n 0.00102244f $X=0.061 $Y=0.1335 $X2=0.111 $Y2=0.135
cc_17 N_4_c_21_n N_Y_c_46_n 2.1777e-19 $X=0.056 $Y=0.216 $X2=0 $Y2=0
cc_18 N_4_c_30_n N_Y_c_46_n 7.34975e-19 $X=0.111 $Y=0.189 $X2=0 $Y2=0
cc_19 N_4_c_35_p N_Y_c_48_n 7.34975e-19 $X=0.111 $Y=0.063 $X2=0 $Y2=0
cc_20 N_4_M2_g N_Y_c_49_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_21 N_4_c_37_p N_Y_c_49_n 0.00114706f $X=0.102 $Y=0.036 $X2=0 $Y2=0
cc_22 N_4_c_38_p N_Y_c_49_n 0.00105983f $X=0.167 $Y=0.135 $X2=0 $Y2=0
cc_23 N_4_M2_g N_Y_c_52_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 N_4_c_40_p N_Y_c_52_n 0.00114706f $X=0.102 $Y=0.234 $X2=0 $Y2=0
cc_25 N_4_c_38_p N_Y_c_52_n 0.00105983f $X=0.167 $Y=0.135 $X2=0 $Y2=0
cc_26 N_4_c_30_n Y 4.97218e-19 $X=0.111 $Y=0.189 $X2=0.081 $Y2=0.135
cc_27 N_4_c_29_n N_Y_c_56_n 4.97218e-19 $X=0.111 $Y=0.081 $X2=0 $Y2=0
cc_28 N_4_c_44_p N_Y_c_57_n 3.15821e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_29 N_4_c_45_p N_Y_c_57_n 0.00103186f $X=0.189 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx2_ASAP7_75t_SRAM.pex.sp.BUFX2_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx3_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:20:02 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx3_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx3_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx3_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:20:02 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX3_ASAP7_75T_SRAM%A 2 5 7 15 VSS
c16 15 VSS 0.0121447f $X=0.061 $Y=0.1335
c17 5 VSS 0.00458972f $X=0.081 $Y=0.135
c18 2 VSS 0.0647198f $X=0.081 $Y=0.0675
r19 15 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r20 5 19 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r21 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX3_ASAP7_75T_SRAM%4 2 5 7 10 15 18 21 23 25 30 33 35 37 38 42 43 44
+ 46 51 52 54 55 56 59 60 69 71 74 VSS
c30 74 VSS 4.62854e-20 $X=0.111 $Y=0.135
c31 71 VSS 0.00161411f $X=0.243 $Y=0.135
c32 69 VSS 7.83125e-19 $X=0.167 $Y=0.135
c33 68 VSS 8.67243e-19 $X=0.145 $Y=0.135
c34 60 VSS 0.00150732f $X=0.111 $Y=0.207
c35 59 VSS 0.0033746f $X=0.111 $Y=0.189
c36 58 VSS 0.00120585f $X=0.111 $Y=0.225
c37 56 VSS 0.00150732f $X=0.111 $Y=0.081
c38 55 VSS 0.00120585f $X=0.111 $Y=0.063
c39 54 VSS 0.00348077f $X=0.111 $Y=0.126
c40 52 VSS 0.00126761f $X=0.0875 $Y=0.234
c41 51 VSS 0.00194782f $X=0.073 $Y=0.234
c42 46 VSS 0.00209231f $X=0.054 $Y=0.234
c43 44 VSS 0.00582115f $X=0.102 $Y=0.234
c44 43 VSS 0.00126761f $X=0.0875 $Y=0.036
c45 42 VSS 0.00194782f $X=0.073 $Y=0.036
c46 38 VSS 0.00635678f $X=0.054 $Y=0.036
c47 37 VSS 0.00209231f $X=0.054 $Y=0.036
c48 35 VSS 0.00582115f $X=0.102 $Y=0.036
c49 33 VSS 0.00635678f $X=0.056 $Y=0.2025
c50 30 VSS 4.5957e-19 $X=0.071 $Y=0.2025
c51 25 VSS 4.5957e-19 $X=0.071 $Y=0.0675
c52 21 VSS 0.00237689f $X=0.243 $Y=0.135
c53 18 VSS 0.0678263f $X=0.243 $Y=0.0675
c54 13 VSS 0.00151182f $X=0.189 $Y=0.135
c55 10 VSS 0.0643964f $X=0.189 $Y=0.0675
c56 5 VSS 0.0012445f $X=0.135 $Y=0.135
c57 2 VSS 0.0621432f $X=0.135 $Y=0.0675
r58 68 69 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.145
+ $Y=0.135 $X2=0.167 $Y2=0.135
r59 66 71 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r60 66 69 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.167 $Y2=0.135
r61 63 68 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.145 $Y2=0.135
r62 61 74 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.12
+ $Y=0.135 $X2=0.111 $Y2=0.135
r63 61 63 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.12
+ $Y=0.135 $X2=0.135 $Y2=0.135
r64 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.189 $X2=0.111 $Y2=0.207
r65 58 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.225 $X2=0.111 $Y2=0.207
r66 57 74 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.144 $X2=0.111 $Y2=0.135
r67 57 59 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.144 $X2=0.111 $Y2=0.189
r68 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.063 $X2=0.111 $Y2=0.081
r69 54 74 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.126 $X2=0.111 $Y2=0.135
r70 54 56 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.126 $X2=0.111 $Y2=0.081
r71 53 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.045 $X2=0.111 $Y2=0.063
r72 51 52 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.073
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r73 46 51 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.073 $Y2=0.234
r74 44 58 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.102 $Y=0.234 $X2=0.111 $Y2=0.225
r75 44 52 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.102
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r76 42 43 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.073
+ $Y=0.036 $X2=0.0875 $Y2=0.036
r77 37 42 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.073 $Y2=0.036
r78 37 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r79 35 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.102 $Y=0.036 $X2=0.111 $Y2=0.045
r80 35 43 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.102
+ $Y=0.036 $X2=0.0875 $Y2=0.036
r81 33 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r82 30 33 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r83 28 38 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r84 25 28 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r85 21 71 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r86 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r87 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r88 13 66 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r89 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r90 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r91 5 63 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r92 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r93 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_BUFX3_ASAP7_75T_SRAM%Y 1 2 6 11 12 15 16 24 29 39 42 44 46 VSS
c14 46 VSS 7.43984e-19 $X=0.297 $Y=0.144
c15 44 VSS 0.00392138f $X=0.2965 $Y=0.1145
c16 42 VSS 0.00392138f $X=0.297 $Y=0.225
c17 40 VSS 4.93225e-19 $X=0.265 $Y=0.234
c18 39 VSS 0.0128846f $X=0.26 $Y=0.234
c19 31 VSS 0.00566632f $X=0.288 $Y=0.234
c20 30 VSS 4.93225e-19 $X=0.265 $Y=0.036
c21 29 VSS 0.0128846f $X=0.26 $Y=0.036
c22 28 VSS 0.00641842f $X=0.27 $Y=0.036
c23 24 VSS 0.00997583f $X=0.162 $Y=0.036
c24 21 VSS 0.00566632f $X=0.288 $Y=0.036
c25 19 VSS 0.00675202f $X=0.268 $Y=0.2025
c26 15 VSS 0.00997583f $X=0.162 $Y=0.2025
c27 11 VSS 6.67211e-19 $X=0.179 $Y=0.2025
c28 9 VSS 3.33606e-19 $X=0.268 $Y=0.0675
c29 1 VSS 6.67211e-19 $X=0.179 $Y=0.0675
r30 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.144
r31 44 45 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1145 $X2=0.297 $Y2=0.126
r32 42 46 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.144
r33 41 44 4.71914 $w=1.8e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.1145
r34 39 40 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.26
+ $Y=0.234 $X2=0.265 $Y2=0.234
r35 37 40 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.265 $Y2=0.234
r36 33 39 6.65432 $w=1.8e-08 $l=9.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.26 $Y2=0.234
r37 31 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.234 $X2=0.297 $Y2=0.225
r38 31 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.27 $Y2=0.234
r39 29 30 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.26
+ $Y=0.036 $X2=0.265 $Y2=0.036
r40 27 30 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.265 $Y2=0.036
r41 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r42 23 29 6.65432 $w=1.8e-08 $l=9.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.26 $Y2=0.036
r43 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r44 21 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r45 21 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.27 $Y2=0.036
r46 19 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r47 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.268 $Y2=0.2025
r48 15 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r49 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r50 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r51 9 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r52 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.268 $Y2=0.0675
r53 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r54 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.0675 $X2=0.162 $Y2=0.0675
r55 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.162 $Y2=0.0675
.ends


* END of "./BUFx3_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx3_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 VSS N_A_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_4_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_4_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 VDD N_A_M4_g N_4_M4_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M5 N_Y_M5_d N_4_M5_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M6 N_Y_M6_d N_4_M6_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M7 N_Y_M7_d N_4_M7_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
*
* 
* .include "BUFx3_ASAP7_75t_SRAM.pex.sp.BUFX3_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx3_ASAP7_75t_SRAM.pex.sp.BUFX3_ASAP7_75T_SRAM.pxi"
* File: BUFx3_ASAP7_75t_SRAM.pex.sp.BUFX3_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:20:02 2017
* 
x_PM_BUFX3_ASAP7_75T_SRAM%A N_A_M0_g N_A_c_2_p N_A_M4_g A VSS
+ PM_BUFX3_ASAP7_75T_SRAM%A
x_PM_BUFX3_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_18_n N_4_M5_g N_4_M2_g N_4_M6_g N_4_M3_g
+ N_4_c_45_p N_4_M7_g N_4_M0_s N_4_M4_s N_4_c_20_n N_4_c_37_p N_4_c_21_n
+ N_4_c_22_n N_4_c_23_n N_4_c_24_n N_4_c_41_p N_4_c_25_n N_4_c_26_n N_4_c_27_n
+ N_4_c_28_n N_4_c_34_p N_4_c_29_n N_4_c_30_n N_4_c_31_n N_4_c_38_p N_4_c_46_p
+ N_4_c_32_n VSS PM_BUFX3_ASAP7_75T_SRAM%4
x_PM_BUFX3_ASAP7_75T_SRAM%Y N_Y_M2_d N_Y_M1_d N_Y_M3_d N_Y_M6_d N_Y_M5_d N_Y_c_47_n
+ N_Y_M7_d N_Y_c_48_n N_Y_c_49_n N_Y_c_53_n N_Y_c_57_n Y N_Y_c_59_n VSS
+ PM_BUFX3_ASAP7_75T_SRAM%Y
cc_1 N_A_M0_g N_4_M1_g 0.00287079f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_4_c_18_n 9.64278e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A_M0_g N_4_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_4 A N_4_c_20_n 0.00198071f $X=0.061 $Y=0.1335 $X2=0.056 $Y2=0.2025
cc_5 A N_4_c_21_n 6.00641e-19 $X=0.061 $Y=0.1335 $X2=0.054 $Y2=0.036
cc_6 A N_4_c_22_n 0.00198071f $X=0.061 $Y=0.1335 $X2=0.054 $Y2=0.036
cc_7 N_A_c_2_p N_4_c_23_n 2.65563e-19 $X=0.081 $Y=0.135 $X2=0.073 $Y2=0.036
cc_8 N_A_M0_g N_4_c_24_n 3.10016e-19 $X=0.081 $Y=0.0675 $X2=0.0875 $Y2=0.036
cc_9 A N_4_c_25_n 6.00641e-19 $X=0.061 $Y=0.1335 $X2=0.054 $Y2=0.234
cc_10 N_A_c_2_p N_4_c_26_n 2.65563e-19 $X=0.081 $Y=0.135 $X2=0.073 $Y2=0.234
cc_11 N_A_M0_g N_4_c_27_n 3.10016e-19 $X=0.081 $Y=0.0675 $X2=0.0875 $Y2=0.234
cc_12 A N_4_c_28_n 7.49723e-19 $X=0.061 $Y=0.1335 $X2=0.111 $Y2=0.126
cc_13 A N_4_c_29_n 3.37664e-19 $X=0.061 $Y=0.1335 $X2=0.111 $Y2=0.081
cc_14 A N_4_c_30_n 7.49723e-19 $X=0.061 $Y=0.1335 $X2=0.111 $Y2=0.189
cc_15 A N_4_c_31_n 3.37664e-19 $X=0.061 $Y=0.1335 $X2=0.111 $Y2=0.207
cc_16 A N_4_c_32_n 0.0010383f $X=0.061 $Y=0.1335 $X2=0.111 $Y2=0.135
cc_17 N_4_c_30_n N_Y_c_47_n 8.06181e-19 $X=0.111 $Y=0.189 $X2=0.061 $Y2=0.1335
cc_18 N_4_c_34_p N_Y_c_48_n 8.06181e-19 $X=0.111 $Y=0.063 $X2=0 $Y2=0
cc_19 N_4_M2_g N_Y_c_49_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_20 N_4_M3_g N_Y_c_49_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_21 N_4_c_37_p N_Y_c_49_n 0.00116333f $X=0.102 $Y=0.036 $X2=0 $Y2=0
cc_22 N_4_c_38_p N_Y_c_49_n 0.00211774f $X=0.167 $Y=0.135 $X2=0 $Y2=0
cc_23 N_4_M2_g N_Y_c_53_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 N_4_M3_g N_Y_c_53_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_25 N_4_c_41_p N_Y_c_53_n 0.00116333f $X=0.102 $Y=0.234 $X2=0 $Y2=0
cc_26 N_4_c_38_p N_Y_c_53_n 0.00211774f $X=0.167 $Y=0.135 $X2=0 $Y2=0
cc_27 N_4_c_30_n N_Y_c_57_n 2.81016e-19 $X=0.111 $Y=0.189 $X2=0 $Y2=0
cc_28 N_4_c_29_n Y 2.81016e-19 $X=0.111 $Y=0.081 $X2=0 $Y2=0
cc_29 N_4_c_45_p N_Y_c_59_n 3.12222e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_30 N_4_c_46_p N_Y_c_59_n 0.00113929f $X=0.243 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx3_ASAP7_75t_SRAM.pex.sp.BUFX3_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx4_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:20:24 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx4_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx4_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx4_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:20:24 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX4_ASAP7_75T_SRAM%A 2 5 7 15 VSS
c16 15 VSS 0.012159f $X=0.061 $Y=0.1355
c17 5 VSS 0.00434738f $X=0.081 $Y=0.135
c18 2 VSS 0.0647198f $X=0.081 $Y=0.054
r19 15 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r20 5 19 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r21 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r22 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX4_ASAP7_75T_SRAM%4 2 5 7 10 15 18 23 26 29 31 33 36 38 41 43 45 50
+ 51 52 54 59 60 62 63 64 67 68 77 82 85 VSS
c31 85 VSS 4.64886e-20 $X=0.111 $Y=0.135
c32 82 VSS 0.00249105f $X=0.297 $Y=0.135
c33 77 VSS 7.83125e-19 $X=0.167 $Y=0.135
c34 76 VSS 8.67243e-19 $X=0.145 $Y=0.135
c35 68 VSS 0.00159137f $X=0.111 $Y=0.207
c36 67 VSS 0.00367238f $X=0.111 $Y=0.189
c37 66 VSS 0.00120585f $X=0.111 $Y=0.225
c38 64 VSS 0.00159137f $X=0.111 $Y=0.081
c39 63 VSS 0.00120585f $X=0.111 $Y=0.063
c40 62 VSS 0.00377913f $X=0.111 $Y=0.126
c41 60 VSS 0.00126761f $X=0.0875 $Y=0.234
c42 59 VSS 0.00195257f $X=0.073 $Y=0.234
c43 54 VSS 0.00209231f $X=0.054 $Y=0.234
c44 52 VSS 0.0057943f $X=0.102 $Y=0.234
c45 51 VSS 0.00126761f $X=0.0875 $Y=0.036
c46 50 VSS 0.00195257f $X=0.073 $Y=0.036
c47 45 VSS 0.00209231f $X=0.054 $Y=0.036
c48 43 VSS 0.0057943f $X=0.102 $Y=0.036
c49 41 VSS 0.00694652f $X=0.056 $Y=0.216
c50 38 VSS 2.6657e-19 $X=0.071 $Y=0.216
c51 36 VSS 0.00660761f $X=0.056 $Y=0.054
c52 33 VSS 2.6657e-19 $X=0.071 $Y=0.054
c53 29 VSS 0.00242908f $X=0.297 $Y=0.135
c54 26 VSS 0.0645347f $X=0.297 $Y=0.0675
c55 21 VSS 0.00123791f $X=0.243 $Y=0.135
c56 18 VSS 0.0644226f $X=0.243 $Y=0.0675
c57 13 VSS 0.00116657f $X=0.189 $Y=0.135
c58 10 VSS 0.0642127f $X=0.189 $Y=0.0675
c59 5 VSS 0.0012445f $X=0.135 $Y=0.135
c60 2 VSS 0.0621464f $X=0.135 $Y=0.0675
r61 79 82 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r62 76 77 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.145
+ $Y=0.135 $X2=0.167 $Y2=0.135
r63 74 79 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r64 74 77 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.167 $Y2=0.135
r65 71 76 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.145 $Y2=0.135
r66 69 85 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.12
+ $Y=0.135 $X2=0.111 $Y2=0.135
r67 69 71 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.12
+ $Y=0.135 $X2=0.135 $Y2=0.135
r68 67 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.189 $X2=0.111 $Y2=0.207
r69 66 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.225 $X2=0.111 $Y2=0.207
r70 65 85 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.144 $X2=0.111 $Y2=0.135
r71 65 67 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.144 $X2=0.111 $Y2=0.189
r72 63 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.063 $X2=0.111 $Y2=0.081
r73 62 85 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.126 $X2=0.111 $Y2=0.135
r74 62 64 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.126 $X2=0.111 $Y2=0.081
r75 61 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.045 $X2=0.111 $Y2=0.063
r76 59 60 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.073
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r77 54 59 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.073 $Y2=0.234
r78 52 66 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.102 $Y=0.234 $X2=0.111 $Y2=0.225
r79 52 60 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.102
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r80 50 51 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.073
+ $Y=0.036 $X2=0.0875 $Y2=0.036
r81 45 50 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.073 $Y2=0.036
r82 43 61 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.102 $Y=0.036 $X2=0.111 $Y2=0.045
r83 43 51 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.102
+ $Y=0.036 $X2=0.0875 $Y2=0.036
r84 41 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r85 38 41 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r86 36 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r87 33 36 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r88 29 82 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r89 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r90 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r91 21 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r92 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r93 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r94 13 74 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r95 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r96 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r97 5 71 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r98 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r99 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_BUFX4_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 15 16 17 24 29 39 44 46 VSS
c15 46 VSS 7.58018e-19 $X=0.348 $Y=0.144
c16 44 VSS 0.00597441f $X=0.3515 $Y=0.1145
c17 42 VSS 0.00597441f $X=0.348 $Y=0.225
c18 40 VSS 0.00211927f $X=0.3265 $Y=0.234
c19 39 VSS 0.0179375f $X=0.314 $Y=0.234
c20 31 VSS 0.00538136f $X=0.339 $Y=0.234
c21 30 VSS 0.00211927f $X=0.3265 $Y=0.036
c22 29 VSS 0.0179375f $X=0.314 $Y=0.036
c23 28 VSS 0.00888988f $X=0.27 $Y=0.036
c24 24 VSS 0.00997633f $X=0.162 $Y=0.036
c25 21 VSS 0.00538136f $X=0.339 $Y=0.036
c26 20 VSS 0.00888988f $X=0.27 $Y=0.2025
c27 16 VSS 6.67211e-19 $X=0.287 $Y=0.2025
c28 15 VSS 0.00978014f $X=0.162 $Y=0.2025
c29 11 VSS 6.67211e-19 $X=0.179 $Y=0.2025
c30 6 VSS 6.67211e-19 $X=0.287 $Y=0.0675
c31 1 VSS 6.67211e-19 $X=0.179 $Y=0.0675
r32 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.348
+ $Y=0.126 $X2=0.348 $Y2=0.144
r33 44 45 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.348
+ $Y=0.1145 $X2=0.348 $Y2=0.126
r34 42 46 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.348
+ $Y=0.225 $X2=0.348 $Y2=0.144
r35 41 44 4.71914 $w=1.8e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.348
+ $Y=0.045 $X2=0.348 $Y2=0.1145
r36 39 40 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.314
+ $Y=0.234 $X2=0.3265 $Y2=0.234
r37 37 39 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.314 $Y2=0.234
r38 33 37 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.27 $Y2=0.234
r39 31 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.339 $Y=0.234 $X2=0.348 $Y2=0.225
r40 31 40 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.339
+ $Y=0.234 $X2=0.3265 $Y2=0.234
r41 29 30 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.314
+ $Y=0.036 $X2=0.3265 $Y2=0.036
r42 27 29 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.314 $Y2=0.036
r43 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r44 23 27 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.27 $Y2=0.036
r45 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r46 21 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.339 $Y=0.036 $X2=0.348 $Y2=0.045
r47 21 30 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.339
+ $Y=0.036 $X2=0.3265 $Y2=0.036
r48 20 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r49 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r50 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r51 15 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r52 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r53 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r54 10 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r55 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r56 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r57 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r58 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.0675 $X2=0.162 $Y2=0.0675
r59 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.162 $Y2=0.0675
.ends


* END of "./BUFx4_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx4_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 VSS N_A_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_4_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_4_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 VDD N_A_M5_g N_4_M5_s VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M6 N_Y_M6_d N_4_M6_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M7 N_Y_M7_d N_4_M7_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M8 N_Y_M8_d N_4_M8_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M9 N_Y_M9_d N_4_M9_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
*
* 
* .include "BUFx4_ASAP7_75t_SRAM.pex.sp.BUFX4_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx4_ASAP7_75t_SRAM.pex.sp.BUFX4_ASAP7_75T_SRAM.pxi"
* File: BUFx4_ASAP7_75t_SRAM.pex.sp.BUFX4_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:20:24 2017
* 
x_PM_BUFX4_ASAP7_75T_SRAM%A N_A_M0_g N_A_c_2_p N_A_M5_g A VSS
+ PM_BUFX4_ASAP7_75T_SRAM%A
x_PM_BUFX4_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_18_n N_4_M6_g N_4_M2_g N_4_M7_g N_4_M3_g
+ N_4_M8_g N_4_M4_g N_4_c_46_p N_4_M9_g N_4_M0_s N_4_c_20_n N_4_M5_s N_4_c_21_n
+ N_4_c_39_p N_4_c_22_n N_4_c_23_n N_4_c_24_n N_4_c_44_p N_4_c_25_n N_4_c_26_n
+ N_4_c_27_n N_4_c_28_n N_4_c_35_p N_4_c_29_n N_4_c_30_n N_4_c_31_n N_4_c_40_p
+ N_4_c_47_p N_4_c_32_n VSS PM_BUFX4_ASAP7_75T_SRAM%4
x_PM_BUFX4_ASAP7_75T_SRAM%Y N_Y_M2_d N_Y_M1_d N_Y_M4_d N_Y_M3_d N_Y_M7_d N_Y_M6_d
+ N_Y_c_48_n N_Y_M9_d N_Y_M8_d N_Y_c_50_n N_Y_c_51_n N_Y_c_56_n Y N_Y_c_61_n VSS
+ PM_BUFX4_ASAP7_75T_SRAM%Y
cc_1 N_A_M0_g N_4_M1_g 0.00287079f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_4_c_18_n 9.64278e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A_M0_g N_4_M2_g 2.34385e-19 $X=0.081 $Y=0.054 $X2=0.189 $Y2=0.0675
cc_4 A N_4_c_20_n 0.00198071f $X=0.061 $Y=0.1355 $X2=0.056 $Y2=0.054
cc_5 A N_4_c_21_n 0.00198071f $X=0.061 $Y=0.1355 $X2=0.056 $Y2=0.216
cc_6 A N_4_c_22_n 6.00641e-19 $X=0.061 $Y=0.1355 $X2=0.054 $Y2=0.036
cc_7 N_A_c_2_p N_4_c_23_n 2.65563e-19 $X=0.081 $Y=0.135 $X2=0.073 $Y2=0.036
cc_8 N_A_M0_g N_4_c_24_n 3.10016e-19 $X=0.081 $Y=0.054 $X2=0.0875 $Y2=0.036
cc_9 A N_4_c_25_n 6.00641e-19 $X=0.061 $Y=0.1355 $X2=0.054 $Y2=0.234
cc_10 N_A_c_2_p N_4_c_26_n 2.65563e-19 $X=0.081 $Y=0.135 $X2=0.073 $Y2=0.234
cc_11 N_A_M0_g N_4_c_27_n 3.10016e-19 $X=0.081 $Y=0.054 $X2=0.0875 $Y2=0.234
cc_12 A N_4_c_28_n 7.49723e-19 $X=0.061 $Y=0.1355 $X2=0.111 $Y2=0.126
cc_13 A N_4_c_29_n 3.37664e-19 $X=0.061 $Y=0.1355 $X2=0.111 $Y2=0.081
cc_14 A N_4_c_30_n 7.49723e-19 $X=0.061 $Y=0.1355 $X2=0.111 $Y2=0.189
cc_15 A N_4_c_31_n 3.37664e-19 $X=0.061 $Y=0.1355 $X2=0.111 $Y2=0.207
cc_16 A N_4_c_32_n 0.00104452f $X=0.061 $Y=0.1355 $X2=0.111 $Y2=0.135
cc_17 N_4_c_21_n N_Y_c_48_n 2.1777e-19 $X=0.056 $Y=0.216 $X2=0.061 $Y2=0.1355
cc_18 N_4_c_30_n N_Y_c_48_n 0.00112297f $X=0.111 $Y=0.189 $X2=0.061 $Y2=0.1355
cc_19 N_4_c_35_p N_Y_c_50_n 0.00112297f $X=0.111 $Y=0.063 $X2=0 $Y2=0
cc_20 N_4_M2_g N_Y_c_51_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_21 N_4_M3_g N_Y_c_51_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_22 N_4_M4_g N_Y_c_51_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_23 N_4_c_39_p N_Y_c_51_n 0.00116998f $X=0.102 $Y=0.036 $X2=0 $Y2=0
cc_24 N_4_c_40_p N_Y_c_51_n 0.00310217f $X=0.167 $Y=0.135 $X2=0 $Y2=0
cc_25 N_4_M2_g N_Y_c_56_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_4_M3_g N_Y_c_56_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_4_M4_g N_Y_c_56_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_28 N_4_c_44_p N_Y_c_56_n 0.00116998f $X=0.102 $Y=0.234 $X2=0 $Y2=0
cc_29 N_4_c_40_p N_Y_c_56_n 0.00310217f $X=0.167 $Y=0.135 $X2=0 $Y2=0
cc_30 N_4_c_46_p N_Y_c_61_n 3.37735e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_31 N_4_c_47_p N_Y_c_61_n 0.00127049f $X=0.297 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx4_ASAP7_75t_SRAM.pex.sp.BUFX4_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx4f_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:20:46 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx4f_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx4f_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx4f_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:20:46 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX4F_ASAP7_75T_SRAM%A 2 7 10 13 15 23 VSS
c19 23 VSS 0.0256137f $X=0.081 $Y=0.135
c20 13 VSS 0.00864439f $X=0.135 $Y=0.135
c21 10 VSS 0.0611086f $X=0.135 $Y=0.0675
c22 2 VSS 0.0654907f $X=0.081 $Y=0.0405
r23 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r24 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r25 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r26 5 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r27 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2295
r28 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0405 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX4F_ASAP7_75T_SRAM%4 2 7 10 15 18 23 26 29 31 33 39 41 45 47 50 52 57
+ 58 60 64 65 69 74 79 83 VSS
c37 80 VSS 0.00199291f $X=0.126 $Y=0.234
c38 79 VSS 0.00263626f $X=0.135 $Y=0.234
c39 74 VSS 0.00209909f $X=0.108 $Y=0.234
c40 70 VSS 0.00199291f $X=0.126 $Y=0.036
c41 69 VSS 0.00263626f $X=0.135 $Y=0.036
c42 65 VSS 0.0107924f $X=0.108 $Y=0.036
c43 64 VSS 0.00209909f $X=0.108 $Y=0.036
c44 60 VSS 2.78189e-19 $X=0.351 $Y=0.135
c45 57 VSS 0.00271998f $X=0.199 $Y=0.135
c46 52 VSS 0.00385172f $X=0.135 $Y=0.225
c47 50 VSS 0.00385172f $X=0.135 $Y=0.126
c48 48 VSS 5.36734e-19 $X=0.108 $Y=0.2295
c49 45 VSS 0.0107924f $X=0.108 $Y=0.2025
c50 42 VSS 0.00368068f $X=0.1125 $Y=0.216
c51 40 VSS 5.36734e-19 $X=0.108 $Y=0.0405
c52 34 VSS 0.00368068f $X=0.1125 $Y=0.054
c53 29 VSS 0.0121429f $X=0.351 $Y=0.135
c54 26 VSS 0.0645347f $X=0.351 $Y=0.0675
c55 18 VSS 0.0644226f $X=0.297 $Y=0.0675
c56 10 VSS 0.0642127f $X=0.243 $Y=0.0675
c57 2 VSS 0.0620458f $X=0.189 $Y=0.0675
r58 80 81 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r59 79 81 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r60 74 80 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r61 70 71 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r62 69 71 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r63 64 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r64 64 65 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r65 57 58 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.199
+ $Y=0.135 $X2=0.221 $Y2=0.135
r66 55 60 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.351 $Y2=0.135
r67 55 58 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.221 $Y2=0.135
r68 53 83 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.135 $Y2=0.135
r69 53 57 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.199 $Y2=0.135
r70 52 79 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.234
r71 51 83 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.135
r72 51 52 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.225
r73 50 83 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.135
r74 49 69 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.036
r75 49 50 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.126
r76 47 48 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2295 $X2=0.108 $Y2=0.2295
r77 45 74 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r78 42 48 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1125 $Y=0.216 $X2=0.108 $Y2=0.2295
r79 42 45 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.1125 $Y=0.216 $X2=0.1125 $Y2=0.189
r80 41 45 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.189 $X2=0.1125 $Y2=0.189
r81 39 40 15.8795 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0405 $X2=0.108 $Y2=0.0405
r82 37 65 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r83 34 40 5.31511 $w=5.4e-08 $l=1.55885e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1125 $Y=0.054 $X2=0.108 $Y2=0.0405
r84 34 37 18.1206 $w=5.4e-08 $l=2.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.1125 $Y=0.054 $X2=0.1125 $Y2=0.081
r85 33 37 8.38915 $w=5.4e-08 $l=1.25e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.081 $X2=0.1125 $Y2=0.081
r86 29 60 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r87 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r88 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r89 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r90 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r91 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r92 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r93 13 55 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r94 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r95 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r96 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r97 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r98 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_BUFX4F_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 29 39 44 46 VSS
c18 46 VSS 7.43984e-19 $X=0.405 $Y=0.144
c19 45 VSS 0.00538213f $X=0.405 $Y=0.126
c20 44 VSS 0.00538213f $X=0.406 $Y=0.153
c21 40 VSS 0.00247117f $X=0.3815 $Y=0.234
c22 39 VSS 0.0177808f $X=0.367 $Y=0.234
c23 31 VSS 0.00566315f $X=0.396 $Y=0.234
c24 30 VSS 0.00247117f $X=0.3815 $Y=0.036
c25 29 VSS 0.0177808f $X=0.367 $Y=0.036
c26 28 VSS 0.00929752f $X=0.324 $Y=0.036
c27 24 VSS 0.00916652f $X=0.216 $Y=0.036
c28 21 VSS 0.00566315f $X=0.396 $Y=0.036
c29 20 VSS 0.00929752f $X=0.324 $Y=0.2025
c30 16 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c31 15 VSS 0.00916652f $X=0.216 $Y=0.2025
c32 11 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c33 6 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c34 1 VSS 5.38922e-19 $X=0.233 $Y=0.0675
r35 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.126 $X2=0.405 $Y2=0.144
r36 44 46 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.153 $X2=0.405 $Y2=0.144
r37 42 44 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.153
r38 41 45 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.126
r39 39 40 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.234 $X2=0.3815 $Y2=0.234
r40 37 39 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.367 $Y2=0.234
r41 33 37 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.324 $Y2=0.234
r42 31 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r43 31 40 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.3815 $Y2=0.234
r44 29 30 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.367
+ $Y=0.036 $X2=0.3815 $Y2=0.036
r45 27 29 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.367 $Y2=0.036
r46 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r47 23 27 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.324 $Y2=0.036
r48 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r49 21 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r50 21 30 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.3815 $Y2=0.036
r51 20 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r52 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r53 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r54 15 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r55 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r56 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r57 10 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r58 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r59 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r60 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r61 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r62 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./BUFx4f_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx4f_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_4_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071 $Y=0.027
M1 N_4_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_4_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_4_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_4_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_4_M6_d N_A_M6_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071 $Y=0.216
M7 N_4_M7_d N_A_M7_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M8 N_Y_M8_d N_4_M8_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M9 N_Y_M9_d N_4_M9_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M10 N_Y_M10_d N_4_M10_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_Y_M11_d N_4_M11_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "BUFx4f_ASAP7_75t_SRAM.pex.sp.BUFX4F_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx4f_ASAP7_75t_SRAM.pex.sp.BUFX4F_ASAP7_75T_SRAM.pxi"
* File: BUFx4f_ASAP7_75t_SRAM.pex.sp.BUFX4F_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:20:46 2017
* 
x_PM_BUFX4F_ASAP7_75T_SRAM%A N_A_M0_g N_A_M6_g N_A_M1_g N_A_c_4_p N_A_M7_g A VSS
+ PM_BUFX4F_ASAP7_75T_SRAM%A
x_PM_BUFX4F_ASAP7_75T_SRAM%4 N_4_M2_g N_4_M8_g N_4_M3_g N_4_M9_g N_4_M4_g N_4_M10_g
+ N_4_M5_g N_4_c_23_n N_4_M11_g N_4_M1_d N_4_M0_d N_4_M7_d N_4_c_24_n N_4_M6_d
+ N_4_c_25_n N_4_c_28_n N_4_c_31_n N_4_c_47_p N_4_c_56_p N_4_c_32_n N_4_c_34_n
+ N_4_c_48_p N_4_c_35_n N_4_c_54_p N_4_c_37_n VSS PM_BUFX4F_ASAP7_75T_SRAM%4
x_PM_BUFX4F_ASAP7_75T_SRAM%Y N_Y_M3_d N_Y_M2_d N_Y_M5_d N_Y_M4_d N_Y_M9_d N_Y_M8_d
+ N_Y_M11_d N_Y_M10_d N_Y_c_61_n N_Y_c_67_n Y N_Y_c_73_n VSS
+ PM_BUFX4F_ASAP7_75T_SRAM%Y
cc_1 N_A_M0_g N_4_M2_g 2.34385e-19 $X=0.081 $Y=0.0405 $X2=0.189 $Y2=0.0675
cc_2 N_A_M1_g N_4_M2_g 0.00287079f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A_M1_g N_4_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_4 N_A_c_4_p N_4_c_23_n 0.00154475f $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.135
cc_5 N_A_c_4_p N_4_c_24_n 7.33389e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_6 N_A_M1_g N_4_c_25_n 6.45702e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.126
cc_7 N_A_c_4_p N_4_c_25_n 4.76064e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.126
cc_8 A N_4_c_25_n 6.94026e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.126
cc_9 N_A_M1_g N_4_c_28_n 6.45702e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.225
cc_10 N_A_c_4_p N_4_c_28_n 4.76064e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.225
cc_11 A N_4_c_28_n 6.94026e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.225
cc_12 N_A_c_4_p N_4_c_31_n 4.61514e-19 $X=0.135 $Y=0.135 $X2=0.199 $Y2=0.135
cc_13 N_A_c_4_p N_4_c_32_n 3.42441e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.036
cc_14 A N_4_c_32_n 5.37037e-19 $X=0.081 $Y=0.135 $X2=0.108 $Y2=0.036
cc_15 N_A_c_4_p N_4_c_34_n 7.33389e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.036
cc_16 N_A_c_4_p N_4_c_35_n 3.42441e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.234
cc_17 A N_4_c_35_n 5.37037e-19 $X=0.081 $Y=0.135 $X2=0.108 $Y2=0.234
cc_18 N_A_c_4_p N_4_c_37_n 0.00101232f $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.135
cc_19 A N_4_c_37_n 0.00105383f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_20 N_4_c_23_n N_Y_M3_d 3.80218e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.0405
cc_21 N_4_c_23_n N_Y_M5_d 3.80218e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.2295
cc_22 N_4_c_23_n N_Y_M9_d 3.80218e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_23 N_4_c_23_n N_Y_M11_d 3.80218e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_24 N_4_M3_g N_Y_c_61_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_25 N_4_M4_g N_Y_c_61_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_4_M5_g N_Y_c_61_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_4_c_23_n N_Y_c_61_n 6.45396e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_28 N_4_c_47_p N_Y_c_61_n 0.0023383f $X=0.221 $Y=0.135 $X2=0 $Y2=0
cc_29 N_4_c_48_p N_Y_c_61_n 3.90464e-19 $X=0.135 $Y=0.036 $X2=0 $Y2=0
cc_30 N_4_M3_g N_Y_c_67_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_4_M4_g N_Y_c_67_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_32 N_4_M5_g N_Y_c_67_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_33 N_4_c_23_n N_Y_c_67_n 6.45396e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_34 N_4_c_47_p N_Y_c_67_n 0.0023383f $X=0.221 $Y=0.135 $X2=0 $Y2=0
cc_35 N_4_c_54_p N_Y_c_67_n 3.90464e-19 $X=0.135 $Y=0.234 $X2=0 $Y2=0
cc_36 N_4_c_23_n N_Y_c_73_n 4.93118e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_56_p N_Y_c_73_n 0.00110084f $X=0.351 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx4f_ASAP7_75t_SRAM.pex.sp.BUFX4F_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx5_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:21:09 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx5_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx5_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx5_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:21:09 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX5_ASAP7_75T_SRAM%A 2 5 7 15 VSS
c16 15 VSS 0.0121447f $X=0.061 $Y=0.1365
c17 5 VSS 0.00459073f $X=0.081 $Y=0.135
c18 2 VSS 0.0647198f $X=0.081 $Y=0.0675
r19 15 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r20 5 19 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r21 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX5_ASAP7_75T_SRAM%4 2 5 7 10 15 18 23 26 31 34 37 39 41 46 49 51 53
+ 54 58 59 60 62 67 68 70 71 72 75 76 85 93 96 VSS
c32 96 VSS 4.66463e-20 $X=0.111 $Y=0.135
c33 93 VSS 0.00356617f $X=0.351 $Y=0.135
c34 85 VSS 7.83125e-19 $X=0.167 $Y=0.135
c35 84 VSS 8.67243e-19 $X=0.145 $Y=0.135
c36 76 VSS 0.00159137f $X=0.111 $Y=0.207
c37 75 VSS 0.00367238f $X=0.111 $Y=0.189
c38 74 VSS 0.00120585f $X=0.111 $Y=0.225
c39 72 VSS 0.00159137f $X=0.111 $Y=0.081
c40 71 VSS 0.00120585f $X=0.111 $Y=0.063
c41 70 VSS 0.0037795f $X=0.111 $Y=0.126
c42 68 VSS 0.00126761f $X=0.0875 $Y=0.234
c43 67 VSS 0.00194782f $X=0.073 $Y=0.234
c44 62 VSS 0.00209231f $X=0.054 $Y=0.234
c45 60 VSS 0.00582115f $X=0.102 $Y=0.234
c46 59 VSS 0.00126761f $X=0.0875 $Y=0.036
c47 58 VSS 0.00194782f $X=0.073 $Y=0.036
c48 54 VSS 0.00635678f $X=0.054 $Y=0.036
c49 53 VSS 0.00209231f $X=0.054 $Y=0.036
c50 51 VSS 0.00582115f $X=0.102 $Y=0.036
c51 49 VSS 0.00635678f $X=0.056 $Y=0.2025
c52 46 VSS 4.5957e-19 $X=0.071 $Y=0.2025
c53 41 VSS 4.5957e-19 $X=0.071 $Y=0.0675
c54 37 VSS 0.00241526f $X=0.351 $Y=0.135
c55 34 VSS 0.0678263f $X=0.351 $Y=0.0675
c56 29 VSS 0.00123791f $X=0.297 $Y=0.135
c57 26 VSS 0.0643964f $X=0.297 $Y=0.0675
c58 21 VSS 0.00112752f $X=0.243 $Y=0.135
c59 18 VSS 0.0642127f $X=0.243 $Y=0.0675
c60 13 VSS 0.00116657f $X=0.189 $Y=0.135
c61 10 VSS 0.0642127f $X=0.189 $Y=0.0675
c62 5 VSS 0.0012445f $X=0.135 $Y=0.135
c63 2 VSS 0.0621491f $X=0.135 $Y=0.0675
r64 90 93 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r65 87 90 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r66 84 85 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.145
+ $Y=0.135 $X2=0.167 $Y2=0.135
r67 82 87 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r68 82 85 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.167 $Y2=0.135
r69 79 84 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.145 $Y2=0.135
r70 77 96 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.12
+ $Y=0.135 $X2=0.111 $Y2=0.135
r71 77 79 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.12
+ $Y=0.135 $X2=0.135 $Y2=0.135
r72 75 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.189 $X2=0.111 $Y2=0.207
r73 74 76 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.225 $X2=0.111 $Y2=0.207
r74 73 96 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.144 $X2=0.111 $Y2=0.135
r75 73 75 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.144 $X2=0.111 $Y2=0.189
r76 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.063 $X2=0.111 $Y2=0.081
r77 70 96 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.126 $X2=0.111 $Y2=0.135
r78 70 72 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.126 $X2=0.111 $Y2=0.081
r79 69 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.111
+ $Y=0.045 $X2=0.111 $Y2=0.063
r80 67 68 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.073
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r81 62 67 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.073 $Y2=0.234
r82 60 74 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.102 $Y=0.234 $X2=0.111 $Y2=0.225
r83 60 68 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.102
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r84 58 59 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.073
+ $Y=0.036 $X2=0.0875 $Y2=0.036
r85 53 58 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.073 $Y2=0.036
r86 53 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r87 51 69 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.102 $Y=0.036 $X2=0.111 $Y2=0.045
r88 51 59 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.102
+ $Y=0.036 $X2=0.0875 $Y2=0.036
r89 49 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r90 46 49 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r91 44 54 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r92 41 44 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r93 37 93 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r94 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r95 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r96 29 90 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r97 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r98 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r99 21 87 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r100 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.2025
r101 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.135
r102 13 82 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r103 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.189 $Y=0.135 $X2=0.189 $Y2=0.2025
r104 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.189 $Y=0.0675 $X2=0.189 $Y2=0.135
r105 5 79 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r106 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r107 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_BUFX5_ASAP7_75T_SRAM%Y 1 2 6 7 11 16 17 20 21 22 26 34 42 55 60 62 VSS
c16 62 VSS 7.43984e-19 $X=0.405 $Y=0.144
c17 60 VSS 0.00406168f $X=0.4075 $Y=0.1145
c18 58 VSS 0.00406168f $X=0.405 $Y=0.225
c19 56 VSS 4.93225e-19 $X=0.373 $Y=0.234
c20 55 VSS 0.024627f $X=0.368 $Y=0.234
c21 44 VSS 0.0056949f $X=0.396 $Y=0.234
c22 43 VSS 4.93225e-19 $X=0.373 $Y=0.036
c23 42 VSS 0.024627f $X=0.368 $Y=0.036
c24 41 VSS 0.00641842f $X=0.378 $Y=0.036
c25 38 VSS 0.00888469f $X=0.27 $Y=0.036
c26 34 VSS 0.00997633f $X=0.162 $Y=0.036
c27 31 VSS 0.0056949f $X=0.396 $Y=0.036
c28 29 VSS 0.00675202f $X=0.376 $Y=0.2025
c29 25 VSS 0.00888469f $X=0.27 $Y=0.2025
c30 21 VSS 6.67211e-19 $X=0.287 $Y=0.2025
c31 20 VSS 0.00997633f $X=0.162 $Y=0.2025
c32 16 VSS 6.67211e-19 $X=0.179 $Y=0.2025
c33 14 VSS 3.33606e-19 $X=0.376 $Y=0.0675
c34 6 VSS 6.67211e-19 $X=0.287 $Y=0.0675
c35 1 VSS 6.67211e-19 $X=0.179 $Y=0.0675
r36 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.126 $X2=0.405 $Y2=0.144
r37 60 61 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.1145 $X2=0.405 $Y2=0.126
r38 58 62 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.144
r39 57 60 4.71914 $w=1.8e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.1145
r40 55 56 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.368
+ $Y=0.234 $X2=0.373 $Y2=0.234
r41 53 56 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.373 $Y2=0.234
r42 50 55 6.65432 $w=1.8e-08 $l=9.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.368 $Y2=0.234
r43 46 50 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.27 $Y2=0.234
r44 44 58 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r45 44 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.378 $Y2=0.234
r46 42 43 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.368
+ $Y=0.036 $X2=0.373 $Y2=0.036
r47 40 43 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.373 $Y2=0.036
r48 40 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r49 37 42 6.65432 $w=1.8e-08 $l=9.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.368 $Y2=0.036
r50 37 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r51 33 37 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.27 $Y2=0.036
r52 33 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r53 31 57 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r54 31 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.378 $Y2=0.036
r55 29 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r56 26 29 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.376 $Y2=0.2025
r57 25 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r58 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r59 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r60 20 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r61 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r62 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r63 14 41 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r64 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.376 $Y2=0.0675
r65 10 38 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r66 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r67 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r68 5 34 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r69 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.0675 $X2=0.162 $Y2=0.0675
r70 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.162 $Y2=0.0675
.ends


* END of "./BUFx5_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx5_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 VSS N_A_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_4_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_4_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_4_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 VDD N_A_M6_g N_4_M6_s VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M7 N_Y_M7_d N_4_M7_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M8 N_Y_M8_d N_4_M8_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M9 N_Y_M9_d N_4_M9_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M10 N_Y_M10_d N_4_M10_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_Y_M11_d N_4_M11_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "BUFx5_ASAP7_75t_SRAM.pex.sp.BUFX5_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx5_ASAP7_75t_SRAM.pex.sp.BUFX5_ASAP7_75T_SRAM.pxi"
* File: BUFx5_ASAP7_75t_SRAM.pex.sp.BUFX5_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:21:09 2017
* 
x_PM_BUFX5_ASAP7_75T_SRAM%A N_A_M0_g N_A_c_2_p N_A_M6_g A VSS
+ PM_BUFX5_ASAP7_75T_SRAM%A
x_PM_BUFX5_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_18_n N_4_M7_g N_4_M2_g N_4_M8_g N_4_M3_g
+ N_4_M9_g N_4_M4_g N_4_M10_g N_4_M5_g N_4_c_47_p N_4_M11_g N_4_M0_s N_4_M6_s
+ N_4_c_20_n N_4_c_39_p N_4_c_21_n N_4_c_22_n N_4_c_23_n N_4_c_24_n N_4_c_45_p
+ N_4_c_25_n N_4_c_26_n N_4_c_27_n N_4_c_28_n N_4_c_34_p N_4_c_29_n N_4_c_30_n
+ N_4_c_31_n N_4_c_40_p N_4_c_48_p N_4_c_32_n VSS PM_BUFX5_ASAP7_75T_SRAM%4
x_PM_BUFX5_ASAP7_75T_SRAM%Y N_Y_M2_d N_Y_M1_d N_Y_M4_d N_Y_M3_d N_Y_M5_d N_Y_M8_d
+ N_Y_M7_d N_Y_c_49_n N_Y_M10_d N_Y_M9_d N_Y_M11_d N_Y_c_50_n N_Y_c_51_n
+ N_Y_c_57_n Y N_Y_c_63_n VSS PM_BUFX5_ASAP7_75T_SRAM%Y
cc_1 N_A_M0_g N_4_M1_g 0.00287079f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_4_c_18_n 9.64278e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A_M0_g N_4_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_4 A N_4_c_20_n 0.00198071f $X=0.061 $Y=0.1365 $X2=0.056 $Y2=0.2025
cc_5 A N_4_c_21_n 6.00641e-19 $X=0.061 $Y=0.1365 $X2=0.054 $Y2=0.036
cc_6 A N_4_c_22_n 0.00198071f $X=0.061 $Y=0.1365 $X2=0.054 $Y2=0.036
cc_7 N_A_c_2_p N_4_c_23_n 2.65563e-19 $X=0.081 $Y=0.135 $X2=0.073 $Y2=0.036
cc_8 N_A_M0_g N_4_c_24_n 3.10016e-19 $X=0.081 $Y=0.0675 $X2=0.0875 $Y2=0.036
cc_9 A N_4_c_25_n 6.00641e-19 $X=0.061 $Y=0.1365 $X2=0.054 $Y2=0.234
cc_10 N_A_c_2_p N_4_c_26_n 2.65563e-19 $X=0.081 $Y=0.135 $X2=0.073 $Y2=0.234
cc_11 N_A_M0_g N_4_c_27_n 3.10016e-19 $X=0.081 $Y=0.0675 $X2=0.0875 $Y2=0.234
cc_12 A N_4_c_28_n 7.49723e-19 $X=0.061 $Y=0.1365 $X2=0.111 $Y2=0.126
cc_13 A N_4_c_29_n 3.37664e-19 $X=0.061 $Y=0.1365 $X2=0.111 $Y2=0.081
cc_14 A N_4_c_30_n 7.49723e-19 $X=0.061 $Y=0.1365 $X2=0.111 $Y2=0.189
cc_15 A N_4_c_31_n 3.37664e-19 $X=0.061 $Y=0.1365 $X2=0.111 $Y2=0.207
cc_16 A N_4_c_32_n 0.00104772f $X=0.061 $Y=0.1365 $X2=0.111 $Y2=0.135
cc_17 N_4_c_30_n N_Y_c_49_n 0.00112297f $X=0.111 $Y=0.189 $X2=0 $Y2=0
cc_18 N_4_c_34_p N_Y_c_50_n 0.00112297f $X=0.111 $Y=0.063 $X2=0 $Y2=0
cc_19 N_4_M2_g N_Y_c_51_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_20 N_4_M3_g N_Y_c_51_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_21 N_4_M4_g N_Y_c_51_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_22 N_4_M5_g N_Y_c_51_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_23 N_4_c_39_p N_Y_c_51_n 0.00117364f $X=0.102 $Y=0.036 $X2=0 $Y2=0
cc_24 N_4_c_40_p N_Y_c_51_n 0.00408661f $X=0.167 $Y=0.135 $X2=0 $Y2=0
cc_25 N_4_M2_g N_Y_c_57_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_4_M3_g N_Y_c_57_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_4_M4_g N_Y_c_57_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_28 N_4_M5_g N_Y_c_57_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_29 N_4_c_45_p N_Y_c_57_n 0.00117364f $X=0.102 $Y=0.234 $X2=0 $Y2=0
cc_30 N_4_c_40_p N_Y_c_57_n 0.00408661f $X=0.167 $Y=0.135 $X2=0 $Y2=0
cc_31 N_4_c_47_p N_Y_c_63_n 3.12222e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_32 N_4_c_48_p N_Y_c_63_n 0.00114293f $X=0.351 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx5_ASAP7_75t_SRAM.pex.sp.BUFX5_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx6f_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:21:31 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx6f_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx6f_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx6f_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:21:31 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX6F_ASAP7_75T_SRAM%A 2 7 10 13 15 26 28 VSS
c19 28 VSS 0.0031408f $X=0.07 $Y=0.135
c20 26 VSS 0.013878f $X=0.053 $Y=0.136
c21 13 VSS 0.00719316f $X=0.135 $Y=0.1345
c22 10 VSS 0.0611108f $X=0.135 $Y=0.0675
c23 2 VSS 0.0653556f $X=0.081 $Y=0.0675
r24 28 29 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.07 $Y=0.135 $X2=0.07
+ $Y2=0.135
r25 26 28 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.053
+ $Y=0.135 $X2=0.07 $Y2=0.135
r26 13 15 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1345 $X2=0.135 $Y2=0.2025
r27 10 13 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1345
r28 5 13 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1345 $X2=0.135 $Y2=0.1345
r29 5 29 9.56522 $w=2.3e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1345 $X2=0.07 $Y2=0.1345
r30 5 7 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1345 $X2=0.081 $Y2=0.2025
r31 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.1345
.ends

.subckt PM_BUFX6F_ASAP7_75T_SRAM%4 2 7 10 15 18 23 26 31 34 39 42 45 47 49 50 54 55
+ 58 60 62 67 68 70 75 77 78 85 86 89 VSS
c43 86 VSS 0.00402867f $X=0.126 $Y=0.234
c44 85 VSS 0.00264717f $X=0.135 $Y=0.234
c45 78 VSS 0.00402695f $X=0.126 $Y=0.036
c46 77 VSS 0.00264717f $X=0.135 $Y=0.036
c47 75 VSS 0.0106764f $X=0.108 $Y=0.036
c48 70 VSS 2.71675e-19 $X=0.405 $Y=0.135
c49 67 VSS 0.00280848f $X=0.202 $Y=0.135
c50 62 VSS 0.00385172f $X=0.135 $Y=0.225
c51 60 VSS 0.00382416f $X=0.135 $Y=0.126
c52 58 VSS 0.0106764f $X=0.108 $Y=0.2025
c53 54 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c54 49 VSS 5.72268e-19 $X=0.125 $Y=0.0675
c55 45 VSS 0.0191506f $X=0.459 $Y=0.135
c56 42 VSS 0.0645347f $X=0.459 $Y=0.0675
c57 34 VSS 0.0644226f $X=0.405 $Y=0.0675
c58 26 VSS 0.0642127f $X=0.351 $Y=0.0675
c59 18 VSS 0.0642127f $X=0.297 $Y=0.0675
c60 10 VSS 0.0642127f $X=0.243 $Y=0.0675
c61 2 VSS 0.0616955f $X=0.189 $Y=0.0675
r62 86 87 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r63 85 87 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r64 82 86 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r65 78 79 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r66 77 79 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r67 74 78 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r68 74 75 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r69 67 68 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.135 $X2=0.2225 $Y2=0.135
r70 65 70 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.405 $Y2=0.135
r71 65 68 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.2225 $Y2=0.135
r72 63 89 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.135 $Y2=0.135
r73 63 67 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.202 $Y2=0.135
r74 62 85 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.234
r75 61 89 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.135
r76 61 62 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.225
r77 60 89 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.135
r78 59 77 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.036
r79 59 60 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.126
r80 58 82 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r81 55 58 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r82 54 58 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r83 53 75 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r84 50 53 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r85 49 53 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r86 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r87 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r88 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r89 37 70 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r90 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r91 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
r92 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r93 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r94 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r95 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r96 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r97 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r98 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r99 13 65 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r100 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.2025
r101 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.135
r102 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r103 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r104 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_BUFX6F_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 21 22 26 27 42 55 60 62 VSS
c24 62 VSS 7.46921e-19 $X=0.513 $Y=0.144
c25 61 VSS 0.00538124f $X=0.513 $Y=0.126
c26 60 VSS 0.00538124f $X=0.514 $Y=0.153
c27 56 VSS 0.00294383f $X=0.4885 $Y=0.234
c28 55 VSS 0.0284173f $X=0.473 $Y=0.234
c29 44 VSS 0.005853f $X=0.504 $Y=0.234
c30 43 VSS 0.00294383f $X=0.4885 $Y=0.036
c31 42 VSS 0.0284173f $X=0.473 $Y=0.036
c32 41 VSS 0.00929752f $X=0.432 $Y=0.036
c33 38 VSS 0.00928955f $X=0.324 $Y=0.036
c34 34 VSS 0.00916652f $X=0.216 $Y=0.036
c35 31 VSS 0.005853f $X=0.504 $Y=0.036
c36 30 VSS 0.00929752f $X=0.432 $Y=0.2025
c37 26 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c38 25 VSS 0.00928955f $X=0.324 $Y=0.2025
c39 21 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c40 20 VSS 0.00916652f $X=0.216 $Y=0.2025
c41 16 VSS 5.72268e-19 $X=0.233 $Y=0.2025
c42 11 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c43 6 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c44 1 VSS 5.72268e-19 $X=0.233 $Y=0.0675
r45 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.126 $X2=0.513 $Y2=0.144
r46 60 62 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.153 $X2=0.513 $Y2=0.144
r47 58 60 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.153
r48 57 61 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.126
r49 55 56 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.473
+ $Y=0.234 $X2=0.4885 $Y2=0.234
r50 53 55 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.473 $Y2=0.234
r51 50 53 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r52 46 50 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.324 $Y2=0.234
r53 44 58 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.234 $X2=0.513 $Y2=0.225
r54 44 56 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.4885 $Y2=0.234
r55 42 43 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.473
+ $Y=0.036 $X2=0.4885 $Y2=0.036
r56 40 42 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.473 $Y2=0.036
r57 40 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r58 37 40 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r59 37 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r60 33 37 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.324 $Y2=0.036
r61 33 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r62 31 57 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.036 $X2=0.513 $Y2=0.045
r63 31 43 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.4885 $Y2=0.036
r64 30 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r65 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r66 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r67 25 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r68 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r69 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r70 20 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r71 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r72 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r73 15 41 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r74 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r75 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r76 10 38 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r77 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r78 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r79 5 34 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r80 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r81 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./BUFx6f_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx6f_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_4_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_4_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_4_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_4_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_4_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_4_M6_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_4_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_4_M8_d N_A_M8_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M9 N_4_M9_d N_A_M9_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M10 N_Y_M10_d N_4_M10_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M11 N_Y_M11_d N_4_M11_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M12 N_Y_M12_d N_4_M12_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M13 N_Y_M13_d N_4_M13_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M14 N_Y_M14_d N_4_M14_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M15 N_Y_M15_d N_4_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "BUFx6f_ASAP7_75t_SRAM.pex.sp.BUFX6F_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx6f_ASAP7_75t_SRAM.pex.sp.BUFX6F_ASAP7_75T_SRAM.pxi"
* File: BUFx6f_ASAP7_75t_SRAM.pex.sp.BUFX6F_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:21:31 2017
* 
x_PM_BUFX6F_ASAP7_75T_SRAM%A N_A_M0_g N_A_M8_g N_A_M1_g N_A_c_4_p N_A_M9_g A
+ N_A_c_19_p VSS PM_BUFX6F_ASAP7_75T_SRAM%A
x_PM_BUFX6F_ASAP7_75T_SRAM%4 N_4_M2_g N_4_M10_g N_4_M3_g N_4_M11_g N_4_M4_g
+ N_4_M12_g N_4_M5_g N_4_M13_g N_4_M6_g N_4_M14_g N_4_M7_g N_4_c_23_n N_4_M15_g
+ N_4_M1_d N_4_M0_d N_4_M9_d N_4_M8_d N_4_c_26_n N_4_c_27_n N_4_c_30_n
+ N_4_c_33_n N_4_c_51_p N_4_c_62_p N_4_c_34_n N_4_c_52_p N_4_c_35_n N_4_c_60_p
+ N_4_c_36_n N_4_c_37_n VSS PM_BUFX6F_ASAP7_75T_SRAM%4
x_PM_BUFX6F_ASAP7_75T_SRAM%Y N_Y_M3_d N_Y_M2_d N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M6_d
+ N_Y_M11_d N_Y_M10_d N_Y_M13_d N_Y_M12_d N_Y_M15_d N_Y_M14_d N_Y_c_69_n
+ N_Y_c_77_n Y N_Y_c_85_n VSS PM_BUFX6F_ASAP7_75T_SRAM%Y
cc_1 N_A_M0_g N_4_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_A_M1_g N_4_M2_g 0.00287079f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A_M1_g N_4_M3_g 2.34385e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_4 N_A_c_4_p N_4_c_23_n 0.00202955f $X=0.135 $Y=0.1345 $X2=0.459 $Y2=0.135
cc_5 N_A_c_4_p N_4_M1_d 3.89905e-19 $X=0.135 $Y=0.1345 $X2=0.125 $Y2=0.0675
cc_6 N_A_c_4_p N_4_M9_d 3.83499e-19 $X=0.135 $Y=0.1345 $X2=0.125 $Y2=0.2025
cc_7 N_A_c_4_p N_4_c_26_n 8.01479e-19 $X=0.135 $Y=0.1345 $X2=0.108 $Y2=0.2025
cc_8 N_A_M1_g N_4_c_27_n 6.21137e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.126
cc_9 N_A_c_4_p N_4_c_27_n 5.0686e-19 $X=0.135 $Y=0.1345 $X2=0.135 $Y2=0.126
cc_10 A N_4_c_27_n 6.86581e-19 $X=0.053 $Y=0.136 $X2=0.135 $Y2=0.126
cc_11 N_A_M1_g N_4_c_30_n 6.45702e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.225
cc_12 N_A_c_4_p N_4_c_30_n 4.76028e-19 $X=0.135 $Y=0.1345 $X2=0.135 $Y2=0.225
cc_13 A N_4_c_30_n 6.94667e-19 $X=0.053 $Y=0.136 $X2=0.135 $Y2=0.225
cc_14 N_A_c_4_p N_4_c_33_n 4.3862e-19 $X=0.135 $Y=0.1345 $X2=0.202 $Y2=0.135
cc_15 N_A_c_4_p N_4_c_34_n 8.45347e-19 $X=0.135 $Y=0.1345 $X2=0.108 $Y2=0.036
cc_16 N_A_c_4_p N_4_c_35_n 3.42736e-19 $X=0.135 $Y=0.1345 $X2=0.126 $Y2=0.036
cc_17 N_A_c_4_p N_4_c_36_n 3.39414e-19 $X=0.135 $Y=0.1345 $X2=0.126 $Y2=0.234
cc_18 N_A_c_4_p N_4_c_37_n 0.00112176f $X=0.135 $Y=0.1345 $X2=0.135 $Y2=0.135
cc_19 N_A_c_19_p N_4_c_37_n 6.83331e-19 $X=0.07 $Y=0.135 $X2=0.135 $Y2=0.135
cc_20 N_4_c_23_n N_Y_M3_d 3.80218e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_21 N_4_c_23_n N_Y_M5_d 3.80218e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_22 N_4_c_23_n N_Y_M7_d 3.80218e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_23 N_4_c_23_n N_Y_M11_d 3.80218e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_24 N_4_c_23_n N_Y_M13_d 3.80218e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_25 N_4_c_23_n N_Y_M15_d 3.80218e-19 $X=0.459 $Y=0.135 $X2=0.053 $Y2=0.136
cc_26 N_4_M3_g N_Y_c_69_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_4_M4_g N_Y_c_69_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_28 N_4_M5_g N_Y_c_69_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_29 N_4_M6_g N_Y_c_69_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_4_M7_g N_Y_c_69_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_4_c_23_n N_Y_c_69_n 9.87293e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_32 N_4_c_51_p N_Y_c_69_n 0.00367654f $X=0.2225 $Y=0.135 $X2=0 $Y2=0
cc_33 N_4_c_52_p N_Y_c_69_n 3.81483e-19 $X=0.135 $Y=0.036 $X2=0 $Y2=0
cc_34 N_4_M3_g N_Y_c_77_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_4_M4_g N_Y_c_77_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_4_M5_g N_Y_c_77_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_4_M6_g N_Y_c_77_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_38 N_4_M7_g N_Y_c_77_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_4_c_23_n N_Y_c_77_n 9.87293e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_40 N_4_c_51_p N_Y_c_77_n 0.00367654f $X=0.2225 $Y=0.135 $X2=0 $Y2=0
cc_41 N_4_c_60_p N_Y_c_77_n 3.81483e-19 $X=0.135 $Y=0.234 $X2=0 $Y2=0
cc_42 N_4_c_23_n N_Y_c_85_n 4.79181e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_43 N_4_c_62_p N_Y_c_85_n 0.0010395f $X=0.405 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx6f_ASAP7_75t_SRAM.pex.sp.BUFX6F_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: BUFx8_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:21:54 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "BUFx8_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./BUFx8_ASAP7_75t_SRAM.pex.sp.pex"
* File: BUFx8_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:21:54 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_BUFX8_ASAP7_75T_SRAM%A 2 7 10 13 15 23 27 VSS
c19 27 VSS 0.00106669f $X=0.081 $Y=0.135
c20 23 VSS 0.0249674f $X=0.0715 $Y=0.134
c21 13 VSS 0.00763526f $X=0.135 $Y=0.135
c22 10 VSS 0.0582189f $X=0.135 $Y=0.054
c23 2 VSS 0.0624608f $X=0.081 $Y=0.054
r24 23 27 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.0715
+ $Y=0.135 $X2=0.081 $Y2=0.135
r25 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r26 10 13 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
r27 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r28 5 27 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r29 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r30 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_BUFX8_ASAP7_75T_SRAM%4 2 7 10 15 18 23 26 31 34 39 42 47 50 55 58 61 63
+ 65 66 69 70 71 74 76 78 83 84 89 93 98 103 108 112 VSS
c49 109 VSS 0.00202053f $X=0.126 $Y=0.234
c50 108 VSS 0.00264832f $X=0.135 $Y=0.234
c51 103 VSS 0.00209506f $X=0.108 $Y=0.234
c52 99 VSS 0.00202053f $X=0.126 $Y=0.036
c53 98 VSS 0.00264832f $X=0.135 $Y=0.036
c54 93 VSS 0.00209506f $X=0.108 $Y=0.036
c55 83 VSS 0.00279153f $X=0.202 $Y=0.135
c56 78 VSS 0.00351237f $X=0.135 $Y=0.225
c57 76 VSS 0.00351237f $X=0.135 $Y=0.126
c58 74 VSS 0.008461f $X=0.108 $Y=0.216
c59 70 VSS 5.3314e-19 $X=0.125 $Y=0.216
c60 69 VSS 0.008461f $X=0.108 $Y=0.054
c61 65 VSS 5.3314e-19 $X=0.125 $Y=0.054
c62 61 VSS 0.0256482f $X=0.567 $Y=0.135
c63 58 VSS 0.0615048f $X=0.567 $Y=0.0675
c64 50 VSS 0.061544f $X=0.513 $Y=0.0675
c65 42 VSS 0.0613551f $X=0.459 $Y=0.0675
c66 34 VSS 0.0613551f $X=0.405 $Y=0.0675
c67 26 VSS 0.0613551f $X=0.351 $Y=0.0675
c68 18 VSS 0.0613551f $X=0.297 $Y=0.0675
c69 10 VSS 0.0613551f $X=0.243 $Y=0.0675
c70 2 VSS 0.0588727f $X=0.189 $Y=0.0675
r71 109 110 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r72 108 110 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r73 103 109 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r74 99 100 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r75 98 100 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r76 93 99 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r77 86 89 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.513 $Y2=0.135
r78 83 84 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.135 $X2=0.2225 $Y2=0.135
r79 81 86 11 $w=1.8e-08 $l=1.62e-07 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.405 $Y2=0.135
r80 81 84 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.2225 $Y2=0.135
r81 79 112 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.135 $Y2=0.135
r82 79 83 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.202 $Y2=0.135
r83 78 108 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.234
r84 77 112 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.135
r85 77 78 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.225
r86 76 112 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.135
r87 75 98 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.036
r88 75 76 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.126
r89 74 103 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r90 71 74 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.216 $X2=0.108 $Y2=0.216
r91 70 74 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.216 $X2=0.108 $Y2=0.216
r92 69 93 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r93 66 69 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.054 $X2=0.108 $Y2=0.054
r94 65 69 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.054 $X2=0.108 $Y2=0.054
r95 61 63 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r96 58 61 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r97 53 61 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r98 53 89 3.03549 $a=6.48e-16 $layer=V0LIG $count=2 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r99 53 55 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r100 50 53 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r101 45 53 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r102 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r103 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r104 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r105 37 86 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r106 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r107 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r108 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r109 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r110 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r111 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r112 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.135 $X2=0.297 $Y2=0.2025
r113 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.0675 $X2=0.297 $Y2=0.135
r114 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r115 13 81 2.02366 $a=9.72e-16 $layer=V0LIG $count=3 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r116 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.2025
r117 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.135
r118 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r119 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r120 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_BUFX8_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 21 22 26 27 31 32 36 37 55 71
+ 76 78 VSS
c30 78 VSS 7.61289e-19 $X=0.621 $Y=0.144
c31 76 VSS 0.00529396f $X=0.6215 $Y=0.113
c32 74 VSS 0.00529396f $X=0.621 $Y=0.225
c33 72 VSS 0.00294383f $X=0.5965 $Y=0.234
c34 71 VSS 0.0399184f $X=0.581 $Y=0.234
c35 57 VSS 0.00586994f $X=0.612 $Y=0.234
c36 56 VSS 0.00294383f $X=0.5965 $Y=0.036
c37 55 VSS 0.0399184f $X=0.581 $Y=0.036
c38 54 VSS 0.00929752f $X=0.54 $Y=0.036
c39 51 VSS 0.00928955f $X=0.432 $Y=0.036
c40 48 VSS 0.00928955f $X=0.324 $Y=0.036
c41 44 VSS 0.00911786f $X=0.216 $Y=0.036
c42 41 VSS 0.00586994f $X=0.612 $Y=0.036
c43 40 VSS 0.00929752f $X=0.54 $Y=0.2025
c44 36 VSS 5.38922e-19 $X=0.557 $Y=0.2025
c45 35 VSS 0.00928955f $X=0.432 $Y=0.2025
c46 31 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c47 30 VSS 0.00928955f $X=0.324 $Y=0.2025
c48 26 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c49 25 VSS 0.00911786f $X=0.216 $Y=0.2025
c50 21 VSS 5.72268e-19 $X=0.233 $Y=0.2025
c51 16 VSS 5.38922e-19 $X=0.557 $Y=0.0675
c52 11 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c53 6 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c54 1 VSS 5.72268e-19 $X=0.233 $Y=0.0675
r55 77 78 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.126 $X2=0.621 $Y2=0.144
r56 76 77 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.113 $X2=0.621 $Y2=0.126
r57 74 78 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.144
r58 73 76 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.113
r59 71 72 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.581
+ $Y=0.234 $X2=0.5965 $Y2=0.234
r60 69 71 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.581 $Y2=0.234
r61 66 69 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.54 $Y2=0.234
r62 63 66 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r63 59 63 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.324 $Y2=0.234
r64 57 74 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r65 57 72 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.5965 $Y2=0.234
r66 55 56 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.581
+ $Y=0.036 $X2=0.5965 $Y2=0.036
r67 53 55 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.581 $Y2=0.036
r68 53 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r69 50 53 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.54 $Y2=0.036
r70 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r71 47 50 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r72 47 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r73 43 47 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.324 $Y2=0.036
r74 43 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r75 41 73 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r76 41 56 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.5965 $Y2=0.036
r77 40 69 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r78 37 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r79 36 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r80 35 66 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r81 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r82 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r83 30 63 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r84 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r85 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r86 25 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r87 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r88 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r89 20 54 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r90 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r91 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r92 15 51 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r93 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r94 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r95 10 48 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r96 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r97 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r98 5 44 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r99 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r100 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./BUFx8_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt BUFx8_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_4_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_4_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_4_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_4_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_4_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_4_M6_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_4_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_4_M8_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_4_M9_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 N_4_M10_d N_A_M10_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M11 N_4_M11_d N_A_M11_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M12 N_Y_M12_d N_4_M12_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M13 N_Y_M13_d N_4_M13_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M14 N_Y_M14_d N_4_M14_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M15 N_Y_M15_d N_4_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M16 N_Y_M16_d N_4_M16_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M17 N_Y_M17_d N_4_M17_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M18 N_Y_M18_d N_4_M18_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M19 N_Y_M19_d N_4_M19_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
*
* 
* .include "BUFx8_ASAP7_75t_SRAM.pex.sp.BUFX8_ASAP7_75T_SRAM.pxi"
* BEGIN of "./BUFx8_ASAP7_75t_SRAM.pex.sp.BUFX8_ASAP7_75T_SRAM.pxi"
* File: BUFx8_ASAP7_75t_SRAM.pex.sp.BUFX8_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:21:54 2017
* 
x_PM_BUFX8_ASAP7_75T_SRAM%A N_A_M0_g N_A_M10_g N_A_M1_g N_A_c_4_p N_A_M11_g A
+ N_A_c_19_p VSS PM_BUFX8_ASAP7_75T_SRAM%A
x_PM_BUFX8_ASAP7_75T_SRAM%4 N_4_M2_g N_4_M12_g N_4_M3_g N_4_M13_g N_4_M4_g
+ N_4_M14_g N_4_M5_g N_4_M15_g N_4_M6_g N_4_M16_g N_4_M7_g N_4_M17_g N_4_M8_g
+ N_4_M18_g N_4_M9_g N_4_c_23_n N_4_M19_g N_4_M1_d N_4_M0_d N_4_c_24_n N_4_M11_d
+ N_4_M10_d N_4_c_25_n N_4_c_26_n N_4_c_29_n N_4_c_32_n N_4_c_55_p N_4_c_68_p
+ N_4_c_33_n N_4_c_56_p N_4_c_35_n N_4_c_66_p N_4_c_37_n VSS
+ PM_BUFX8_ASAP7_75T_SRAM%4
x_PM_BUFX8_ASAP7_75T_SRAM%Y N_Y_M3_d N_Y_M2_d N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M6_d
+ N_Y_M9_d N_Y_M8_d N_Y_M13_d N_Y_M12_d N_Y_M15_d N_Y_M14_d N_Y_M17_d N_Y_M16_d
+ N_Y_M19_d N_Y_M18_d N_Y_c_77_n N_Y_c_87_n Y N_Y_c_98_n VSS
+ PM_BUFX8_ASAP7_75T_SRAM%Y
cc_1 N_A_M0_g N_4_M2_g 2.13359e-19 $X=0.081 $Y=0.054 $X2=0.189 $Y2=0.0675
cc_2 N_A_M1_g N_4_M2_g 0.00268443f $X=0.135 $Y=0.054 $X2=0.189 $Y2=0.0675
cc_3 N_A_M1_g N_4_M3_g 2.13359e-19 $X=0.135 $Y=0.054 $X2=0.243 $Y2=0.0675
cc_4 N_A_c_4_p N_4_c_23_n 0.00154814f $X=0.135 $Y=0.135 $X2=0.567 $Y2=0.135
cc_5 N_A_c_4_p N_4_c_24_n 3.91995e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.054
cc_6 N_A_c_4_p N_4_c_25_n 3.91995e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.216
cc_7 N_A_M1_g N_4_c_26_n 7.69468e-19 $X=0.135 $Y=0.054 $X2=0.135 $Y2=0.126
cc_8 N_A_c_4_p N_4_c_26_n 4.76064e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.126
cc_9 A N_4_c_26_n 0.0010108f $X=0.0715 $Y=0.134 $X2=0.135 $Y2=0.126
cc_10 N_A_M1_g N_4_c_29_n 7.69468e-19 $X=0.135 $Y=0.054 $X2=0.135 $Y2=0.225
cc_11 N_A_c_4_p N_4_c_29_n 4.76064e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.225
cc_12 A N_4_c_29_n 0.0010108f $X=0.0715 $Y=0.134 $X2=0.135 $Y2=0.225
cc_13 N_A_c_4_p N_4_c_32_n 5.49367e-19 $X=0.135 $Y=0.135 $X2=0.202 $Y2=0.135
cc_14 N_A_c_4_p N_4_c_33_n 3.3231e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.036
cc_15 A N_4_c_33_n 5.37037e-19 $X=0.0715 $Y=0.134 $X2=0.108 $Y2=0.036
cc_16 N_A_c_4_p N_4_c_35_n 3.3231e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.234
cc_17 A N_4_c_35_n 5.37037e-19 $X=0.0715 $Y=0.134 $X2=0.108 $Y2=0.234
cc_18 N_A_c_4_p N_4_c_37_n 0.00102271f $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.135
cc_19 N_A_c_19_p N_4_c_37_n 0.00105996f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_20 N_4_c_23_n N_Y_M3_d 3.80218e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.054
cc_21 N_4_c_23_n N_Y_M5_d 3.80218e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.216
cc_22 N_4_c_23_n N_Y_M7_d 3.80218e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_23 N_4_c_23_n N_Y_M9_d 3.80218e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_24 N_4_c_23_n N_Y_M13_d 3.80218e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_25 N_4_c_23_n N_Y_M15_d 3.80218e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.135
cc_26 N_4_c_23_n N_Y_M17_d 3.80218e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_27 N_4_c_23_n N_Y_M19_d 3.80218e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.135
cc_28 N_4_M3_g N_Y_c_77_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_29 N_4_M4_g N_Y_c_77_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_4_M5_g N_Y_c_77_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_31 N_4_M6_g N_Y_c_77_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_32 N_4_M7_g N_Y_c_77_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_33 N_4_M8_g N_Y_c_77_n 4.28653e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_34 N_4_M9_g N_Y_c_77_n 4.28653e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_4_c_23_n N_Y_c_77_n 0.00140144f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_36 N_4_c_55_p N_Y_c_77_n 0.00512201f $X=0.2225 $Y=0.135 $X2=0 $Y2=0
cc_37 N_4_c_56_p N_Y_c_77_n 3.8417e-19 $X=0.135 $Y=0.036 $X2=0 $Y2=0
cc_38 N_4_M3_g N_Y_c_87_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_4_M4_g N_Y_c_87_n 4.28653e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_40 N_4_M5_g N_Y_c_87_n 4.28653e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_41 N_4_M6_g N_Y_c_87_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_42 N_4_M7_g N_Y_c_87_n 4.28653e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_4_M8_g N_Y_c_87_n 4.28653e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_4_M9_g N_Y_c_87_n 4.28653e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_45 N_4_c_23_n N_Y_c_87_n 0.00140144f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_46 N_4_c_55_p N_Y_c_87_n 0.00512201f $X=0.2225 $Y=0.135 $X2=0 $Y2=0
cc_47 N_4_c_66_p N_Y_c_87_n 3.8417e-19 $X=0.135 $Y=0.234 $X2=0 $Y2=0
cc_48 N_4_c_23_n Y 4.27377e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_49 N_4_c_68_p N_Y_c_98_n 8.73292e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0

* END of "./BUFx8_ASAP7_75t_SRAM.pex.sp.BUFX8_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVx11_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:32:45 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVx11_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVx11_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVx11_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:32:45 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVX11_ASAP7_75T_SRAM%A 2 7 10 15 18 23 26 31 34 39 42 47 50 55 58 63 66
+ 71 74 79 82 85 87 95 VSS
c45 95 VSS 0.0275187f $X=0.063 $Y=0.1355
c46 85 VSS 0.0581303f $X=0.621 $Y=0.135
c47 82 VSS 0.0678263f $X=0.621 $Y=0.0675
c48 74 VSS 0.0643964f $X=0.567 $Y=0.0675
c49 66 VSS 0.0642127f $X=0.513 $Y=0.0675
c50 58 VSS 0.0642127f $X=0.459 $Y=0.0675
c51 50 VSS 0.0642127f $X=0.405 $Y=0.0675
c52 42 VSS 0.0642127f $X=0.351 $Y=0.0675
c53 34 VSS 0.0642127f $X=0.297 $Y=0.0675
c54 26 VSS 0.0642127f $X=0.243 $Y=0.0675
c55 18 VSS 0.0642127f $X=0.189 $Y=0.0675
c56 10 VSS 0.0644226f $X=0.135 $Y=0.0675
c57 2 VSS 0.0655089f $X=0.081 $Y=0.0675
r58 95 99 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r59 85 87 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r60 82 85 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
r61 77 85 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.567
+ $Y=0.135 $X2=0.621 $Y2=0.135
r62 77 79 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r63 74 77 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r64 69 77 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r65 69 71 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r66 66 69 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
r67 61 69 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r68 61 63 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r69 58 61 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r70 53 61 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r71 53 55 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r72 50 53 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
r73 45 53 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r74 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r75 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r76 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r77 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r78 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r79 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r80 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r81 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r82 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r83 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r84 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r85 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r86 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r87 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r88 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r89 5 99 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r90 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r91 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVX11_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 21 22 26 31 32 35 36 37 40
+ 41 42 45 46 47 50 51 52 55 56 61 64 68 71 74 77 81 104 VSS
c45 104 VSS 0.00874911f $X=0.6775 $Y=0.1475
c46 81 VSS 0.0676509f $X=0.666 $Y=0.234
c47 80 VSS 0.00692279f $X=0.648 $Y=0.036
c48 77 VSS 0.00928905f $X=0.54 $Y=0.036
c49 74 VSS 0.00928955f $X=0.432 $Y=0.036
c50 71 VSS 0.00928955f $X=0.324 $Y=0.036
c51 68 VSS 0.00928954f $X=0.216 $Y=0.036
c52 64 VSS 0.00904082f $X=0.108 $Y=0.036
c53 61 VSS 0.0676509f $X=0.666 $Y=0.036
c54 59 VSS 0.00726838f $X=0.646 $Y=0.2025
c55 55 VSS 0.00928905f $X=0.54 $Y=0.2025
c56 51 VSS 5.38922e-19 $X=0.557 $Y=0.2025
c57 50 VSS 0.00928955f $X=0.432 $Y=0.2025
c58 46 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c59 45 VSS 0.00928955f $X=0.324 $Y=0.2025
c60 41 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c61 40 VSS 0.00928954f $X=0.216 $Y=0.2025
c62 36 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c63 35 VSS 0.00904082f $X=0.108 $Y=0.2025
c64 31 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c65 29 VSS 3.45593e-19 $X=0.646 $Y=0.0675
c66 21 VSS 5.38922e-19 $X=0.557 $Y=0.0675
c67 16 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c68 11 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c69 6 VSS 5.38922e-19 $X=0.233 $Y=0.0675
c70 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r71 102 104 5.26235 $w=1.8e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.675
+ $Y=0.225 $X2=0.675 $Y2=0.1475
r72 101 104 6.95988 $w=1.8e-08 $l=1.025e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.675 $Y=0.045 $X2=0.675 $Y2=0.1475
r73 96 99 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.648 $Y2=0.234
r74 93 96 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.54 $Y2=0.234
r75 90 93 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r76 87 90 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.324 $Y2=0.234
r77 83 87 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.216 $Y2=0.234
r78 81 102 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.234 $X2=0.675 $Y2=0.225
r79 81 99 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.234 $X2=0.648 $Y2=0.234
r80 79 80 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036 $X2=0.648
+ $Y2=0.036
r81 76 79 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.648 $Y2=0.036
r82 76 77 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r83 73 76 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.54 $Y2=0.036
r84 73 74 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r85 70 73 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r86 70 71 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r87 67 70 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.324 $Y2=0.036
r88 67 68 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r89 63 67 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.216 $Y2=0.036
r90 63 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r91 61 101 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.666 $Y=0.036 $X2=0.675 $Y2=0.045
r92 61 79 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.036 $X2=0.648 $Y2=0.036
r93 59 99 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234 $X2=0.648
+ $Y2=0.234
r94 56 59 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.646 $Y2=0.2025
r95 55 96 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r96 52 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r97 51 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r98 50 93 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r99 47 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r100 46 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r101 45 90 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r102 42 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r103 41 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r104 40 87 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r105 37 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r106 36 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r107 35 83 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r108 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r109 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r110 29 80 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r111 26 29 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.646 $Y2=0.0675
r112 25 77 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r113 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r114 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r115 20 74 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r116 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r117 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r118 15 71 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r119 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r120 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r121 10 68 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.216 $Y=0.0675 $X2=0.216 $Y2=0.036
r122 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r123 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r124 5 64 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r125 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r126 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./INVx11_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVx11_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_A_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_A_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_A_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_A_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_A_M6_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_A_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_A_M8_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_A_M9_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 N_Y_M10_d N_A_M10_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M11 N_Y_M11_d N_A_M11_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M12 N_Y_M12_d N_A_M12_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M13 N_Y_M13_d N_A_M13_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M14 N_Y_M14_d N_A_M14_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M15 N_Y_M15_d N_A_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M16 N_Y_M16_d N_A_M16_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M17 N_Y_M17_d N_A_M17_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M18 N_Y_M18_d N_A_M18_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M19 N_Y_M19_d N_A_M19_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M20 N_Y_M20_d N_A_M20_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M21 N_Y_M21_d N_A_M21_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
*
* 
* .include "INVx11_ASAP7_75t_SRAM.pex.sp.INVX11_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVx11_ASAP7_75t_SRAM.pex.sp.INVX11_ASAP7_75T_SRAM.pxi"
* File: INVx11_ASAP7_75t_SRAM.pex.sp.INVX11_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:32:45 2017
* 
x_PM_INVX11_ASAP7_75T_SRAM%A N_A_M0_g N_A_M11_g N_A_M1_g N_A_M12_g N_A_M2_g
+ N_A_M13_g N_A_M3_g N_A_M14_g N_A_M4_g N_A_M15_g N_A_M5_g N_A_M16_g N_A_M6_g
+ N_A_M17_g N_A_M7_g N_A_M18_g N_A_M8_g N_A_M19_g N_A_M9_g N_A_M20_g N_A_M10_g
+ N_A_c_1_p N_A_M21_g A VSS PM_INVX11_ASAP7_75T_SRAM%A
x_PM_INVX11_ASAP7_75T_SRAM%Y N_Y_M1_d N_Y_M0_d N_Y_M3_d N_Y_M2_d N_Y_M5_d N_Y_M4_d
+ N_Y_M7_d N_Y_M6_d N_Y_M9_d N_Y_M8_d N_Y_M10_d N_Y_M12_d N_Y_M11_d N_Y_c_52_n
+ N_Y_M14_d N_Y_M13_d N_Y_c_54_n N_Y_M16_d N_Y_M15_d N_Y_c_56_n N_Y_M18_d
+ N_Y_M17_d N_Y_c_58_n N_Y_M20_d N_Y_M19_d N_Y_c_60_n N_Y_M21_d N_Y_c_61_n
+ N_Y_c_73_n N_Y_c_74_n N_Y_c_75_n N_Y_c_76_n N_Y_c_77_n N_Y_c_78_n Y VSS
+ PM_INVX11_ASAP7_75T_SRAM%Y
cc_1 N_A_c_1_p N_Y_M1_d 3.80663e-19 $X=0.621 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_2 N_A_c_1_p N_Y_M3_d 3.80663e-19 $X=0.621 $Y=0.135 $X2=0.233 $Y2=0.0675
cc_3 N_A_c_1_p N_Y_M5_d 3.80663e-19 $X=0.621 $Y=0.135 $X2=0.341 $Y2=0.0675
cc_4 N_A_c_1_p N_Y_M7_d 3.80663e-19 $X=0.621 $Y=0.135 $X2=0.449 $Y2=0.0675
cc_5 N_A_c_1_p N_Y_M9_d 3.80663e-19 $X=0.621 $Y=0.135 $X2=0.557 $Y2=0.0675
cc_6 N_A_c_1_p N_Y_M12_d 3.80663e-19 $X=0.621 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_7 N_A_c_1_p N_Y_c_52_n 8.00061e-19 $X=0.621 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_8 N_A_c_1_p N_Y_M14_d 3.80663e-19 $X=0.621 $Y=0.135 $X2=0.233 $Y2=0.2025
cc_9 N_A_c_1_p N_Y_c_54_n 8.00061e-19 $X=0.621 $Y=0.135 $X2=0.216 $Y2=0.2025
cc_10 N_A_c_1_p N_Y_M16_d 3.80663e-19 $X=0.621 $Y=0.135 $X2=0.341 $Y2=0.2025
cc_11 N_A_c_1_p N_Y_c_56_n 8.00061e-19 $X=0.621 $Y=0.135 $X2=0.324 $Y2=0.2025
cc_12 N_A_c_1_p N_Y_M18_d 3.80663e-19 $X=0.621 $Y=0.135 $X2=0.449 $Y2=0.2025
cc_13 N_A_c_1_p N_Y_c_58_n 8.00061e-19 $X=0.621 $Y=0.135 $X2=0.432 $Y2=0.2025
cc_14 N_A_c_1_p N_Y_M20_d 3.80663e-19 $X=0.621 $Y=0.135 $X2=0.557 $Y2=0.2025
cc_15 N_A_c_1_p N_Y_c_60_n 8.00061e-19 $X=0.621 $Y=0.135 $X2=0.54 $Y2=0.2025
cc_16 N_A_M1_g N_Y_c_61_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.666 $Y2=0.036
cc_17 N_A_M2_g N_Y_c_61_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.666 $Y2=0.036
cc_18 N_A_M3_g N_Y_c_61_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.666 $Y2=0.036
cc_19 N_A_M4_g N_Y_c_61_n 4.59284e-19 $X=0.297 $Y=0.0675 $X2=0.666 $Y2=0.036
cc_20 N_A_M5_g N_Y_c_61_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.666 $Y2=0.036
cc_21 N_A_M6_g N_Y_c_61_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0.666 $Y2=0.036
cc_22 N_A_M7_g N_Y_c_61_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.666 $Y2=0.036
cc_23 N_A_M8_g N_Y_c_61_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.666 $Y2=0.036
cc_24 N_A_M9_g N_Y_c_61_n 4.59284e-19 $X=0.567 $Y=0.0675 $X2=0.666 $Y2=0.036
cc_25 N_A_M10_g N_Y_c_61_n 4.59284e-19 $X=0.621 $Y=0.0675 $X2=0.666 $Y2=0.036
cc_26 N_A_c_1_p N_Y_c_61_n 0.00679508f $X=0.621 $Y=0.135 $X2=0.666 $Y2=0.036
cc_27 A N_Y_c_61_n 5.33309e-19 $X=0.063 $Y=0.1355 $X2=0.666 $Y2=0.036
cc_28 N_A_c_1_p N_Y_c_73_n 8.00061e-19 $X=0.621 $Y=0.135 $X2=0.108 $Y2=0.036
cc_29 N_A_c_1_p N_Y_c_74_n 8.00061e-19 $X=0.621 $Y=0.135 $X2=0.216 $Y2=0.036
cc_30 N_A_c_1_p N_Y_c_75_n 8.00061e-19 $X=0.621 $Y=0.135 $X2=0.324 $Y2=0.036
cc_31 N_A_c_1_p N_Y_c_76_n 8.00061e-19 $X=0.621 $Y=0.135 $X2=0.432 $Y2=0.036
cc_32 N_A_c_1_p N_Y_c_77_n 8.00061e-19 $X=0.621 $Y=0.135 $X2=0.54 $Y2=0.036
cc_33 N_A_M1_g N_Y_c_78_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.666 $Y2=0.234
cc_34 N_A_M2_g N_Y_c_78_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.666 $Y2=0.234
cc_35 N_A_M3_g N_Y_c_78_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.666 $Y2=0.234
cc_36 N_A_M4_g N_Y_c_78_n 4.59284e-19 $X=0.297 $Y=0.0675 $X2=0.666 $Y2=0.234
cc_37 N_A_M5_g N_Y_c_78_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.666 $Y2=0.234
cc_38 N_A_M6_g N_Y_c_78_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0.666 $Y2=0.234
cc_39 N_A_M7_g N_Y_c_78_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.666 $Y2=0.234
cc_40 N_A_M8_g N_Y_c_78_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.666 $Y2=0.234
cc_41 N_A_M9_g N_Y_c_78_n 4.59284e-19 $X=0.567 $Y=0.0675 $X2=0.666 $Y2=0.234
cc_42 N_A_M10_g N_Y_c_78_n 4.59284e-19 $X=0.621 $Y=0.0675 $X2=0.666 $Y2=0.234
cc_43 N_A_c_1_p N_Y_c_78_n 0.00679508f $X=0.621 $Y=0.135 $X2=0.666 $Y2=0.234
cc_44 A N_Y_c_78_n 5.33309e-19 $X=0.063 $Y=0.1355 $X2=0.666 $Y2=0.234
cc_45 N_A_c_1_p Y 0.00101871f $X=0.621 $Y=0.135 $X2=0.6775 $Y2=0.1475

* END of "./INVx11_ASAP7_75t_SRAM.pex.sp.INVX11_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVx13_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:33:07 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVx13_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVx13_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVx13_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:33:07 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVX13_ASAP7_75T_SRAM%A 2 7 10 15 18 23 26 31 34 39 42 47 50 55 58 63 66
+ 71 74 79 82 87 90 95 98 101 103 115 VSS
c53 115 VSS 0.0275217f $X=0.066 $Y=0.1365
c54 101 VSS 0.0683982f $X=0.729 $Y=0.135
c55 98 VSS 0.0678263f $X=0.729 $Y=0.0675
c56 90 VSS 0.0643964f $X=0.675 $Y=0.0675
c57 82 VSS 0.0642127f $X=0.621 $Y=0.0675
c58 74 VSS 0.0642127f $X=0.567 $Y=0.0675
c59 66 VSS 0.0642127f $X=0.513 $Y=0.0675
c60 58 VSS 0.0642127f $X=0.459 $Y=0.0675
c61 50 VSS 0.0642127f $X=0.405 $Y=0.0675
c62 42 VSS 0.0642127f $X=0.351 $Y=0.0675
c63 34 VSS 0.0642127f $X=0.297 $Y=0.0675
c64 26 VSS 0.0642127f $X=0.243 $Y=0.0675
c65 18 VSS 0.0642127f $X=0.189 $Y=0.0675
c66 10 VSS 0.0644226f $X=0.135 $Y=0.0675
c67 2 VSS 0.0655089f $X=0.081 $Y=0.0675
r68 112 115 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135
+ $X2=0.064 $Y2=0.135
r69 101 103 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.135 $X2=0.729 $Y2=0.2025
r70 98 101 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.135
r71 93 101 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.729 $Y2=0.135
r72 93 95 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.2025
r73 90 93 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0675 $X2=0.675 $Y2=0.135
r74 85 93 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621
+ $Y=0.135 $X2=0.675 $Y2=0.135
r75 85 87 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r76 82 85 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
r77 77 85 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.567
+ $Y=0.135 $X2=0.621 $Y2=0.135
r78 77 79 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r79 74 77 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r80 69 77 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r81 69 71 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r82 66 69 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
r83 61 69 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r84 61 63 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r85 58 61 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r86 53 61 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r87 53 55 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r88 50 53 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
r89 45 53 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r90 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r91 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r92 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r93 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r94 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r95 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r96 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r97 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r98 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r99 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r100 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.189 $Y=0.0675 $X2=0.189 $Y2=0.135
r101 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r102 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r103 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r104 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r105 5 112 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r106 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r107 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVX13_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 21 22 26 27 31 36 37 40 41
+ 42 45 46 47 50 51 52 55 56 57 60 61 62 65 66 71 74 78 81 84 87 90 94 120 VSS
c53 120 VSS 0.00874864f $X=0.7825 $Y=0.1475
c54 94 VSS 0.0796806f $X=0.774 $Y=0.234
c55 93 VSS 0.00692279f $X=0.756 $Y=0.036
c56 90 VSS 0.00928905f $X=0.648 $Y=0.036
c57 87 VSS 0.00928955f $X=0.54 $Y=0.036
c58 84 VSS 0.00928955f $X=0.432 $Y=0.036
c59 81 VSS 0.00928955f $X=0.324 $Y=0.036
c60 78 VSS 0.00928954f $X=0.216 $Y=0.036
c61 74 VSS 0.00904082f $X=0.108 $Y=0.036
c62 71 VSS 0.0796806f $X=0.774 $Y=0.036
c63 69 VSS 0.00730645f $X=0.754 $Y=0.2025
c64 65 VSS 0.00928905f $X=0.648 $Y=0.2025
c65 61 VSS 5.38922e-19 $X=0.665 $Y=0.2025
c66 60 VSS 0.00928955f $X=0.54 $Y=0.2025
c67 56 VSS 5.38922e-19 $X=0.557 $Y=0.2025
c68 55 VSS 0.00928955f $X=0.432 $Y=0.2025
c69 51 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c70 50 VSS 0.00928955f $X=0.324 $Y=0.2025
c71 46 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c72 45 VSS 0.00928954f $X=0.216 $Y=0.2025
c73 41 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c74 40 VSS 0.00904082f $X=0.108 $Y=0.2025
c75 36 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c76 34 VSS 3.8366e-19 $X=0.754 $Y=0.0675
c77 26 VSS 5.38922e-19 $X=0.665 $Y=0.0675
c78 21 VSS 5.38922e-19 $X=0.557 $Y=0.0675
c79 16 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c80 11 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c81 6 VSS 5.38922e-19 $X=0.233 $Y=0.0675
c82 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r83 118 120 5.26235 $w=1.8e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.783
+ $Y=0.225 $X2=0.783 $Y2=0.1475
r84 117 120 6.95988 $w=1.8e-08 $l=1.025e-07 $layer=M1 $thickness=3.6e-08
+ $X=0.783 $Y=0.045 $X2=0.783 $Y2=0.1475
r85 112 115 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.756 $Y2=0.234
r86 109 112 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.648 $Y2=0.234
r87 106 109 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.54 $Y2=0.234
r88 103 106 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r89 100 103 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.324 $Y2=0.234
r90 96 100 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.216 $Y2=0.234
r91 94 118 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.774 $Y=0.234 $X2=0.783 $Y2=0.225
r92 94 115 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.234 $X2=0.756 $Y2=0.234
r93 92 93 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r94 89 92 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.756 $Y2=0.036
r95 89 90 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036 $X2=0.648
+ $Y2=0.036
r96 86 89 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.648 $Y2=0.036
r97 86 87 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r98 83 86 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.54 $Y2=0.036
r99 83 84 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r100 80 83 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r101 80 81 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r102 77 80 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.324 $Y2=0.036
r103 77 78 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r104 73 77 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.216 $Y2=0.036
r105 73 74 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r106 71 117 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.774 $Y=0.036 $X2=0.783 $Y2=0.045
r107 71 92 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.774
+ $Y=0.036 $X2=0.756 $Y2=0.036
r108 69 115 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234
+ $X2=0.756 $Y2=0.234
r109 66 69 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.754 $Y2=0.2025
r110 65 112 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234
+ $X2=0.648 $Y2=0.234
r111 62 65 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.648 $Y2=0.2025
r112 61 65 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.648 $Y2=0.2025
r113 60 109 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r114 57 60 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r115 56 60 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r116 55 106 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r117 52 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r118 51 55 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r119 50 103 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r120 47 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r121 46 50 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r122 45 100 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r123 42 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r124 41 45 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r125 40 96 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r126 37 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r127 36 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r128 34 93 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.756 $Y=0.0675 $X2=0.756 $Y2=0.036
r129 31 34 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.754 $Y2=0.0675
r130 30 90 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.648 $Y=0.0675 $X2=0.648 $Y2=0.036
r131 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.648 $Y2=0.0675
r132 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0675 $X2=0.648 $Y2=0.0675
r133 25 87 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r134 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r135 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r136 20 84 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r137 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r138 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r139 15 81 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r140 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r141 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r142 10 78 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.216 $Y=0.0675 $X2=0.216 $Y2=0.036
r143 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r144 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r145 5 74 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r146 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r147 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./INVx13_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVx13_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_A_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_A_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_A_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_A_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_A_M6_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_A_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_A_M8_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_A_M9_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 N_Y_M10_d N_A_M10_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M11 N_Y_M11_d N_A_M11_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M12 N_Y_M12_d N_A_M12_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M13 N_Y_M13_d N_A_M13_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M14 N_Y_M14_d N_A_M14_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M15 N_Y_M15_d N_A_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M16 N_Y_M16_d N_A_M16_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M17 N_Y_M17_d N_A_M17_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M18 N_Y_M18_d N_A_M18_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M19 N_Y_M19_d N_A_M19_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M20 N_Y_M20_d N_A_M20_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M21 N_Y_M21_d N_A_M21_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M22 N_Y_M22_d N_A_M22_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M23 N_Y_M23_d N_A_M23_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M24 N_Y_M24_d N_A_M24_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
M25 N_Y_M25_d N_A_M25_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
*
* 
* .include "INVx13_ASAP7_75t_SRAM.pex.sp.INVX13_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVx13_ASAP7_75t_SRAM.pex.sp.INVX13_ASAP7_75T_SRAM.pxi"
* File: INVx13_ASAP7_75t_SRAM.pex.sp.INVX13_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:33:07 2017
* 
x_PM_INVX13_ASAP7_75T_SRAM%A N_A_M0_g N_A_M13_g N_A_M1_g N_A_M14_g N_A_M2_g
+ N_A_M15_g N_A_M3_g N_A_M16_g N_A_M4_g N_A_M17_g N_A_M5_g N_A_M18_g N_A_M6_g
+ N_A_M19_g N_A_M7_g N_A_M20_g N_A_M8_g N_A_M21_g N_A_M9_g N_A_M22_g N_A_M10_g
+ N_A_M23_g N_A_M11_g N_A_M24_g N_A_M12_g N_A_c_1_p N_A_M25_g A VSS
+ PM_INVX13_ASAP7_75T_SRAM%A
x_PM_INVX13_ASAP7_75T_SRAM%Y N_Y_M1_d N_Y_M0_d N_Y_M3_d N_Y_M2_d N_Y_M5_d N_Y_M4_d
+ N_Y_M7_d N_Y_M6_d N_Y_M9_d N_Y_M8_d N_Y_M11_d N_Y_M10_d N_Y_M12_d N_Y_M14_d
+ N_Y_M13_d N_Y_c_61_n N_Y_M16_d N_Y_M15_d N_Y_c_63_n N_Y_M18_d N_Y_M17_d
+ N_Y_c_65_n N_Y_M20_d N_Y_M19_d N_Y_c_67_n N_Y_M22_d N_Y_M21_d N_Y_c_69_n
+ N_Y_M24_d N_Y_M23_d N_Y_c_71_n N_Y_M25_d N_Y_c_72_n N_Y_c_86_n N_Y_c_87_n
+ N_Y_c_88_n N_Y_c_89_n N_Y_c_90_n N_Y_c_91_n N_Y_c_92_n Y VSS
+ PM_INVX13_ASAP7_75T_SRAM%Y
cc_1 N_A_c_1_p N_Y_M1_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_2 N_A_c_1_p N_Y_M3_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.233 $Y2=0.0675
cc_3 N_A_c_1_p N_Y_M5_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.341 $Y2=0.0675
cc_4 N_A_c_1_p N_Y_M7_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.449 $Y2=0.0675
cc_5 N_A_c_1_p N_Y_M9_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.557 $Y2=0.0675
cc_6 N_A_c_1_p N_Y_M11_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.665 $Y2=0.0675
cc_7 N_A_c_1_p N_Y_M14_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_8 N_A_c_1_p N_Y_c_61_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_9 N_A_c_1_p N_Y_M16_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.233 $Y2=0.2025
cc_10 N_A_c_1_p N_Y_c_63_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.216 $Y2=0.2025
cc_11 N_A_c_1_p N_Y_M18_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.341 $Y2=0.2025
cc_12 N_A_c_1_p N_Y_c_65_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.324 $Y2=0.2025
cc_13 N_A_c_1_p N_Y_M20_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.449 $Y2=0.2025
cc_14 N_A_c_1_p N_Y_c_67_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.432 $Y2=0.2025
cc_15 N_A_c_1_p N_Y_M22_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.557 $Y2=0.2025
cc_16 N_A_c_1_p N_Y_c_69_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.54 $Y2=0.2025
cc_17 N_A_c_1_p N_Y_M24_d 3.80663e-19 $X=0.729 $Y=0.135 $X2=0.665 $Y2=0.2025
cc_18 N_A_c_1_p N_Y_c_71_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.648 $Y2=0.2025
cc_19 N_A_M1_g N_Y_c_72_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_20 N_A_M2_g N_Y_c_72_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_21 N_A_M3_g N_Y_c_72_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_22 N_A_M4_g N_Y_c_72_n 4.59284e-19 $X=0.297 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_23 N_A_M5_g N_Y_c_72_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_24 N_A_M6_g N_Y_c_72_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_25 N_A_M7_g N_Y_c_72_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_26 N_A_M8_g N_Y_c_72_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_27 N_A_M9_g N_Y_c_72_n 4.59284e-19 $X=0.567 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_28 N_A_M10_g N_Y_c_72_n 4.59284e-19 $X=0.621 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_29 N_A_M11_g N_Y_c_72_n 4.59284e-19 $X=0.675 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_30 N_A_M12_g N_Y_c_72_n 4.59284e-19 $X=0.729 $Y=0.0675 $X2=0.774 $Y2=0.036
cc_31 N_A_c_1_p N_Y_c_72_n 0.00817348f $X=0.729 $Y=0.135 $X2=0.774 $Y2=0.036
cc_32 A N_Y_c_72_n 5.33584e-19 $X=0.066 $Y=0.1365 $X2=0.774 $Y2=0.036
cc_33 N_A_c_1_p N_Y_c_86_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.108 $Y2=0.036
cc_34 N_A_c_1_p N_Y_c_87_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.216 $Y2=0.036
cc_35 N_A_c_1_p N_Y_c_88_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.324 $Y2=0.036
cc_36 N_A_c_1_p N_Y_c_89_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.432 $Y2=0.036
cc_37 N_A_c_1_p N_Y_c_90_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.54 $Y2=0.036
cc_38 N_A_c_1_p N_Y_c_91_n 8.00061e-19 $X=0.729 $Y=0.135 $X2=0.648 $Y2=0.036
cc_39 N_A_M1_g N_Y_c_92_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_40 N_A_M2_g N_Y_c_92_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_41 N_A_M3_g N_Y_c_92_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_42 N_A_M4_g N_Y_c_92_n 4.59284e-19 $X=0.297 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_43 N_A_M5_g N_Y_c_92_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_44 N_A_M6_g N_Y_c_92_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_45 N_A_M7_g N_Y_c_92_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_46 N_A_M8_g N_Y_c_92_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_47 N_A_M9_g N_Y_c_92_n 4.59284e-19 $X=0.567 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_48 N_A_M10_g N_Y_c_92_n 4.59284e-19 $X=0.621 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_49 N_A_M11_g N_Y_c_92_n 4.59284e-19 $X=0.675 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_50 N_A_M12_g N_Y_c_92_n 4.59284e-19 $X=0.729 $Y=0.0675 $X2=0.774 $Y2=0.234
cc_51 N_A_c_1_p N_Y_c_92_n 0.00817348f $X=0.729 $Y=0.135 $X2=0.774 $Y2=0.234
cc_52 A N_Y_c_92_n 5.33584e-19 $X=0.066 $Y=0.1365 $X2=0.774 $Y2=0.234
cc_53 N_A_c_1_p Y 0.00103293f $X=0.729 $Y=0.135 $X2=0.7825 $Y2=0.1475

* END of "./INVx13_ASAP7_75t_SRAM.pex.sp.INVX13_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVx1_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:33:30 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVx1_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVx1_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVx1_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:33:30 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVX1_ASAP7_75T_SRAM%A 2 7 15 19 VSS
c5 19 VSS 9.16094e-19 $X=0.064 $Y=0.135
c6 15 VSS 0.0241737f $X=0.047 $Y=0.1365
c7 5 VSS 0.00713947f $X=0.081 $Y=0.135
c8 2 VSS 0.0702997f $X=0.081 $Y=0.0675
r9 19 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r10 15 19 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.047
+ $Y=0.135 $X2=0.064 $Y2=0.135
r11 5 20 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r12 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r13 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVX1_ASAP7_75T_SRAM%Y 1 6 12 14 16 22 30 VSS
c5 30 VSS 0.00413618f $X=0.126 $Y=0.234
c6 29 VSS 0.00278493f $X=0.135 $Y=0.234
c7 22 VSS 0.00413618f $X=0.126 $Y=0.036
c8 21 VSS 0.00278493f $X=0.135 $Y=0.036
c9 19 VSS 0.0065018f $X=0.108 $Y=0.036
c10 16 VSS 7.74764e-19 $X=0.135 $Y=0.144
c11 14 VSS 0.00405481f $X=0.1355 $Y=0.1145
c12 12 VSS 0.0038739f $X=0.135 $Y=0.225
c13 9 VSS 0.00688074f $X=0.106 $Y=0.2025
c14 4 VSS 3.7894e-19 $X=0.106 $Y=0.0675
r15 30 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r16 29 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r17 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r18 22 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r19 21 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r20 18 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r21 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r22 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.144
r23 14 15 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.1145 $X2=0.135 $Y2=0.126
r24 12 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.234
r25 12 16 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.144
r26 11 21 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.036
r27 11 14 4.71914 $w=1.8e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.1145
r28 9 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r29 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.2025 $X2=0.106 $Y2=0.2025
r30 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r31 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.106 $Y2=0.0675
.ends


* END of "./INVx1_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVx1_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
*
* 
* .include "INVx1_ASAP7_75t_SRAM.pex.sp.INVX1_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVx1_ASAP7_75t_SRAM.pex.sp.INVX1_ASAP7_75T_SRAM.pxi"
* File: INVx1_ASAP7_75t_SRAM.pex.sp.INVX1_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:33:30 2017
* 
x_PM_INVX1_ASAP7_75T_SRAM%A N_A_M0_g N_A_M1_g A N_A_c_3_p VSS
+ PM_INVX1_ASAP7_75T_SRAM%A
x_PM_INVX1_ASAP7_75T_SRAM%Y N_Y_M0_d N_Y_M1_d N_Y_c_6_n Y N_Y_c_8_n N_Y_c_9_n
+ N_Y_c_10_n VSS PM_INVX1_ASAP7_75T_SRAM%Y
cc_1 A N_Y_c_6_n 6.7994e-19 $X=0.047 $Y=0.1365 $X2=0.135 $Y2=0.225
cc_2 A Y 6.7994e-19 $X=0.047 $Y=0.1365 $X2=0.1355 $Y2=0.1145
cc_3 N_A_c_3_p N_Y_c_8_n 5.19281e-19 $X=0.064 $Y=0.135 $X2=0.135 $Y2=0.144
cc_4 A N_Y_c_9_n 5.53308e-19 $X=0.047 $Y=0.1365 $X2=0.126 $Y2=0.036
cc_5 A N_Y_c_10_n 5.53308e-19 $X=0.047 $Y=0.1365 $X2=0.126 $Y2=0.234

* END of "./INVx1_ASAP7_75t_SRAM.pex.sp.INVX1_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVx2_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:33:52 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVx2_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVx2_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVx2_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:33:52 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVX2_ASAP7_75T_SRAM%A 2 7 10 13 15 23 VSS
c13 28 VSS 4.99695e-19 $X=0.055 $Y=0.135
c14 27 VSS 9.69018e-19 $X=0.046 $Y=0.135
c15 25 VSS 6.28633e-19 $X=0.064 $Y=0.135
c16 23 VSS 0.0241049f $X=0.042 $Y=0.1345
c17 13 VSS 0.00898269f $X=0.135 $Y=0.135
c18 10 VSS 0.0641916f $X=0.135 $Y=0.0675
c19 2 VSS 0.0651658f $X=0.081 $Y=0.0675
r20 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.055 $Y2=0.135
r21 25 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.135 $X2=0.055 $Y2=0.135
r22 25 26 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r23 23 27 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.042
+ $Y=0.135 $X2=0.046 $Y2=0.135
r24 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r25 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r26 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r27 5 26 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r28 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r29 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVX2_ASAP7_75T_SRAM%Y 1 2 6 7 10 11 14 16 24 25 VSS
c13 26 VSS 9.75657e-19 $X=0.189 $Y=0.144
c14 25 VSS 0.0047383f $X=0.189 $Y=0.126
c15 24 VSS 0.0047383f $X=0.189 $Y=0.1475
c16 16 VSS 0.0145004f $X=0.18 $Y=0.234
c17 14 VSS 0.00904881f $X=0.108 $Y=0.036
c18 11 VSS 0.0145004f $X=0.18 $Y=0.036
c19 10 VSS 0.00904881f $X=0.108 $Y=0.2025
c20 6 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c21 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r22 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.144
r23 24 26 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.1475 $X2=0.189 $Y2=0.144
r24 22 24 5.26235 $w=1.8e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.1475
r25 21 25 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.126
r26 16 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.234 $X2=0.189 $Y2=0.225
r27 16 18 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.108 $Y2=0.234
r28 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r29 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r30 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.108 $Y2=0.036
r31 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r32 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r33 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r34 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r35 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r36 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./INVx2_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVx2_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_A_M2_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M3 N_Y_M3_d N_A_M3_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
*
* 
* .include "INVx2_ASAP7_75t_SRAM.pex.sp.INVX2_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVx2_ASAP7_75t_SRAM.pex.sp.INVX2_ASAP7_75T_SRAM.pxi"
* File: INVx2_ASAP7_75t_SRAM.pex.sp.INVX2_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:33:52 2017
* 
x_PM_INVX2_ASAP7_75T_SRAM%A N_A_M0_g N_A_M2_g N_A_M1_g N_A_c_1_p N_A_M3_g A VSS
+ PM_INVX2_ASAP7_75T_SRAM%A
x_PM_INVX2_ASAP7_75T_SRAM%Y N_Y_M1_d N_Y_M0_d N_Y_M3_d N_Y_M2_d N_Y_c_16_n
+ N_Y_c_17_n N_Y_c_20_n N_Y_c_21_n Y N_Y_c_25_n VSS PM_INVX2_ASAP7_75T_SRAM%Y
cc_1 N_A_c_1_p N_Y_M1_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_2 N_A_c_1_p N_Y_M3_d 3.80663e-19 $X=0.135 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_3 N_A_c_1_p N_Y_c_16_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_4 N_A_M1_g N_Y_c_17_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.18 $Y2=0.036
cc_5 N_A_c_1_p N_Y_c_17_n 5.51214e-19 $X=0.135 $Y=0.135 $X2=0.18 $Y2=0.036
cc_6 A N_Y_c_17_n 5.24213e-19 $X=0.042 $Y=0.1345 $X2=0.18 $Y2=0.036
cc_7 N_A_c_1_p N_Y_c_20_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.108 $Y2=0.036
cc_8 N_A_M1_g N_Y_c_21_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.18 $Y2=0.234
cc_9 N_A_c_1_p N_Y_c_21_n 5.51214e-19 $X=0.135 $Y=0.135 $X2=0.18 $Y2=0.234
cc_10 A N_Y_c_21_n 5.24213e-19 $X=0.042 $Y=0.1345 $X2=0.18 $Y2=0.234
cc_11 A Y 2.97507e-19 $X=0.042 $Y=0.1345 $X2=0.189 $Y2=0.1475
cc_12 N_A_c_1_p N_Y_c_25_n 5.14102e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.126
cc_13 A N_Y_c_25_n 2.97507e-19 $X=0.042 $Y=0.1345 $X2=0.189 $Y2=0.126

* END of "./INVx2_ASAP7_75t_SRAM.pex.sp.INVX2_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVx3_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:34:14 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVx3_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVx3_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVx3_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:34:14 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVX3_ASAP7_75T_SRAM%A 2 7 10 15 18 21 23 31 VSS
c13 31 VSS 0.0276577f $X=0.062 $Y=0.1335
c14 21 VSS 0.0172079f $X=0.189 $Y=0.135
c15 18 VSS 0.0678263f $X=0.189 $Y=0.0675
c16 10 VSS 0.0646063f $X=0.135 $Y=0.0675
c17 2 VSS 0.0655089f $X=0.081 $Y=0.0675
r18 31 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r19 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r20 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r21 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r22 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r23 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r24 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r25 5 35 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVX3_ASAP7_75T_SRAM%Y 1 2 6 11 12 15 16 21 24 29 40 41 VSS
c13 42 VSS 8.99665e-19 $X=0.243 $Y=0.144
c14 41 VSS 0.00398275f $X=0.243 $Y=0.126
c15 40 VSS 0.00398275f $X=0.2445 $Y=0.1465
c16 29 VSS 0.01958f $X=0.234 $Y=0.234
c17 28 VSS 0.00692279f $X=0.216 $Y=0.036
c18 24 VSS 0.00904032f $X=0.108 $Y=0.036
c19 21 VSS 0.01958f $X=0.234 $Y=0.036
c20 19 VSS 0.00726838f $X=0.214 $Y=0.2025
c21 15 VSS 0.00904032f $X=0.108 $Y=0.2025
c22 11 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c23 9 VSS 3.45593e-19 $X=0.214 $Y=0.0675
c24 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r25 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.144
r26 40 42 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.1465 $X2=0.243 $Y2=0.144
r27 38 40 5.33025 $w=1.8e-08 $l=7.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.1465
r28 37 41 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.126
r29 31 35 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.216 $Y2=0.234
r30 29 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r31 29 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r32 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r33 23 27 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.216 $Y2=0.036
r34 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r35 21 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r36 21 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r37 19 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r38 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.214 $Y2=0.2025
r39 15 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r40 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r41 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r42 9 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r43 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.214 $Y2=0.0675
r44 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r45 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r46 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./INVx3_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVx3_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_A_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_A_M3_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M4 N_Y_M4_d N_A_M4_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M5 N_Y_M5_d N_A_M5_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
*
* 
* .include "INVx3_ASAP7_75t_SRAM.pex.sp.INVX3_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVx3_ASAP7_75t_SRAM.pex.sp.INVX3_ASAP7_75T_SRAM.pxi"
* File: INVx3_ASAP7_75t_SRAM.pex.sp.INVX3_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:34:14 2017
* 
x_PM_INVX3_ASAP7_75T_SRAM%A N_A_M0_g N_A_M3_g N_A_M1_g N_A_M4_g N_A_M2_g N_A_c_1_p
+ N_A_M5_g A VSS PM_INVX3_ASAP7_75T_SRAM%A
x_PM_INVX3_ASAP7_75T_SRAM%Y N_Y_M1_d N_Y_M0_d N_Y_M2_d N_Y_M4_d N_Y_M3_d N_Y_c_16_n
+ N_Y_M5_d N_Y_c_17_n N_Y_c_21_n N_Y_c_22_n Y N_Y_c_26_n VSS
+ PM_INVX3_ASAP7_75T_SRAM%Y
cc_1 N_A_c_1_p N_Y_M1_d 3.80663e-19 $X=0.189 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_2 N_A_c_1_p N_Y_M4_d 3.80663e-19 $X=0.189 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_3 N_A_c_1_p N_Y_c_16_n 8.00061e-19 $X=0.189 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_4 N_A_M1_g N_Y_c_17_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.234 $Y2=0.036
cc_5 N_A_M2_g N_Y_c_17_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.234 $Y2=0.036
cc_6 N_A_c_1_p N_Y_c_17_n 0.00134609f $X=0.189 $Y=0.135 $X2=0.234 $Y2=0.036
cc_7 A N_Y_c_17_n 5.28865e-19 $X=0.062 $Y=0.1335 $X2=0.234 $Y2=0.036
cc_8 N_A_c_1_p N_Y_c_21_n 8.00061e-19 $X=0.189 $Y=0.135 $X2=0.108 $Y2=0.036
cc_9 N_A_M1_g N_Y_c_22_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.234 $Y2=0.234
cc_10 N_A_M2_g N_Y_c_22_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.234 $Y2=0.234
cc_11 N_A_c_1_p N_Y_c_22_n 0.00134609f $X=0.189 $Y=0.135 $X2=0.234 $Y2=0.234
cc_12 A N_Y_c_22_n 5.28865e-19 $X=0.062 $Y=0.1335 $X2=0.234 $Y2=0.234
cc_13 N_A_c_1_p N_Y_c_26_n 5.51266e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.126

* END of "./INVx3_ASAP7_75t_SRAM.pex.sp.INVX3_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVx4_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:34:37 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVx4_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVx4_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVx4_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:34:37 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVX4_ASAP7_75T_SRAM%A 2 7 10 15 18 23 26 29 31 39 VSS
c19 39 VSS 0.0276205f $X=0.062 $Y=0.1345
c20 29 VSS 0.0190713f $X=0.243 $Y=0.135
c21 26 VSS 0.0645347f $X=0.243 $Y=0.0675
c22 18 VSS 0.0644226f $X=0.189 $Y=0.0675
c23 10 VSS 0.0644226f $X=0.135 $Y=0.0675
c24 2 VSS 0.0655089f $X=0.081 $Y=0.0675
r25 39 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r26 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r27 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r28 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r29 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r30 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r31 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r32 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r33 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r34 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r35 5 43 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r36 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r37 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVX4_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 15 16 17 20 21 24 28 29 40 41 VSS
c19 42 VSS 7.62145e-19 $X=0.297 $Y=0.144
c20 41 VSS 0.00529405f $X=0.297 $Y=0.126
c21 40 VSS 0.00529405f $X=0.2965 $Y=0.1465
c22 29 VSS 0.0266097f $X=0.288 $Y=0.234
c23 28 VSS 0.00929751f $X=0.216 $Y=0.036
c24 24 VSS 0.00904081f $X=0.108 $Y=0.036
c25 21 VSS 0.0266097f $X=0.288 $Y=0.036
c26 20 VSS 0.00929751f $X=0.216 $Y=0.2025
c27 16 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c28 15 VSS 0.00904081f $X=0.108 $Y=0.2025
c29 11 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c30 6 VSS 5.38922e-19 $X=0.233 $Y=0.0675
c31 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r32 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.144
r33 40 42 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1465 $X2=0.297 $Y2=0.144
r34 38 40 5.33025 $w=1.8e-08 $l=7.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.1465
r35 37 41 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.126
r36 31 35 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.216 $Y2=0.234
r37 29 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.234 $X2=0.297 $Y2=0.225
r38 29 35 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.216 $Y2=0.234
r39 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r40 23 27 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.216 $Y2=0.036
r41 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r42 21 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r43 21 27 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.216 $Y2=0.036
r44 20 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r45 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r46 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r47 15 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r48 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r49 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r50 10 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r51 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r52 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r53 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r54 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r55 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./INVx4_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVx4_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_A_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_A_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_A_M4_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M5 N_Y_M5_d N_A_M5_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M6 N_Y_M6_d N_A_M6_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M7 N_Y_M7_d N_A_M7_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
*
* 
* .include "INVx4_ASAP7_75t_SRAM.pex.sp.INVX4_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVx4_ASAP7_75t_SRAM.pex.sp.INVX4_ASAP7_75T_SRAM.pxi"
* File: INVx4_ASAP7_75t_SRAM.pex.sp.INVX4_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:34:37 2017
* 
x_PM_INVX4_ASAP7_75T_SRAM%A N_A_M0_g N_A_M4_g N_A_M1_g N_A_M5_g N_A_M2_g N_A_M6_g
+ N_A_M3_g N_A_c_1_p N_A_M7_g A VSS PM_INVX4_ASAP7_75T_SRAM%A
x_PM_INVX4_ASAP7_75T_SRAM%Y N_Y_M1_d N_Y_M0_d N_Y_M3_d N_Y_M2_d N_Y_M5_d N_Y_M4_d
+ N_Y_c_23_n N_Y_M7_d N_Y_M6_d N_Y_c_25_n N_Y_c_26_n N_Y_c_31_n N_Y_c_32_n
+ N_Y_c_33_n Y N_Y_c_38_n VSS PM_INVX4_ASAP7_75T_SRAM%Y
cc_1 N_A_c_1_p N_Y_M1_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_2 N_A_c_1_p N_Y_M3_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.233 $Y2=0.0675
cc_3 N_A_c_1_p N_Y_M5_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_4 N_A_c_1_p N_Y_c_23_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_5 N_A_c_1_p N_Y_M7_d 3.80663e-19 $X=0.243 $Y=0.135 $X2=0.233 $Y2=0.2025
cc_6 N_A_c_1_p N_Y_c_25_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.216 $Y2=0.2025
cc_7 N_A_M1_g N_Y_c_26_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.288 $Y2=0.036
cc_8 N_A_M2_g N_Y_c_26_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.288 $Y2=0.036
cc_9 N_A_M3_g N_Y_c_26_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.288 $Y2=0.036
cc_10 N_A_c_1_p N_Y_c_26_n 0.00191346f $X=0.243 $Y=0.135 $X2=0.288 $Y2=0.036
cc_11 A N_Y_c_26_n 5.30329e-19 $X=0.062 $Y=0.1345 $X2=0.288 $Y2=0.036
cc_12 N_A_c_1_p N_Y_c_31_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.108 $Y2=0.036
cc_13 N_A_c_1_p N_Y_c_32_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.216 $Y2=0.036
cc_14 N_A_M1_g N_Y_c_33_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.288 $Y2=0.234
cc_15 N_A_M2_g N_Y_c_33_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.288 $Y2=0.234
cc_16 N_A_M3_g N_Y_c_33_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.288 $Y2=0.234
cc_17 N_A_c_1_p N_Y_c_33_n 0.00191346f $X=0.243 $Y=0.135 $X2=0.288 $Y2=0.234
cc_18 A N_Y_c_33_n 5.30329e-19 $X=0.062 $Y=0.1345 $X2=0.288 $Y2=0.234
cc_19 N_A_c_1_p N_Y_c_38_n 5.76695e-19 $X=0.243 $Y=0.135 $X2=0.297 $Y2=0.126

* END of "./INVx4_ASAP7_75t_SRAM.pex.sp.INVX4_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVx5_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:34:59 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVx5_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVx5_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVx5_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:34:59 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVX5_ASAP7_75T_SRAM%A 2 7 10 15 18 23 26 31 34 37 39 51 VSS
c21 51 VSS 0.0275217f $X=0.066 $Y=0.1345
c22 37 VSS 0.0276912f $X=0.297 $Y=0.135
c23 34 VSS 0.0678263f $X=0.297 $Y=0.0675
c24 26 VSS 0.0643964f $X=0.243 $Y=0.0675
c25 18 VSS 0.0642127f $X=0.189 $Y=0.0675
c26 10 VSS 0.0644226f $X=0.135 $Y=0.0675
c27 2 VSS 0.0655089f $X=0.081 $Y=0.0675
r28 48 51 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r29 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r30 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r31 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r32 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r33 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r34 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r35 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r36 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r37 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r38 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r39 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r40 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r41 5 48 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r42 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r43 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVX5_ASAP7_75T_SRAM%Y 1 2 6 7 11 16 17 20 21 22 25 26 31 34 38 42 56 57
+ VSS
c21 58 VSS 7.62145e-19 $X=0.351 $Y=0.144
c22 57 VSS 0.00398275f $X=0.351 $Y=0.126
c23 56 VSS 0.00398275f $X=0.3515 $Y=0.1475
c24 42 VSS 0.0315875f $X=0.342 $Y=0.234
c25 41 VSS 0.00692279f $X=0.324 $Y=0.036
c26 38 VSS 0.00928904f $X=0.216 $Y=0.036
c27 34 VSS 0.00904082f $X=0.108 $Y=0.036
c28 31 VSS 0.0315875f $X=0.342 $Y=0.036
c29 29 VSS 0.00726838f $X=0.322 $Y=0.2025
c30 25 VSS 0.00928904f $X=0.216 $Y=0.2025
c31 21 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c32 20 VSS 0.00904082f $X=0.108 $Y=0.2025
c33 16 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c34 14 VSS 3.45593e-19 $X=0.322 $Y=0.0675
c35 6 VSS 5.38922e-19 $X=0.233 $Y=0.0675
c36 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r37 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.144
r38 56 58 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1475 $X2=0.351 $Y2=0.144
r39 54 56 5.26235 $w=1.8e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.1475
r40 53 57 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.126
r41 48 51 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.324 $Y2=0.234
r42 44 48 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.216 $Y2=0.234
r43 42 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.234 $X2=0.351 $Y2=0.225
r44 42 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.324 $Y2=0.234
r45 40 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r46 37 40 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.324 $Y2=0.036
r47 37 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r48 33 37 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.216 $Y2=0.036
r49 33 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r50 31 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.036 $X2=0.351 $Y2=0.045
r51 31 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.324 $Y2=0.036
r52 29 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r53 26 29 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.322 $Y2=0.2025
r54 25 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r55 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r56 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r57 20 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r58 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r59 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r60 14 41 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r61 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.322 $Y2=0.0675
r62 10 38 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r63 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r64 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r65 5 34 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r66 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r67 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./INVx5_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVx5_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_A_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_A_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_A_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_A_M5_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M6 N_Y_M6_d N_A_M6_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M7 N_Y_M7_d N_A_M7_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M8 N_Y_M8_d N_A_M8_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M9 N_Y_M9_d N_A_M9_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
*
* 
* .include "INVx5_ASAP7_75t_SRAM.pex.sp.INVX5_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVx5_ASAP7_75t_SRAM.pex.sp.INVX5_ASAP7_75T_SRAM.pxi"
* File: INVx5_ASAP7_75t_SRAM.pex.sp.INVX5_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:34:59 2017
* 
x_PM_INVX5_ASAP7_75T_SRAM%A N_A_M0_g N_A_M5_g N_A_M1_g N_A_M6_g N_A_M2_g N_A_M7_g
+ N_A_M3_g N_A_M8_g N_A_M4_g N_A_c_1_p N_A_M9_g A VSS PM_INVX5_ASAP7_75T_SRAM%A
x_PM_INVX5_ASAP7_75T_SRAM%Y N_Y_M1_d N_Y_M0_d N_Y_M3_d N_Y_M2_d N_Y_M4_d N_Y_M6_d
+ N_Y_M5_d N_Y_c_25_n N_Y_M8_d N_Y_M7_d N_Y_c_27_n N_Y_M9_d N_Y_c_28_n
+ N_Y_c_34_n N_Y_c_35_n N_Y_c_36_n Y N_Y_c_42_n VSS PM_INVX5_ASAP7_75T_SRAM%Y
cc_1 N_A_c_1_p N_Y_M1_d 3.80663e-19 $X=0.297 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_2 N_A_c_1_p N_Y_M3_d 3.80663e-19 $X=0.297 $Y=0.135 $X2=0.233 $Y2=0.0675
cc_3 N_A_c_1_p N_Y_M6_d 3.80663e-19 $X=0.297 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_4 N_A_c_1_p N_Y_c_25_n 8.00061e-19 $X=0.297 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_5 N_A_c_1_p N_Y_M8_d 3.80663e-19 $X=0.297 $Y=0.135 $X2=0.233 $Y2=0.2025
cc_6 N_A_c_1_p N_Y_c_27_n 8.00061e-19 $X=0.297 $Y=0.135 $X2=0.216 $Y2=0.2025
cc_7 N_A_M1_g N_Y_c_28_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.342 $Y2=0.036
cc_8 N_A_M2_g N_Y_c_28_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.342 $Y2=0.036
cc_9 N_A_M3_g N_Y_c_28_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.342 $Y2=0.036
cc_10 N_A_M4_g N_Y_c_28_n 4.59284e-19 $X=0.297 $Y=0.0675 $X2=0.342 $Y2=0.036
cc_11 N_A_c_1_p N_Y_c_28_n 0.00270834f $X=0.297 $Y=0.135 $X2=0.342 $Y2=0.036
cc_12 A N_Y_c_28_n 5.31238e-19 $X=0.066 $Y=0.1345 $X2=0.342 $Y2=0.036
cc_13 N_A_c_1_p N_Y_c_34_n 8.00061e-19 $X=0.297 $Y=0.135 $X2=0.108 $Y2=0.036
cc_14 N_A_c_1_p N_Y_c_35_n 8.00061e-19 $X=0.297 $Y=0.135 $X2=0.216 $Y2=0.036
cc_15 N_A_M1_g N_Y_c_36_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.342 $Y2=0.234
cc_16 N_A_M2_g N_Y_c_36_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.342 $Y2=0.234
cc_17 N_A_M3_g N_Y_c_36_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.342 $Y2=0.234
cc_18 N_A_M4_g N_Y_c_36_n 4.59284e-19 $X=0.297 $Y=0.0675 $X2=0.342 $Y2=0.234
cc_19 N_A_c_1_p N_Y_c_36_n 0.00270834f $X=0.297 $Y=0.135 $X2=0.342 $Y2=0.234
cc_20 A N_Y_c_36_n 5.31238e-19 $X=0.066 $Y=0.1345 $X2=0.342 $Y2=0.234
cc_21 N_A_c_1_p N_Y_c_42_n 0.00100412f $X=0.297 $Y=0.135 $X2=0.351 $Y2=0.126

* END of "./INVx5_ASAP7_75t_SRAM.pex.sp.INVX5_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVx6_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:35:21 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVx6_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVx6_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVx6_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:35:21 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVX6_ASAP7_75T_SRAM%A 2 7 10 15 18 23 26 31 34 39 42 45 47 59 VSS
c27 59 VSS 0.0275217f $X=0.066 $Y=0.1355
c28 45 VSS 0.0295445f $X=0.351 $Y=0.135
c29 42 VSS 0.0645347f $X=0.351 $Y=0.0675
c30 34 VSS 0.0644226f $X=0.297 $Y=0.0675
c31 26 VSS 0.0642127f $X=0.243 $Y=0.0675
c32 18 VSS 0.0642127f $X=0.189 $Y=0.0675
c33 10 VSS 0.0644226f $X=0.135 $Y=0.0675
c34 2 VSS 0.0655089f $X=0.081 $Y=0.0675
r35 56 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r36 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r37 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r38 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r39 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r40 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r41 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r42 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r43 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r44 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r45 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r46 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r47 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r48 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r49 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r50 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r51 5 56 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r52 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r53 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVX6_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 20 21 22 25 26 27 30 31 34 38
+ 41 42 56 VSS
c27 56 VSS 0.0113717f $X=0.4035 $Y=0.1475
c28 42 VSS 0.0386536f $X=0.396 $Y=0.234
c29 41 VSS 0.00929752f $X=0.324 $Y=0.036
c30 38 VSS 0.00928952f $X=0.216 $Y=0.036
c31 34 VSS 0.00904082f $X=0.108 $Y=0.036
c32 31 VSS 0.0386536f $X=0.396 $Y=0.036
c33 30 VSS 0.00929752f $X=0.324 $Y=0.2025
c34 26 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c35 25 VSS 0.00928952f $X=0.216 $Y=0.2025
c36 21 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c37 20 VSS 0.00904082f $X=0.108 $Y=0.2025
c38 16 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c39 11 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c40 6 VSS 5.38922e-19 $X=0.233 $Y=0.0675
c41 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r42 54 56 5.26235 $w=1.8e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.1475
r43 53 56 6.95988 $w=1.8e-08 $l=1.025e-07 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.1475
r44 48 51 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.324 $Y2=0.234
r45 44 48 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.216 $Y2=0.234
r46 42 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r47 42 51 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.324 $Y2=0.234
r48 40 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r49 37 40 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.324 $Y2=0.036
r50 37 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r51 33 37 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.216 $Y2=0.036
r52 33 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r53 31 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r54 31 40 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.324 $Y2=0.036
r55 30 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r56 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r57 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r58 25 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r59 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r60 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r61 20 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r62 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r63 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r64 15 41 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r65 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r66 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r67 10 38 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r68 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r69 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r70 5 34 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r71 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r72 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./INVx6_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVx6_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_A_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_A_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_A_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_A_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_A_M6_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M7 N_Y_M7_d N_A_M7_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M8 N_Y_M8_d N_A_M8_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M9 N_Y_M9_d N_A_M9_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M10 N_Y_M10_d N_A_M10_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_Y_M11_d N_A_M11_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "INVx6_ASAP7_75t_SRAM.pex.sp.INVX6_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVx6_ASAP7_75t_SRAM.pex.sp.INVX6_ASAP7_75T_SRAM.pxi"
* File: INVx6_ASAP7_75t_SRAM.pex.sp.INVX6_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:35:21 2017
* 
x_PM_INVX6_ASAP7_75T_SRAM%A N_A_M0_g N_A_M6_g N_A_M1_g N_A_M7_g N_A_M2_g N_A_M8_g
+ N_A_M3_g N_A_M9_g N_A_M4_g N_A_M10_g N_A_M5_g N_A_c_1_p N_A_M11_g A VSS
+ PM_INVX6_ASAP7_75T_SRAM%A
x_PM_INVX6_ASAP7_75T_SRAM%Y N_Y_M1_d N_Y_M0_d N_Y_M3_d N_Y_M2_d N_Y_M5_d N_Y_M4_d
+ N_Y_M7_d N_Y_M6_d N_Y_c_32_n N_Y_M9_d N_Y_M8_d N_Y_c_34_n N_Y_M11_d N_Y_M10_d
+ N_Y_c_36_n N_Y_c_37_n N_Y_c_44_n N_Y_c_45_n N_Y_c_46_n N_Y_c_47_n Y VSS
+ PM_INVX6_ASAP7_75T_SRAM%Y
cc_1 N_A_c_1_p N_Y_M1_d 3.80663e-19 $X=0.351 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_2 N_A_c_1_p N_Y_M3_d 3.80663e-19 $X=0.351 $Y=0.135 $X2=0.233 $Y2=0.0675
cc_3 N_A_c_1_p N_Y_M5_d 3.80663e-19 $X=0.351 $Y=0.135 $X2=0.341 $Y2=0.0675
cc_4 N_A_c_1_p N_Y_M7_d 3.80663e-19 $X=0.351 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_5 N_A_c_1_p N_Y_c_32_n 8.00061e-19 $X=0.351 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_6 N_A_c_1_p N_Y_M9_d 3.80663e-19 $X=0.351 $Y=0.135 $X2=0.233 $Y2=0.2025
cc_7 N_A_c_1_p N_Y_c_34_n 8.00061e-19 $X=0.351 $Y=0.135 $X2=0.216 $Y2=0.2025
cc_8 N_A_c_1_p N_Y_M11_d 3.80663e-19 $X=0.351 $Y=0.135 $X2=0.341 $Y2=0.2025
cc_9 N_A_c_1_p N_Y_c_36_n 8.00061e-19 $X=0.351 $Y=0.135 $X2=0.324 $Y2=0.2025
cc_10 N_A_M1_g N_Y_c_37_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.396 $Y2=0.036
cc_11 N_A_M2_g N_Y_c_37_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.396 $Y2=0.036
cc_12 N_A_M3_g N_Y_c_37_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.396 $Y2=0.036
cc_13 N_A_M4_g N_Y_c_37_n 4.59284e-19 $X=0.297 $Y=0.0675 $X2=0.396 $Y2=0.036
cc_14 N_A_M5_g N_Y_c_37_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.396 $Y2=0.036
cc_15 N_A_c_1_p N_Y_c_37_n 0.00327571f $X=0.351 $Y=0.135 $X2=0.396 $Y2=0.036
cc_16 A N_Y_c_37_n 5.31858e-19 $X=0.066 $Y=0.1355 $X2=0.396 $Y2=0.036
cc_17 N_A_c_1_p N_Y_c_44_n 8.00061e-19 $X=0.351 $Y=0.135 $X2=0.108 $Y2=0.036
cc_18 N_A_c_1_p N_Y_c_45_n 8.00061e-19 $X=0.351 $Y=0.135 $X2=0.216 $Y2=0.036
cc_19 N_A_c_1_p N_Y_c_46_n 8.00061e-19 $X=0.351 $Y=0.135 $X2=0.324 $Y2=0.036
cc_20 N_A_M1_g N_Y_c_47_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.396 $Y2=0.234
cc_21 N_A_M2_g N_Y_c_47_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.396 $Y2=0.234
cc_22 N_A_M3_g N_Y_c_47_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.396 $Y2=0.234
cc_23 N_A_M4_g N_Y_c_47_n 4.59284e-19 $X=0.297 $Y=0.0675 $X2=0.396 $Y2=0.234
cc_24 N_A_M5_g N_Y_c_47_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.396 $Y2=0.234
cc_25 N_A_c_1_p N_Y_c_47_n 0.00327571f $X=0.351 $Y=0.135 $X2=0.396 $Y2=0.234
cc_26 A N_Y_c_47_n 5.31858e-19 $X=0.066 $Y=0.1355 $X2=0.396 $Y2=0.234
cc_27 N_A_c_1_p Y 0.00101646f $X=0.351 $Y=0.135 $X2=0.4035 $Y2=0.1475

* END of "./INVx6_ASAP7_75t_SRAM.pex.sp.INVX6_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVx8_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:35:44 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVx8_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVx8_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVx8_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:35:44 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVX8_ASAP7_75T_SRAM%A 2 7 10 15 18 23 26 31 34 39 42 47 50 55 58 61 63
+ 71 VSS
c35 71 VSS 0.0275313f $X=0.062 $Y=0.1315
c36 61 VSS 0.0396921f $X=0.459 $Y=0.135
c37 58 VSS 0.0645347f $X=0.459 $Y=0.0675
c38 50 VSS 0.0644226f $X=0.405 $Y=0.0675
c39 42 VSS 0.0642127f $X=0.351 $Y=0.0675
c40 34 VSS 0.0642127f $X=0.297 $Y=0.0675
c41 26 VSS 0.0642127f $X=0.243 $Y=0.0675
c42 18 VSS 0.0642127f $X=0.189 $Y=0.0675
c43 10 VSS 0.0644226f $X=0.135 $Y=0.0675
c44 2 VSS 0.0655089f $X=0.081 $Y=0.0675
r45 71 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r46 61 63 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r47 58 61 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r48 53 61 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r49 53 55 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r50 50 53 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
r51 45 53 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r52 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r53 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r54 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r55 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r56 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r57 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r58 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r59 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r60 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r61 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r62 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r63 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r64 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r65 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r66 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r67 5 75 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r68 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r69 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVX8_ASAP7_75T_SRAM%Y 1 2 6 7 11 12 16 17 21 22 25 26 27 30 31 32 35 36
+ 37 40 41 44 48 51 54 55 72 VSS
c35 72 VSS 0.0113717f $X=0.513 $Y=0.1475
c36 55 VSS 0.0506904f $X=0.504 $Y=0.234
c37 54 VSS 0.00929752f $X=0.432 $Y=0.036
c38 51 VSS 0.00928953f $X=0.324 $Y=0.036
c39 48 VSS 0.00928954f $X=0.216 $Y=0.036
c40 44 VSS 0.00904082f $X=0.108 $Y=0.036
c41 41 VSS 0.0506904f $X=0.504 $Y=0.036
c42 40 VSS 0.00929752f $X=0.432 $Y=0.2025
c43 36 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c44 35 VSS 0.00928953f $X=0.324 $Y=0.2025
c45 31 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c46 30 VSS 0.00928954f $X=0.216 $Y=0.2025
c47 26 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c48 25 VSS 0.00904082f $X=0.108 $Y=0.2025
c49 21 VSS 5.72268e-19 $X=0.125 $Y=0.2025
c50 16 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c51 11 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c52 6 VSS 5.38922e-19 $X=0.233 $Y=0.0675
c53 1 VSS 5.72268e-19 $X=0.125 $Y=0.0675
r54 70 72 5.26235 $w=1.8e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.1475
r55 69 72 6.95988 $w=1.8e-08 $l=1.025e-07 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.1475
r56 64 67 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r57 61 64 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.324 $Y2=0.234
r58 57 61 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.216 $Y2=0.234
r59 55 70 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.234 $X2=0.513 $Y2=0.225
r60 55 67 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.432 $Y2=0.234
r61 53 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r62 50 53 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r63 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r64 47 50 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.324 $Y2=0.036
r65 47 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r66 43 47 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.216 $Y2=0.036
r67 43 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r68 41 69 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.036 $X2=0.513 $Y2=0.045
r69 41 53 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.432 $Y2=0.036
r70 40 67 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r71 37 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r72 36 40 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r73 35 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r74 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r75 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r76 30 61 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r77 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r78 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r79 25 57 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r80 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r81 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r82 20 54 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r83 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r84 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r85 15 51 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r86 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r87 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r88 10 48 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r89 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r90 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r91 5 44 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r92 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r93 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./INVx8_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVx8_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_A_M2_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_A_M3_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_A_M4_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_A_M5_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_A_M6_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_A_M7_g VSS VSS NMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_A_M8_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M9 N_Y_M9_d N_A_M9_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M10 N_Y_M10_d N_A_M10_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M11 N_Y_M11_d N_A_M11_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M12 N_Y_M12_d N_A_M12_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M13 N_Y_M13_d N_A_M13_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M14 N_Y_M14_d N_A_M14_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M15 N_Y_M15_d N_A_M15_g VDD VDD PMOS_SRAM L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "INVx8_ASAP7_75t_SRAM.pex.sp.INVX8_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVx8_ASAP7_75t_SRAM.pex.sp.INVX8_ASAP7_75T_SRAM.pxi"
* File: INVx8_ASAP7_75t_SRAM.pex.sp.INVX8_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:35:44 2017
* 
x_PM_INVX8_ASAP7_75T_SRAM%A N_A_M0_g N_A_M8_g N_A_M1_g N_A_M9_g N_A_M2_g N_A_M10_g
+ N_A_M3_g N_A_M11_g N_A_M4_g N_A_M12_g N_A_M5_g N_A_M13_g N_A_M6_g N_A_M14_g
+ N_A_M7_g N_A_c_1_p N_A_M15_g A VSS PM_INVX8_ASAP7_75T_SRAM%A
x_PM_INVX8_ASAP7_75T_SRAM%Y N_Y_M1_d N_Y_M0_d N_Y_M3_d N_Y_M2_d N_Y_M5_d N_Y_M4_d
+ N_Y_M7_d N_Y_M6_d N_Y_M9_d N_Y_M8_d N_Y_c_41_n N_Y_M11_d N_Y_M10_d N_Y_c_43_n
+ N_Y_M13_d N_Y_M12_d N_Y_c_45_n N_Y_M15_d N_Y_M14_d N_Y_c_47_n N_Y_c_48_n
+ N_Y_c_57_n N_Y_c_58_n N_Y_c_59_n N_Y_c_60_n N_Y_c_61_n Y VSS
+ PM_INVX8_ASAP7_75T_SRAM%Y
cc_1 N_A_c_1_p N_Y_M1_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.125 $Y2=0.0675
cc_2 N_A_c_1_p N_Y_M3_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.233 $Y2=0.0675
cc_3 N_A_c_1_p N_Y_M5_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.341 $Y2=0.0675
cc_4 N_A_c_1_p N_Y_M7_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.449 $Y2=0.0675
cc_5 N_A_c_1_p N_Y_M9_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.125 $Y2=0.2025
cc_6 N_A_c_1_p N_Y_c_41_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.108 $Y2=0.2025
cc_7 N_A_c_1_p N_Y_M11_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.233 $Y2=0.2025
cc_8 N_A_c_1_p N_Y_c_43_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.216 $Y2=0.2025
cc_9 N_A_c_1_p N_Y_M13_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.341 $Y2=0.2025
cc_10 N_A_c_1_p N_Y_c_45_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.324 $Y2=0.2025
cc_11 N_A_c_1_p N_Y_M15_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.449 $Y2=0.2025
cc_12 N_A_c_1_p N_Y_c_47_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.432 $Y2=0.2025
cc_13 N_A_M1_g N_Y_c_48_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.504 $Y2=0.036
cc_14 N_A_M2_g N_Y_c_48_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.504 $Y2=0.036
cc_15 N_A_M3_g N_Y_c_48_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.504 $Y2=0.036
cc_16 N_A_M4_g N_Y_c_48_n 4.59284e-19 $X=0.297 $Y=0.0675 $X2=0.504 $Y2=0.036
cc_17 N_A_M5_g N_Y_c_48_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.504 $Y2=0.036
cc_18 N_A_M6_g N_Y_c_48_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0.504 $Y2=0.036
cc_19 N_A_M7_g N_Y_c_48_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.504 $Y2=0.036
cc_20 N_A_c_1_p N_Y_c_48_n 0.00463796f $X=0.459 $Y=0.135 $X2=0.504 $Y2=0.036
cc_21 A N_Y_c_48_n 5.32649e-19 $X=0.062 $Y=0.1315 $X2=0.504 $Y2=0.036
cc_22 N_A_c_1_p N_Y_c_57_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.108 $Y2=0.036
cc_23 N_A_c_1_p N_Y_c_58_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.216 $Y2=0.036
cc_24 N_A_c_1_p N_Y_c_59_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.324 $Y2=0.036
cc_25 N_A_c_1_p N_Y_c_60_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.432 $Y2=0.036
cc_26 N_A_M1_g N_Y_c_61_n 4.59284e-19 $X=0.135 $Y=0.0675 $X2=0.504 $Y2=0.234
cc_27 N_A_M2_g N_Y_c_61_n 4.59284e-19 $X=0.189 $Y=0.0675 $X2=0.504 $Y2=0.234
cc_28 N_A_M3_g N_Y_c_61_n 4.59284e-19 $X=0.243 $Y=0.0675 $X2=0.504 $Y2=0.234
cc_29 N_A_M4_g N_Y_c_61_n 4.59284e-19 $X=0.297 $Y=0.0675 $X2=0.504 $Y2=0.234
cc_30 N_A_M5_g N_Y_c_61_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.504 $Y2=0.234
cc_31 N_A_M6_g N_Y_c_61_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0.504 $Y2=0.234
cc_32 N_A_M7_g N_Y_c_61_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.504 $Y2=0.234
cc_33 N_A_c_1_p N_Y_c_61_n 0.00463796f $X=0.459 $Y=0.135 $X2=0.504 $Y2=0.234
cc_34 A N_Y_c_61_n 5.32649e-19 $X=0.062 $Y=0.1315 $X2=0.504 $Y2=0.234
cc_35 N_A_c_1_p Y 0.0010177f $X=0.459 $Y=0.135 $X2=0.513 $Y2=0.1475

* END of "./INVx8_ASAP7_75t_SRAM.pex.sp.INVX8_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVxp33_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:36:06 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVxp33_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVxp33_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVxp33_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:36:06 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVXP33_ASAP7_75T_SRAM%A 2 7 13 15 18 21 VSS
c3 21 VSS 0.00752511f $X=0.018 $Y=0.135
c4 18 VSS 0.00262293f $X=0.064 $Y=0.135
c5 13 VSS 0.00685663f $X=0.018 $Y=0.144
c6 5 VSS 0.00597435f $X=0.081 $Y=0.135
c7 2 VSS 0.0702997f $X=0.081 $Y=0.0405
r8 18 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r9 16 21 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r10 16 18 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.064 $Y2=0.135
r11 13 21 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r12 13 15 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1495
r13 5 19 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r14 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2295
r15 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0405 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVXP33_ASAP7_75T_SRAM%Y 1 6 12 14 16 VSS
c3 30 VSS 0.00457827f $X=0.126 $Y=0.234
c4 29 VSS 0.00278493f $X=0.135 $Y=0.234
c5 22 VSS 0.00457655f $X=0.126 $Y=0.036
c6 21 VSS 0.00278493f $X=0.135 $Y=0.036
c7 16 VSS 7.74764e-19 $X=0.135 $Y=0.144
c8 14 VSS 0.00465839f $X=0.1355 $Y=0.1145
c9 12 VSS 0.00447748f $X=0.135 $Y=0.225
c10 9 VSS 0.00426628f $X=0.106 $Y=0.2295
c11 4 VSS 0.00426628f $X=0.106 $Y=0.0405
r12 30 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r13 29 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r14 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r15 22 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r16 21 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r17 18 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r18 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.144
r19 14 15 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.1145 $X2=0.135 $Y2=0.126
r20 12 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.234
r21 12 16 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.144
r22 11 21 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.036
r23 11 14 4.71914 $w=1.8e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.1145
r24 9 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r25 6 9 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.2295 $X2=0.106 $Y2=0.2295
r26 4 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r27 1 4 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0405 $X2=0.106 $Y2=0.0405
.ends


* END of "./INVxp33_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVxp33_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VDD VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071 $Y=0.216
*
* 
* .include "INVxp33_ASAP7_75t_SRAM.pex.sp.INVXP33_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVxp33_ASAP7_75t_SRAM.pex.sp.INVXP33_ASAP7_75T_SRAM.pxi"
* File: INVxp33_ASAP7_75t_SRAM.pex.sp.INVXP33_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:36:06 2017
* 
x_PM_INVXP33_ASAP7_75T_SRAM%A N_A_M0_g N_A_M1_g N_A_c_1_p A N_A_c_3_p N_A_c_2_p VSS
+ PM_INVXP33_ASAP7_75T_SRAM%A
x_PM_INVXP33_ASAP7_75T_SRAM%Y N_Y_M0_d N_Y_M1_d N_Y_c_4_n Y N_Y_c_6_n VSS
+ PM_INVXP33_ASAP7_75T_SRAM%Y
cc_1 N_A_c_1_p N_Y_c_4_n 0.00137512f $X=0.018 $Y=0.144 $X2=0.135 $Y2=0.225
cc_2 N_A_c_2_p Y 0.00137274f $X=0.018 $Y=0.135 $X2=0.1355 $Y2=0.1145
cc_3 N_A_c_3_p N_Y_c_6_n 5.19281e-19 $X=0.064 $Y=0.135 $X2=0.135 $Y2=0.144

* END of "./INVxp33_ASAP7_75t_SRAM.pex.sp.INVXP33_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: INVxp67_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:36:29 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "INVxp67_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./INVxp67_ASAP7_75t_SRAM.pex.sp.pex"
* File: INVxp67_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:36:29 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_INVXP67_ASAP7_75T_SRAM%A 2 7 18 20 VSS
c3 20 VSS 0.00259832f $X=0.064 $Y=0.135
c4 18 VSS 0.014046f $X=0.04 $Y=0.1375
c5 5 VSS 0.00613135f $X=0.081 $Y=0.135
c6 2 VSS 0.0702997f $X=0.081 $Y=0.054
r7 20 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r8 18 20 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.135 $X2=0.064 $Y2=0.135
r9 5 21 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r10 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r11 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_INVXP67_ASAP7_75T_SRAM%Y 1 6 12 14 16 VSS
c3 30 VSS 0.00453062f $X=0.126 $Y=0.234
c4 29 VSS 0.00278493f $X=0.135 $Y=0.234
c5 22 VSS 0.0045289f $X=0.126 $Y=0.036
c6 21 VSS 0.00278493f $X=0.135 $Y=0.036
c7 16 VSS 7.74764e-19 $X=0.135 $Y=0.144
c8 14 VSS 0.0043566f $X=0.1355 $Y=0.1145
c9 12 VSS 0.00417569f $X=0.135 $Y=0.225
c10 9 VSS 0.00549433f $X=0.106 $Y=0.216
c11 4 VSS 0.00549433f $X=0.106 $Y=0.054
r12 30 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r13 29 31 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r14 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r15 22 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r16 21 23 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r17 18 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r18 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.144
r19 14 15 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.1145 $X2=0.135 $Y2=0.126
r20 12 29 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.234
r21 12 16 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.144
r22 11 21 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.036
r23 11 14 4.71914 $w=1.8e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.1145
r24 9 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r25 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.216 $X2=0.106 $Y2=0.216
r26 4 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r27 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.054 $X2=0.106 $Y2=0.054
.ends


* END of "./INVxp67_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt INVxp67_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
*
* 
* .include "INVxp67_ASAP7_75t_SRAM.pex.sp.INVXP67_ASAP7_75T_SRAM.pxi"
* BEGIN of "./INVxp67_ASAP7_75t_SRAM.pex.sp.INVXP67_ASAP7_75T_SRAM.pxi"
* File: INVxp67_ASAP7_75t_SRAM.pex.sp.INVXP67_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:36:29 2017
* 
x_PM_INVXP67_ASAP7_75T_SRAM%A N_A_M0_g N_A_M1_g A N_A_c_3_p VSS
+ PM_INVXP67_ASAP7_75T_SRAM%A
x_PM_INVXP67_ASAP7_75T_SRAM%Y N_Y_M0_d N_Y_M1_d N_Y_c_4_n Y N_Y_c_6_n VSS
+ PM_INVXP67_ASAP7_75T_SRAM%Y
cc_1 A N_Y_c_4_n 0.00102711f $X=0.04 $Y=0.1375 $X2=0.135 $Y2=0.225
cc_2 A Y 0.00102556f $X=0.04 $Y=0.1375 $X2=0.1355 $Y2=0.1145
cc_3 N_A_c_3_p N_Y_c_6_n 5.19281e-19 $X=0.064 $Y=0.135 $X2=0.135 $Y2=0.144

* END of "./INVxp67_ASAP7_75t_SRAM.pex.sp.INVXP67_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: HB1xp67_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:30:07 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "HB1xp67_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./HB1xp67_ASAP7_75t_SRAM.pex.sp.pex"
* File: HB1xp67_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:30:07 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_HB1XP67_ASAP7_75T_SRAM%A 2 5 7 16 21 28 VSS
c14 28 VSS 0.00623497f $X=0.018 $Y=0.135
c15 24 VSS 5.0748e-19 $X=0.055 $Y=0.135
c16 23 VSS 0.00109101f $X=0.046 $Y=0.135
c17 21 VSS 4.75057e-19 $X=0.064 $Y=0.135
c18 16 VSS 0.00553592f $X=0.019 $Y=0.1495
c19 5 VSS 0.0045218f $X=0.081 $Y=0.135
c20 2 VSS 0.0663428f $X=0.081 $Y=0.0405
r21 23 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.055 $Y2=0.135
r22 21 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.064
+ $Y=0.135 $X2=0.055 $Y2=0.135
r23 21 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r24 19 28 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r25 19 23 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.046 $Y2=0.135
r26 13 28 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r27 13 16 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1495
r28 5 22 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r29 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2295
r30 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0405 $X2=0.081 $Y2=0.135
.ends

.subckt PM_HB1XP67_ASAP7_75T_SRAM%4 2 5 7 9 14 19 21 26 27 28 30 35 36 38 39 40 43
+ 44 48 51 56 63 VSS
c23 64 VSS 3.34713e-19 $X=0.126 $Y=0.162
c24 63 VSS 3.75831e-19 $X=0.117 $Y=0.162
c25 62 VSS 4.939e-19 $X=0.135 $Y=0.162
c26 58 VSS 3.34713e-19 $X=0.126 $Y=0.108
c27 57 VSS 3.75831e-19 $X=0.117 $Y=0.108
c28 56 VSS 4.939e-19 $X=0.135 $Y=0.108
c29 53 VSS 1.53902e-19 $X=0.135 $Y=0.1485
c30 51 VSS 5.41721e-21 $X=0.135 $Y=0.1305
c31 50 VSS 3.03024e-19 $X=0.135 $Y=0.126
c32 48 VSS 5.41721e-21 $X=0.135 $Y=0.135
c33 46 VSS 3.77561e-20 $X=0.135 $Y=0.153
c34 44 VSS 0.00179951f $X=0.108 $Y=0.207
c35 43 VSS 4.31818e-19 $X=0.108 $Y=0.189
c36 42 VSS 0.00119316f $X=0.108 $Y=0.225
c37 40 VSS 0.00179951f $X=0.108 $Y=0.081
c38 39 VSS 0.00119316f $X=0.108 $Y=0.063
c39 38 VSS 4.31818e-19 $X=0.108 $Y=0.099
c40 36 VSS 9.17922e-19 $X=0.0885 $Y=0.234
c41 35 VSS 0.00257781f $X=0.078 $Y=0.234
c42 30 VSS 0.00219602f $X=0.054 $Y=0.234
c43 28 VSS 0.00489465f $X=0.099 $Y=0.234
c44 27 VSS 9.17922e-19 $X=0.0885 $Y=0.036
c45 26 VSS 0.00257781f $X=0.078 $Y=0.036
c46 21 VSS 0.00219602f $X=0.054 $Y=0.036
c47 19 VSS 0.00489465f $X=0.099 $Y=0.036
c48 17 VSS 0.00435822f $X=0.056 $Y=0.2295
c49 14 VSS 2.67274e-19 $X=0.071 $Y=0.2295
c50 12 VSS 0.00435822f $X=0.056 $Y=0.0405
c51 9 VSS 2.67274e-19 $X=0.071 $Y=0.0405
c52 5 VSS 0.00185592f $X=0.135 $Y=0.135
c53 2 VSS 0.0661191f $X=0.135 $Y=0.054
r54 63 64 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.162 $X2=0.126 $Y2=0.162
r55 62 64 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.162 $X2=0.126 $Y2=0.162
r56 60 63 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.162 $X2=0.117 $Y2=0.162
r57 57 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.108 $X2=0.126 $Y2=0.108
r58 56 58 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.108 $X2=0.126 $Y2=0.108
r59 54 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.108 $X2=0.117 $Y2=0.108
r60 52 53 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.1485
r61 50 51 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.1305
r62 48 52 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r63 48 51 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.1305
r64 46 62 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.153 $X2=0.135 $Y2=0.162
r65 46 53 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.153 $X2=0.135 $Y2=0.1485
r66 45 56 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.117 $X2=0.135 $Y2=0.108
r67 45 50 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.117 $X2=0.135 $Y2=0.126
r68 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.189 $X2=0.108 $Y2=0.207
r69 42 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.225 $X2=0.108 $Y2=0.207
r70 41 60 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.171 $X2=0.108 $Y2=0.162
r71 41 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.171 $X2=0.108 $Y2=0.189
r72 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.063 $X2=0.108 $Y2=0.081
r73 38 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.099 $X2=0.108 $Y2=0.108
r74 38 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.099 $X2=0.108 $Y2=0.081
r75 37 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.045 $X2=0.108 $Y2=0.063
r76 35 36 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.234 $X2=0.0885 $Y2=0.234
r77 30 35 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.078 $Y2=0.234
r78 28 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.099 $Y=0.234 $X2=0.108 $Y2=0.225
r79 28 36 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.234 $X2=0.0885 $Y2=0.234
r80 26 27 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.036 $X2=0.0885 $Y2=0.036
r81 21 26 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.078 $Y2=0.036
r82 19 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.099 $Y=0.036 $X2=0.108 $Y2=0.045
r83 19 27 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.036 $X2=0.0885 $Y2=0.036
r84 17 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r85 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2295 $X2=0.056 $Y2=0.2295
r86 12 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r87 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0405 $X2=0.056 $Y2=0.0405
r88 5 48 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r89 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r90 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_HB1XP67_ASAP7_75T_SRAM%Y 1 4 6 9 12 14 15 16 18 24 32 VSS
c9 32 VSS 0.00407364f $X=0.18 $Y=0.234
c10 31 VSS 0.00278493f $X=0.189 $Y=0.234
c11 24 VSS 0.00407364f $X=0.18 $Y=0.036
c12 23 VSS 0.00278493f $X=0.189 $Y=0.036
c13 18 VSS 0.00128813f $X=0.189 $Y=0.198
c14 16 VSS 0.00122153f $X=0.189 $Y=0.12425
c15 15 VSS 0.00263333f $X=0.189 $Y=0.099
c16 14 VSS 0.00208512f $X=0.19 $Y=0.1495
c17 12 VSS 0.00134931f $X=0.189 $Y=0.225
c18 9 VSS 0.00562876f $X=0.16 $Y=0.216
c19 4 VSS 0.00562876f $X=0.16 $Y=0.054
r20 32 33 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r21 31 33 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.1845 $Y2=0.234
r22 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r23 24 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r24 23 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.036 $X2=0.1845 $Y2=0.036
r25 20 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r26 17 18 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.171 $X2=0.189 $Y2=0.198
r27 15 16 1.71451 $w=1.8e-08 $l=2.525e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.099 $X2=0.189 $Y2=0.12425
r28 14 17 1.45988 $w=1.8e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.1495 $X2=0.189 $Y2=0.171
r29 14 16 1.71451 $w=1.8e-08 $l=2.525e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.1495 $X2=0.189 $Y2=0.12425
r30 12 31 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.234
r31 12 18 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.198
r32 11 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.036
r33 11 15 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.099
r34 9 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r35 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.216 $X2=0.16 $Y2=0.216
r36 4 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r37 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.054 $X2=0.16 $Y2=0.054
.ends


* END of "./HB1xp67_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt HB1xp67_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 VSS N_A_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_4_M1_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VDD N_A_M2_g N_4_M2_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071 $Y=0.216
M3 N_Y_M3_d N_4_M3_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
*
* 
* .include "HB1xp67_ASAP7_75t_SRAM.pex.sp.HB1XP67_ASAP7_75T_SRAM.pxi"
* BEGIN of "./HB1xp67_ASAP7_75t_SRAM.pex.sp.HB1XP67_ASAP7_75T_SRAM.pxi"
* File: HB1xp67_ASAP7_75t_SRAM.pex.sp.HB1XP67_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:30:07 2017
* 
x_PM_HB1XP67_ASAP7_75T_SRAM%A N_A_M0_g N_A_c_2_p N_A_M2_g A N_A_c_13_p N_A_c_3_p
+ VSS PM_HB1XP67_ASAP7_75T_SRAM%A
x_PM_HB1XP67_ASAP7_75T_SRAM%4 N_4_M1_g N_4_c_16_n N_4_M3_g N_4_M0_s N_4_M2_s
+ N_4_c_36_p N_4_c_17_n N_4_c_18_n N_4_c_19_n N_4_c_37_p N_4_c_20_n N_4_c_21_n
+ N_4_c_22_n N_4_c_23_n N_4_c_29_p N_4_c_24_n N_4_c_25_n N_4_c_26_n N_4_c_32_p
+ N_4_c_27_n N_4_c_34_p N_4_c_28_n VSS PM_HB1XP67_ASAP7_75T_SRAM%4
x_PM_HB1XP67_ASAP7_75T_SRAM%Y N_Y_M1_d N_Y_c_38_n N_Y_M3_d N_Y_c_39_n N_Y_c_40_n Y
+ N_Y_c_42_n N_Y_c_43_n N_Y_c_44_n N_Y_c_45_n N_Y_c_46_n VSS
+ PM_HB1XP67_ASAP7_75T_SRAM%Y
cc_1 N_A_M0_g N_4_M1_g 0.00287079f $X=0.081 $Y=0.0405 $X2=0.135 $Y2=0.054
cc_2 N_A_c_2_p N_4_c_16_n 0.0011f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A_c_3_p N_4_c_17_n 5.65154e-19 $X=0.018 $Y=0.135 $X2=0.054 $Y2=0.036
cc_4 N_A_c_2_p N_4_c_18_n 2.28446e-19 $X=0.081 $Y=0.135 $X2=0.078 $Y2=0.036
cc_5 N_A_M0_g N_4_c_19_n 2.41124e-19 $X=0.081 $Y=0.0405 $X2=0.0885 $Y2=0.036
cc_6 A N_4_c_20_n 5.65154e-19 $X=0.019 $Y=0.1495 $X2=0.054 $Y2=0.234
cc_7 N_A_c_2_p N_4_c_21_n 2.28446e-19 $X=0.081 $Y=0.135 $X2=0.078 $Y2=0.234
cc_8 N_A_M0_g N_4_c_22_n 2.41124e-19 $X=0.081 $Y=0.0405 $X2=0.0885 $Y2=0.234
cc_9 N_A_c_3_p N_4_c_23_n 0.00102037f $X=0.018 $Y=0.135 $X2=0.108 $Y2=0.099
cc_10 N_A_c_3_p N_4_c_24_n 5.34348e-19 $X=0.018 $Y=0.135 $X2=0.108 $Y2=0.081
cc_11 A N_4_c_25_n 5.13477e-19 $X=0.019 $Y=0.1495 $X2=0.108 $Y2=0.189
cc_12 A N_4_c_26_n 5.34348e-19 $X=0.019 $Y=0.1495 $X2=0.108 $Y2=0.207
cc_13 N_A_c_13_p N_4_c_27_n 4.18081e-19 $X=0.064 $Y=0.135 $X2=0.135 $Y2=0.1305
cc_14 A N_4_c_28_n 5.13477e-19 $X=0.019 $Y=0.1495 $X2=0.117 $Y2=0.162
cc_15 N_4_c_29_p N_Y_c_38_n 2.54174e-19 $X=0.108 $Y=0.063 $X2=0.081 $Y2=0.135
cc_16 N_4_c_26_n N_Y_c_39_n 2.54174e-19 $X=0.108 $Y=0.207 $X2=0 $Y2=0
cc_17 N_4_c_26_n N_Y_c_40_n 5.20276e-19 $X=0.108 $Y=0.207 $X2=0 $Y2=0
cc_18 N_4_c_32_p Y 0.00182786f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_19 N_4_c_29_p N_Y_c_42_n 0.00103841f $X=0.108 $Y=0.063 $X2=0.018 $Y2=0.1495
cc_20 N_4_c_34_p N_Y_c_43_n 0.00182786f $X=0.135 $Y=0.108 $X2=0.019 $Y2=0.1495
cc_21 N_4_c_25_n N_Y_c_44_n 5.20276e-19 $X=0.108 $Y=0.189 $X2=0 $Y2=0
cc_22 N_4_c_36_p N_Y_c_45_n 8.87733e-19 $X=0.099 $Y=0.036 $X2=0.055 $Y2=0.135
cc_23 N_4_c_37_p N_Y_c_46_n 8.87733e-19 $X=0.099 $Y=0.234 $X2=0 $Y2=0

* END of "./HB1xp67_ASAP7_75t_SRAM.pex.sp.HB1XP67_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: HB2xp67_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:30:30 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "HB2xp67_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./HB2xp67_ASAP7_75t_SRAM.pex.sp.pex"
* File: HB2xp67_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:30:30 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_HB2XP67_ASAP7_75T_SRAM%A 2 7 10 13 15 22 25 27 28 32 VSS
c30 32 VSS 0.00632726f $X=0.018 $Y=0.135
c31 28 VSS 3.72004e-19 $X=0.0635 $Y=0.135
c32 27 VSS 7.68869e-19 $X=0.046 $Y=0.135
c33 25 VSS 1.82386e-19 $X=0.081 $Y=0.135
c34 22 VSS 0.00561056f $X=0.021 $Y=0.1495
c35 13 VSS 0.00566049f $X=0.135 $Y=0.135
c36 10 VSS 0.0597072f $X=0.135 $Y=0.0405
c37 2 VSS 0.0659264f $X=0.081 $Y=0.0405
r38 27 28 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r39 25 28 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r40 23 32 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r41 23 27 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.046 $Y2=0.135
r42 19 32 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r43 19 22 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1495
r44 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2295
r45 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0405 $X2=0.135 $Y2=0.135
r46 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r47 5 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r48 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2295
r49 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0405 $X2=0.081 $Y2=0.135
.ends

.subckt PM_HB2XP67_ASAP7_75T_SRAM%4 2 5 7 9 14 19 21 26 28 30 35 38 39 40 43 44 47
+ 51 VSS
c36 47 VSS 0.00297943f $X=0.189 $Y=0.135
c37 44 VSS 3.34321e-19 $X=0.135 $Y=0.207
c38 43 VSS 5.00212e-19 $X=0.135 $Y=0.189
c39 42 VSS 6.9932e-19 $X=0.135 $Y=0.225
c40 40 VSS 3.34321e-19 $X=0.135 $Y=0.081
c41 39 VSS 6.9932e-19 $X=0.135 $Y=0.063
c42 38 VSS 5.00212e-19 $X=0.135 $Y=0.126
c43 36 VSS 0.00154104f $X=0.1105 $Y=0.234
c44 35 VSS 0.00363755f $X=0.095 $Y=0.234
c45 30 VSS 0.00186632f $X=0.054 $Y=0.234
c46 28 VSS 0.00445717f $X=0.126 $Y=0.234
c47 27 VSS 0.00154104f $X=0.1105 $Y=0.036
c48 26 VSS 0.00363755f $X=0.095 $Y=0.036
c49 21 VSS 0.00186632f $X=0.054 $Y=0.036
c50 19 VSS 0.00445717f $X=0.126 $Y=0.036
c51 17 VSS 0.00302864f $X=0.056 $Y=0.2295
c52 14 VSS 2.67274e-19 $X=0.071 $Y=0.2295
c53 12 VSS 0.00302864f $X=0.056 $Y=0.0405
c54 9 VSS 2.67274e-19 $X=0.071 $Y=0.0405
c55 5 VSS 0.00242288f $X=0.189 $Y=0.135
c56 2 VSS 0.0634914f $X=0.189 $Y=0.054
r57 45 51 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.135 $Y2=0.135
r58 45 47 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.189 $Y2=0.135
r59 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.135 $Y2=0.207
r60 42 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.207
r61 41 51 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.135
r62 41 43 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.189
r63 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.063 $X2=0.135 $Y2=0.081
r64 38 51 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.135
r65 38 40 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.081
r66 37 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.063
r67 35 36 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.234 $X2=0.1105 $Y2=0.234
r68 30 35 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.095 $Y2=0.234
r69 28 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.126 $Y=0.234 $X2=0.135 $Y2=0.225
r70 28 36 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1105 $Y2=0.234
r71 26 27 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.036 $X2=0.1105 $Y2=0.036
r72 21 26 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.095 $Y2=0.036
r73 19 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.126 $Y=0.036 $X2=0.135 $Y2=0.045
r74 19 27 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.1105 $Y2=0.036
r75 17 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r76 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2295 $X2=0.056 $Y2=0.2295
r77 12 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r78 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0405 $X2=0.056 $Y2=0.0405
r79 5 47 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r80 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r81 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_HB2XP67_ASAP7_75T_SRAM%Y 1 6 12 14 15 16 18 28 VSS
c6 34 VSS 0.00270568f $X=0.234 $Y=0.234
c7 33 VSS 0.00278493f $X=0.243 $Y=0.234
c8 28 VSS 0.00142361f $X=0.216 $Y=0.234
c9 24 VSS 0.00270568f $X=0.234 $Y=0.036
c10 23 VSS 0.00278493f $X=0.243 $Y=0.036
c11 18 VSS 0.00142361f $X=0.216 $Y=0.036
c12 16 VSS 7.46953e-19 $X=0.243 $Y=0.144
c13 15 VSS 0.00420929f $X=0.243 $Y=0.126
c14 12 VSS 0.00420929f $X=0.243 $Y=0.225
c15 9 VSS 0.00547789f $X=0.214 $Y=0.216
c16 4 VSS 0.00547789f $X=0.214 $Y=0.054
r17 34 35 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.2385 $Y2=0.234
r18 33 35 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.234 $X2=0.2385 $Y2=0.234
r19 28 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.234 $Y2=0.234
r20 24 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.2385 $Y2=0.036
r21 23 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.036 $X2=0.2385 $Y2=0.036
r22 18 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.234 $Y2=0.036
r23 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.144
r24 14 16 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.1495 $X2=0.243 $Y2=0.144
r25 12 33 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.234
r26 12 14 5.12654 $w=1.8e-08 $l=7.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.225 $X2=0.243 $Y2=0.1495
r27 11 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.036
r28 11 15 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.126
r29 9 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r30 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.216 $X2=0.214 $Y2=0.216
r31 4 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r32 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.054 $X2=0.214 $Y2=0.054
.ends

.subckt PM_HB2XP67_ASAP7_75T_SRAM%6 1 2 VSS
c0 1 VSS 0.00190998f $X=0.125 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0405 $X2=0.091 $Y2=0.0405
.ends

.subckt PM_HB2XP67_ASAP7_75T_SRAM%7 1 2 VSS
c0 1 VSS 0.00190998f $X=0.125 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2295 $X2=0.091 $Y2=0.2295
.ends


* END of "./HB2xp67_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt HB2xp67_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_6_M0_d N_A_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071
+ $Y=0.027
M1 VSS N_A_M1_g N_6_M1_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_4_M2_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 N_7_M3_d N_A_M3_g N_4_M3_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071
+ $Y=0.216
M4 VDD N_A_M4_g N_7_M4_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.125 $Y=0.216
M5 N_Y_M5_d N_4_M5_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.189
*
* 
* .include "HB2xp67_ASAP7_75t_SRAM.pex.sp.HB2XP67_ASAP7_75T_SRAM.pxi"
* BEGIN of "./HB2xp67_ASAP7_75t_SRAM.pex.sp.HB2XP67_ASAP7_75T_SRAM.pxi"
* File: HB2xp67_ASAP7_75t_SRAM.pex.sp.HB2XP67_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:30:30 2017
* 
x_PM_HB2XP67_ASAP7_75T_SRAM%A N_A_M0_g N_A_M3_g N_A_M1_g N_A_c_3_p N_A_M4_g A
+ N_A_c_10_p N_A_c_5_p N_A_c_6_p N_A_c_7_p VSS PM_HB2XP67_ASAP7_75T_SRAM%A
x_PM_HB2XP67_ASAP7_75T_SRAM%4 N_4_M2_g N_4_c_33_n N_4_M5_g N_4_M0_s N_4_M3_s
+ N_4_c_34_n N_4_c_35_n N_4_c_38_n N_4_c_41_n N_4_c_42_n N_4_c_45_n N_4_c_48_n
+ N_4_c_62_p N_4_c_51_n N_4_c_53_n N_4_c_56_n N_4_c_58_n N_4_c_59_n VSS
+ PM_HB2XP67_ASAP7_75T_SRAM%4
x_PM_HB2XP67_ASAP7_75T_SRAM%Y N_Y_M2_d N_Y_M5_d N_Y_c_67_n Y N_Y_c_68_n N_Y_c_69_n
+ N_Y_c_71_n N_Y_c_72_n VSS PM_HB2XP67_ASAP7_75T_SRAM%Y
x_PM_HB2XP67_ASAP7_75T_SRAM%6 N_6_M1_s N_6_M0_d VSS PM_HB2XP67_ASAP7_75T_SRAM%6
x_PM_HB2XP67_ASAP7_75T_SRAM%7 N_7_M4_s N_7_M3_d VSS PM_HB2XP67_ASAP7_75T_SRAM%7
cc_1 N_A_M0_g N_4_M2_g 2.13359e-19 $X=0.081 $Y=0.0405 $X2=0.189 $Y2=0.054
cc_2 N_A_M1_g N_4_M2_g 0.00268443f $X=0.135 $Y=0.0405 $X2=0.189 $Y2=0.054
cc_3 N_A_c_3_p N_4_c_33_n 0.00146414f $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_4 N_A_M1_g N_4_c_34_n 2.0666e-19 $X=0.135 $Y=0.0405 $X2=0.126 $Y2=0.036
cc_5 N_A_c_5_p N_4_c_35_n 3.03951e-19 $X=0.046 $Y=0.135 $X2=0.054 $Y2=0.036
cc_6 N_A_c_6_p N_4_c_35_n 3.03951e-19 $X=0.0635 $Y=0.135 $X2=0.054 $Y2=0.036
cc_7 N_A_c_7_p N_4_c_35_n 5.65154e-19 $X=0.018 $Y=0.135 $X2=0.054 $Y2=0.036
cc_8 N_A_M0_g N_4_c_38_n 4.28653e-19 $X=0.081 $Y=0.0405 $X2=0.095 $Y2=0.036
cc_9 N_A_c_3_p N_4_c_38_n 5.79344e-19 $X=0.135 $Y=0.135 $X2=0.095 $Y2=0.036
cc_10 N_A_c_10_p N_4_c_38_n 3.03951e-19 $X=0.081 $Y=0.135 $X2=0.095 $Y2=0.036
cc_11 N_A_M1_g N_4_c_41_n 2.0666e-19 $X=0.135 $Y=0.0405 $X2=0.126 $Y2=0.234
cc_12 A N_4_c_42_n 5.65154e-19 $X=0.021 $Y=0.1495 $X2=0.054 $Y2=0.234
cc_13 N_A_c_5_p N_4_c_42_n 3.03951e-19 $X=0.046 $Y=0.135 $X2=0.054 $Y2=0.234
cc_14 N_A_c_6_p N_4_c_42_n 3.03951e-19 $X=0.0635 $Y=0.135 $X2=0.054 $Y2=0.234
cc_15 N_A_M0_g N_4_c_45_n 4.28653e-19 $X=0.081 $Y=0.0405 $X2=0.095 $Y2=0.234
cc_16 N_A_c_3_p N_4_c_45_n 5.79344e-19 $X=0.135 $Y=0.135 $X2=0.095 $Y2=0.234
cc_17 N_A_c_10_p N_4_c_45_n 3.03951e-19 $X=0.081 $Y=0.135 $X2=0.095 $Y2=0.234
cc_18 N_A_M1_g N_4_c_48_n 6.5784e-19 $X=0.135 $Y=0.0405 $X2=0.135 $Y2=0.126
cc_19 N_A_c_3_p N_4_c_48_n 4.98151e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.126
cc_20 N_A_c_7_p N_4_c_48_n 8.16844e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.126
cc_21 N_A_M1_g N_4_c_51_n 2.9698e-19 $X=0.135 $Y=0.0405 $X2=0.135 $Y2=0.081
cc_22 N_A_c_7_p N_4_c_51_n 4.46275e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.081
cc_23 N_A_M1_g N_4_c_53_n 6.5784e-19 $X=0.135 $Y=0.0405 $X2=0.135 $Y2=0.189
cc_24 N_A_c_3_p N_4_c_53_n 4.98151e-19 $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.189
cc_25 A N_4_c_53_n 8.16844e-19 $X=0.021 $Y=0.1495 $X2=0.135 $Y2=0.189
cc_26 N_A_M1_g N_4_c_56_n 2.9698e-19 $X=0.135 $Y=0.0405 $X2=0.135 $Y2=0.207
cc_27 A N_4_c_56_n 4.46275e-19 $X=0.021 $Y=0.1495 $X2=0.135 $Y2=0.207
cc_28 N_A_c_3_p N_4_c_58_n 5.49466e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_29 N_A_c_3_p N_4_c_59_n 0.00101917f $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.135
cc_30 N_A_c_10_p N_4_c_59_n 9.16541e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_31 N_4_c_53_n N_Y_c_67_n 0.00116014f $X=0.135 $Y=0.189 $X2=0.135 $Y2=0.135
cc_32 N_4_c_62_p N_Y_c_68_n 0.00116014f $X=0.135 $Y=0.063 $X2=0.135 $Y2=0.2295
cc_33 N_4_c_33_n N_Y_c_69_n 3.15821e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_34 N_4_c_58_n N_Y_c_69_n 0.00102675f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_35 N_4_c_34_n N_Y_c_71_n 3.74279e-19 $X=0.126 $Y=0.036 $X2=0 $Y2=0
cc_36 N_4_c_41_n N_Y_c_72_n 3.74279e-19 $X=0.126 $Y=0.234 $X2=0.0635 $Y2=0.135

* END of "./HB2xp67_ASAP7_75t_SRAM.pex.sp.HB2XP67_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: HB3xp67_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:30:52 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "HB3xp67_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./HB3xp67_ASAP7_75t_SRAM.pex.sp.pex"
* File: HB3xp67_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:30:52 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_HB3XP67_ASAP7_75T_SRAM%A 2 7 10 15 18 21 23 30 33 35 36 40 VSS
c34 40 VSS 0.00666046f $X=0.018 $Y=0.135
c35 36 VSS 3.72004e-19 $X=0.0635 $Y=0.135
c36 35 VSS 7.68869e-19 $X=0.046 $Y=0.135
c37 33 VSS 1.33597e-19 $X=0.081 $Y=0.135
c38 30 VSS 0.00594377f $X=0.02 $Y=0.1585
c39 21 VSS 0.00842093f $X=0.189 $Y=0.135
c40 18 VSS 0.0622999f $X=0.189 $Y=0.0405
c41 10 VSS 0.065668f $X=0.135 $Y=0.0405
c42 2 VSS 0.0689204f $X=0.081 $Y=0.0405
r43 35 36 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r44 33 36 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r45 31 40 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r46 31 35 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.046 $Y2=0.135
r47 27 40 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r48 27 30 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1585
r49 21 23 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2295
r50 18 21 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0405 $X2=0.189 $Y2=0.135
r51 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r52 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2295
r53 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0405 $X2=0.135 $Y2=0.135
r54 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r55 5 33 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r56 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2295
r57 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0405 $X2=0.081 $Y2=0.135
.ends

.subckt PM_HB3XP67_ASAP7_75T_SRAM%4 2 5 7 9 14 19 21 26 27 28 30 35 36 38 39 40 43
+ 44 47 51 VSS
c40 47 VSS 0.00297943f $X=0.243 $Y=0.135
c41 44 VSS 3.85561e-19 $X=0.189 $Y=0.207
c42 43 VSS 6.55088e-19 $X=0.189 $Y=0.189
c43 42 VSS 4.4335e-19 $X=0.189 $Y=0.225
c44 40 VSS 3.85561e-19 $X=0.189 $Y=0.081
c45 39 VSS 4.4335e-19 $X=0.189 $Y=0.063
c46 38 VSS 6.55088e-19 $X=0.189 $Y=0.126
c47 36 VSS 0.00408275f $X=0.1375 $Y=0.234
c48 35 VSS 0.00363755f $X=0.095 $Y=0.234
c49 30 VSS 0.00188634f $X=0.054 $Y=0.234
c50 28 VSS 0.00654982f $X=0.18 $Y=0.234
c51 27 VSS 0.00408275f $X=0.1375 $Y=0.036
c52 26 VSS 0.00363755f $X=0.095 $Y=0.036
c53 21 VSS 0.00188634f $X=0.054 $Y=0.036
c54 19 VSS 0.00654982f $X=0.18 $Y=0.036
c55 17 VSS 0.00231457f $X=0.056 $Y=0.2295
c56 14 VSS 2.67274e-19 $X=0.071 $Y=0.2295
c57 12 VSS 0.00231457f $X=0.056 $Y=0.0405
c58 9 VSS 2.67274e-19 $X=0.071 $Y=0.0405
c59 5 VSS 0.00237409f $X=0.243 $Y=0.135
c60 2 VSS 0.0664863f $X=0.243 $Y=0.054
r61 45 51 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.135 $X2=0.189 $Y2=0.135
r62 45 47 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.135 $X2=0.243 $Y2=0.135
r63 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.207
r64 42 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.207
r65 41 51 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.135
r66 41 43 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.189
r67 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.063 $X2=0.189 $Y2=0.081
r68 38 51 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.135
r69 38 40 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.081
r70 37 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r71 35 36 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.234 $X2=0.1375 $Y2=0.234
r72 30 35 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.095 $Y2=0.234
r73 28 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.234 $X2=0.189 $Y2=0.225
r74 28 36 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1375 $Y2=0.234
r75 26 27 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.036 $X2=0.1375 $Y2=0.036
r76 21 26 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.095 $Y2=0.036
r77 19 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r78 19 27 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1375 $Y2=0.036
r79 17 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r80 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2295 $X2=0.056 $Y2=0.2295
r81 12 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r82 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0405 $X2=0.056 $Y2=0.0405
r83 5 47 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r84 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r85 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_HB3XP67_ASAP7_75T_SRAM%Y 1 6 12 14 15 16 18 28 VSS
c6 34 VSS 0.00270568f $X=0.288 $Y=0.234
c7 33 VSS 0.00278493f $X=0.297 $Y=0.234
c8 28 VSS 0.00142361f $X=0.27 $Y=0.234
c9 24 VSS 0.00270568f $X=0.288 $Y=0.036
c10 23 VSS 0.00278493f $X=0.297 $Y=0.036
c11 18 VSS 0.00142361f $X=0.27 $Y=0.036
c12 16 VSS 7.46953e-19 $X=0.297 $Y=0.144
c13 15 VSS 0.00420929f $X=0.297 $Y=0.126
c14 12 VSS 0.00420929f $X=0.297 $Y=0.225
c15 9 VSS 0.00547789f $X=0.268 $Y=0.216
c16 4 VSS 0.00547789f $X=0.268 $Y=0.054
r17 34 35 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.2925 $Y2=0.234
r18 33 35 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.234 $X2=0.2925 $Y2=0.234
r19 28 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.288 $Y2=0.234
r20 24 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.2925 $Y2=0.036
r21 23 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.036 $X2=0.2925 $Y2=0.036
r22 18 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.288 $Y2=0.036
r23 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.144
r24 14 16 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1585 $X2=0.297 $Y2=0.144
r25 12 33 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.234
r26 12 14 4.51543 $w=1.8e-08 $l=6.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.1585
r27 11 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.036
r28 11 15 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.126
r29 9 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r30 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.216 $X2=0.268 $Y2=0.216
r31 4 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r32 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.054 $X2=0.268 $Y2=0.054
.ends

.subckt PM_HB3XP67_ASAP7_75T_SRAM%6 1 2 VSS
c0 1 VSS 0.00192428f $X=0.125 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0405 $X2=0.091 $Y2=0.0405
.ends

.subckt PM_HB3XP67_ASAP7_75T_SRAM%7 1 2 VSS
c0 1 VSS 0.00194494f $X=0.179 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0405 $X2=0.145 $Y2=0.0405
.ends

.subckt PM_HB3XP67_ASAP7_75T_SRAM%8 1 2 VSS
c0 1 VSS 0.00192428f $X=0.125 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2295 $X2=0.091 $Y2=0.2295
.ends

.subckt PM_HB3XP67_ASAP7_75T_SRAM%9 1 2 VSS
c0 1 VSS 0.00194494f $X=0.179 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2295 $X2=0.145 $Y2=0.2295
.ends


* END of "./HB3xp67_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt HB3xp67_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_6_M0_d N_A_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071
+ $Y=0.027
M1 N_7_M1_d N_A_M1_g N_6_M1_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.125
+ $Y=0.027
M2 VSS N_A_M2_g N_7_M2_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_4_M3_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 N_8_M4_d N_A_M4_g N_4_M4_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071
+ $Y=0.216
M5 N_9_M5_d N_A_M5_g N_8_M5_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.125
+ $Y=0.216
M6 VDD N_A_M6_g N_9_M6_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.179 $Y=0.216
M7 N_Y_M7_d N_4_M7_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.189
*
* 
* .include "HB3xp67_ASAP7_75t_SRAM.pex.sp.HB3XP67_ASAP7_75T_SRAM.pxi"
* BEGIN of "./HB3xp67_ASAP7_75t_SRAM.pex.sp.HB3XP67_ASAP7_75T_SRAM.pxi"
* File: HB3xp67_ASAP7_75t_SRAM.pex.sp.HB3XP67_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:30:52 2017
* 
x_PM_HB3XP67_ASAP7_75T_SRAM%A N_A_M0_g N_A_M4_g N_A_M1_g N_A_M5_g N_A_M2_g
+ N_A_c_3_p N_A_M6_g A N_A_c_11_p N_A_c_6_p N_A_c_7_p N_A_c_8_p VSS
+ PM_HB3XP67_ASAP7_75T_SRAM%A
x_PM_HB3XP67_ASAP7_75T_SRAM%4 N_4_M3_g N_4_c_37_n N_4_M7_g N_4_M0_s N_4_M4_s
+ N_4_c_38_n N_4_c_40_n N_4_c_43_n N_4_c_46_n N_4_c_47_n N_4_c_49_n N_4_c_52_n
+ N_4_c_55_n N_4_c_56_n N_4_c_70_p N_4_c_59_n N_4_c_61_n N_4_c_64_n N_4_c_66_n
+ N_4_c_67_n VSS PM_HB3XP67_ASAP7_75T_SRAM%4
x_PM_HB3XP67_ASAP7_75T_SRAM%Y N_Y_M3_d N_Y_M7_d N_Y_c_75_n Y N_Y_c_76_n N_Y_c_77_n
+ N_Y_c_79_n N_Y_c_80_n VSS PM_HB3XP67_ASAP7_75T_SRAM%Y
x_PM_HB3XP67_ASAP7_75T_SRAM%6 N_6_M1_s N_6_M0_d VSS PM_HB3XP67_ASAP7_75T_SRAM%6
x_PM_HB3XP67_ASAP7_75T_SRAM%7 N_7_M2_s N_7_M1_d VSS PM_HB3XP67_ASAP7_75T_SRAM%7
x_PM_HB3XP67_ASAP7_75T_SRAM%8 N_8_M5_s N_8_M4_d VSS PM_HB3XP67_ASAP7_75T_SRAM%8
x_PM_HB3XP67_ASAP7_75T_SRAM%9 N_9_M6_s N_9_M5_d VSS PM_HB3XP67_ASAP7_75T_SRAM%9
cc_1 N_A_M1_g N_4_M3_g 2.34385e-19 $X=0.135 $Y=0.0405 $X2=0.243 $Y2=0.054
cc_2 N_A_M2_g N_4_M3_g 0.00287079f $X=0.189 $Y=0.0405 $X2=0.243 $Y2=0.054
cc_3 N_A_c_3_p N_4_c_37_n 0.0014668f $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.135
cc_4 N_A_M1_g N_4_c_38_n 2.00459e-19 $X=0.135 $Y=0.0405 $X2=0.18 $Y2=0.036
cc_5 N_A_M2_g N_4_c_38_n 2.0666e-19 $X=0.189 $Y=0.0405 $X2=0.18 $Y2=0.036
cc_6 N_A_c_6_p N_4_c_40_n 3.03951e-19 $X=0.046 $Y=0.135 $X2=0.054 $Y2=0.036
cc_7 N_A_c_7_p N_4_c_40_n 3.03951e-19 $X=0.0635 $Y=0.135 $X2=0.054 $Y2=0.036
cc_8 N_A_c_8_p N_4_c_40_n 5.65154e-19 $X=0.018 $Y=0.135 $X2=0.054 $Y2=0.036
cc_9 N_A_M0_g N_4_c_43_n 4.28653e-19 $X=0.081 $Y=0.0405 $X2=0.095 $Y2=0.036
cc_10 N_A_c_3_p N_4_c_43_n 0.00132028f $X=0.189 $Y=0.135 $X2=0.095 $Y2=0.036
cc_11 N_A_c_11_p N_4_c_43_n 3.03951e-19 $X=0.081 $Y=0.135 $X2=0.095 $Y2=0.036
cc_12 N_A_M1_g N_4_c_46_n 3.45619e-19 $X=0.135 $Y=0.0405 $X2=0.1375 $Y2=0.036
cc_13 N_A_M1_g N_4_c_47_n 2.00459e-19 $X=0.135 $Y=0.0405 $X2=0.18 $Y2=0.234
cc_14 N_A_M2_g N_4_c_47_n 2.0666e-19 $X=0.189 $Y=0.0405 $X2=0.18 $Y2=0.234
cc_15 A N_4_c_49_n 5.65154e-19 $X=0.02 $Y=0.1585 $X2=0.054 $Y2=0.234
cc_16 N_A_c_6_p N_4_c_49_n 3.03951e-19 $X=0.046 $Y=0.135 $X2=0.054 $Y2=0.234
cc_17 N_A_c_7_p N_4_c_49_n 3.03951e-19 $X=0.0635 $Y=0.135 $X2=0.054 $Y2=0.234
cc_18 N_A_M0_g N_4_c_52_n 4.28653e-19 $X=0.081 $Y=0.0405 $X2=0.095 $Y2=0.234
cc_19 N_A_c_3_p N_4_c_52_n 0.00132028f $X=0.189 $Y=0.135 $X2=0.095 $Y2=0.234
cc_20 N_A_c_11_p N_4_c_52_n 3.03951e-19 $X=0.081 $Y=0.135 $X2=0.095 $Y2=0.234
cc_21 N_A_M1_g N_4_c_55_n 3.45619e-19 $X=0.135 $Y=0.0405 $X2=0.1375 $Y2=0.234
cc_22 N_A_M2_g N_4_c_56_n 7.88673e-19 $X=0.189 $Y=0.0405 $X2=0.189 $Y2=0.126
cc_23 N_A_c_3_p N_4_c_56_n 5.09138e-19 $X=0.189 $Y=0.135 $X2=0.189 $Y2=0.126
cc_24 N_A_c_8_p N_4_c_56_n 4.86282e-19 $X=0.018 $Y=0.135 $X2=0.189 $Y2=0.126
cc_25 N_A_M2_g N_4_c_59_n 3.58231e-19 $X=0.189 $Y=0.0405 $X2=0.189 $Y2=0.081
cc_26 N_A_c_8_p N_4_c_59_n 2.85111e-19 $X=0.018 $Y=0.135 $X2=0.189 $Y2=0.081
cc_27 N_A_M2_g N_4_c_61_n 7.88673e-19 $X=0.189 $Y=0.0405 $X2=0.189 $Y2=0.189
cc_28 N_A_c_3_p N_4_c_61_n 5.09138e-19 $X=0.189 $Y=0.135 $X2=0.189 $Y2=0.189
cc_29 A N_4_c_61_n 4.86282e-19 $X=0.02 $Y=0.1585 $X2=0.189 $Y2=0.189
cc_30 N_A_M2_g N_4_c_64_n 3.58231e-19 $X=0.189 $Y=0.0405 $X2=0.189 $Y2=0.207
cc_31 A N_4_c_64_n 2.85111e-19 $X=0.02 $Y=0.1585 $X2=0.189 $Y2=0.207
cc_32 N_A_c_3_p N_4_c_66_n 5.49186e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.135
cc_33 N_A_c_3_p N_4_c_67_n 0.00129387f $X=0.189 $Y=0.135 $X2=0.189 $Y2=0.135
cc_34 N_A_c_11_p N_4_c_67_n 2.96499e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_35 N_4_c_61_n N_Y_c_75_n 0.00115681f $X=0.189 $Y=0.189 $X2=0.135 $Y2=0.135
cc_36 N_4_c_70_p N_Y_c_76_n 0.00115681f $X=0.189 $Y=0.063 $X2=0.135 $Y2=0.2295
cc_37 N_4_c_37_n N_Y_c_77_n 3.15821e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_38 N_4_c_66_n N_Y_c_77_n 0.00102675f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_39 N_4_c_38_n N_Y_c_79_n 3.78293e-19 $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.0405
cc_40 N_4_c_47_n N_Y_c_80_n 3.78293e-19 $X=0.18 $Y=0.234 $X2=0 $Y2=0

* END of "./HB3xp67_ASAP7_75t_SRAM.pex.sp.HB3XP67_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

* File: HB4xp67_ASAP7_75t_SRAM.pex.sp
* Created: Tue Sep  5 12:31:14 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "HB4xp67_ASAP7_75t_SRAM.pex.sp.pex"
* BEGIN of "./HB4xp67_ASAP7_75t_SRAM.pex.sp.pex"
* File: HB4xp67_ASAP7_75t_SRAM.pex.sp.pex
* Created: Tue Sep  5 12:31:14 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_HB4XP67_ASAP7_75T_SRAM%A 2 7 10 15 18 23 26 29 31 38 41 43 44 48 VSS
c37 48 VSS 0.00527166f $X=0.018 $Y=0.135
c38 44 VSS 3.72004e-19 $X=0.0635 $Y=0.135
c39 43 VSS 7.23977e-19 $X=0.046 $Y=0.135
c40 41 VSS 1.33597e-19 $X=0.081 $Y=0.135
c41 38 VSS 0.00594103f $X=0.021 $Y=0.1565
c42 29 VSS 0.0118251f $X=0.243 $Y=0.135
c43 26 VSS 0.0629072f $X=0.243 $Y=0.0405
c44 18 VSS 0.0649884f $X=0.189 $Y=0.0405
c45 10 VSS 0.0654789f $X=0.135 $Y=0.0405
c46 2 VSS 0.0687797f $X=0.081 $Y=0.0405
r47 43 44 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.046
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r48 41 44 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0635 $Y2=0.135
r49 39 48 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r50 39 43 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.046 $Y2=0.135
r51 35 48 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r52 35 38 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.1565
r53 29 31 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2295
r54 26 29 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0405 $X2=0.243 $Y2=0.135
r55 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r56 21 23 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2295
r57 18 21 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0405 $X2=0.189 $Y2=0.135
r58 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r59 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2295
r60 10 13 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0405 $X2=0.135 $Y2=0.135
r61 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r62 5 41 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r63 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2295
r64 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0405 $X2=0.081 $Y2=0.135
.ends

.subckt PM_HB4XP67_ASAP7_75T_SRAM%4 2 5 7 9 14 19 21 26 27 28 30 35 36 38 39 40 42
+ 43 44 47 51 VSS
c41 47 VSS 0.00472678f $X=0.297 $Y=0.135
c42 44 VSS 3.30481e-19 $X=0.189 $Y=0.207
c43 43 VSS 7.9698e-19 $X=0.189 $Y=0.189
c44 42 VSS 2.81339e-19 $X=0.189 $Y=0.225
c45 40 VSS 3.13346e-19 $X=0.189 $Y=0.099
c46 39 VSS 8.6896e-19 $X=0.189 $Y=0.081
c47 38 VSS 4.66155e-19 $X=0.189 $Y=0.126
c48 36 VSS 0.00408275f $X=0.1375 $Y=0.234
c49 35 VSS 0.00363755f $X=0.095 $Y=0.234
c50 30 VSS 0.00188634f $X=0.054 $Y=0.234
c51 28 VSS 0.00689504f $X=0.18 $Y=0.234
c52 27 VSS 0.00408275f $X=0.1375 $Y=0.036
c53 26 VSS 0.00363755f $X=0.095 $Y=0.036
c54 21 VSS 0.00189187f $X=0.054 $Y=0.036
c55 19 VSS 0.00689504f $X=0.18 $Y=0.036
c56 17 VSS 0.00231457f $X=0.056 $Y=0.2295
c57 14 VSS 2.67274e-19 $X=0.071 $Y=0.2295
c58 12 VSS 0.00231786f $X=0.056 $Y=0.0405
c59 9 VSS 2.67274e-19 $X=0.071 $Y=0.0405
c60 5 VSS 0.00239754f $X=0.297 $Y=0.135
c61 2 VSS 0.0664863f $X=0.297 $Y=0.054
r62 45 51 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.135 $X2=0.189 $Y2=0.135
r63 45 47 6.72222 $w=1.8e-08 $l=9.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.135 $X2=0.297 $Y2=0.135
r64 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.207
r65 42 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.207
r66 41 51 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.135
r67 41 43 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.189
r68 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.081 $X2=0.189 $Y2=0.099
r69 38 51 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.135
r70 38 40 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.126 $X2=0.189 $Y2=0.099
r71 37 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.081
r72 35 36 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.234 $X2=0.1375 $Y2=0.234
r73 30 35 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.095 $Y2=0.234
r74 28 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.234 $X2=0.189 $Y2=0.225
r75 28 36 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.1375 $Y2=0.234
r76 26 27 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.036 $X2=0.1375 $Y2=0.036
r77 21 26 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.095 $Y2=0.036
r78 19 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r79 19 27 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.1375 $Y2=0.036
r80 17 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r81 14 17 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2295 $X2=0.056 $Y2=0.2295
r82 12 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r83 9 12 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0405 $X2=0.056 $Y2=0.0405
r84 5 47 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r85 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r86 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
.ends

.subckt PM_HB4XP67_ASAP7_75T_SRAM%Y 1 6 12 14 16 VSS
c4 34 VSS 0.00270568f $X=0.342 $Y=0.234
c5 33 VSS 0.00278493f $X=0.351 $Y=0.234
c6 28 VSS 0.00176131f $X=0.324 $Y=0.234
c7 24 VSS 0.00270568f $X=0.342 $Y=0.036
c8 23 VSS 0.00278493f $X=0.351 $Y=0.036
c9 18 VSS 0.00176131f $X=0.324 $Y=0.036
c10 16 VSS 7.46953e-19 $X=0.351 $Y=0.144
c11 14 VSS 0.00448156f $X=0.3515 $Y=0.1145
c12 12 VSS 0.00448156f $X=0.351 $Y=0.225
c13 9 VSS 0.00547928f $X=0.322 $Y=0.216
c14 4 VSS 0.00547928f $X=0.322 $Y=0.054
r15 34 35 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.3465 $Y2=0.234
r16 33 35 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.234 $X2=0.3465 $Y2=0.234
r17 28 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.342 $Y2=0.234
r18 24 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.3465 $Y2=0.036
r19 23 25 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.036 $X2=0.3465 $Y2=0.036
r20 18 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r21 15 16 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.144
r22 14 15 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1145 $X2=0.351 $Y2=0.126
r23 12 33 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.234
r24 12 16 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.144
r25 11 23 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.036
r26 11 14 4.71914 $w=1.8e-08 $l=6.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.1145
r27 9 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r28 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.216 $X2=0.322 $Y2=0.216
r29 4 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r30 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.054 $X2=0.322 $Y2=0.054
.ends

.subckt PM_HB4XP67_ASAP7_75T_SRAM%6 1 2 VSS
c0 1 VSS 0.00192428f $X=0.125 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0405 $X2=0.091 $Y2=0.0405
.ends

.subckt PM_HB4XP67_ASAP7_75T_SRAM%7 1 2 VSS
c0 1 VSS 0.00194494f $X=0.179 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0405 $X2=0.145 $Y2=0.0405
.ends

.subckt PM_HB4XP67_ASAP7_75T_SRAM%8 1 2 VSS
c0 1 VSS 0.00214045f $X=0.233 $Y=0.0405
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0405 $X2=0.199 $Y2=0.0405
.ends

.subckt PM_HB4XP67_ASAP7_75T_SRAM%9 1 2 VSS
c0 1 VSS 0.00192428f $X=0.125 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2295 $X2=0.091 $Y2=0.2295
.ends

.subckt PM_HB4XP67_ASAP7_75T_SRAM%10 1 2 VSS
c0 1 VSS 0.00194494f $X=0.179 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2295 $X2=0.145 $Y2=0.2295
.ends

.subckt PM_HB4XP67_ASAP7_75T_SRAM%11 1 2 VSS
c0 1 VSS 0.00214045f $X=0.233 $Y=0.2295
r1 1 2 50.3704 $w=2.7e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2295 $X2=0.199 $Y2=0.2295
.ends


* END of "./HB4xp67_ASAP7_75t_SRAM.pex.sp.pex"
* 
.subckt HB4xp67_ASAP7_75t_SRAM  VSS VDD A Y
* 
* Y	Y
* A	A
M0 N_6_M0_d N_A_M0_g N_4_M0_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071
+ $Y=0.027
M1 N_7_M1_d N_A_M1_g N_6_M1_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.125
+ $Y=0.027
M2 N_8_M2_d N_A_M2_g N_7_M2_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.179
+ $Y=0.027
M3 VSS N_A_M3_g N_8_M3_s VSS NMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_4_M4_g VSS VSS NMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.287 $Y=0.027
M5 N_9_M5_d N_A_M5_g N_4_M5_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.071
+ $Y=0.216
M6 N_10_M6_d N_A_M6_g N_9_M6_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.125
+ $Y=0.216
M7 N_11_M7_d N_A_M7_g N_10_M7_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.179
+ $Y=0.216
M8 VDD N_A_M8_g N_11_M8_s VDD PMOS_SRAM L=2e-08 W=2.7e-08 NFIN=1 $X=0.233
+ $Y=0.216
M9 N_Y_M9_d N_4_M9_g VDD VDD PMOS_SRAM L=2e-08 W=5.4e-08 NFIN=2 $X=0.287 $Y=0.189
*
* 
* .include "HB4xp67_ASAP7_75t_SRAM.pex.sp.HB4XP67_ASAP7_75T_SRAM.pxi"
* BEGIN of "./HB4xp67_ASAP7_75t_SRAM.pex.sp.HB4XP67_ASAP7_75T_SRAM.pxi"
* File: HB4xp67_ASAP7_75t_SRAM.pex.sp.HB4XP67_ASAP7_75T_SRAM.pxi
* Created: Tue Sep  5 12:31:14 2017
* 
x_PM_HB4XP67_ASAP7_75T_SRAM%A N_A_M0_g N_A_M5_g N_A_M1_g N_A_M6_g N_A_M2_g N_A_M7_g
+ N_A_M3_g N_A_c_3_p N_A_M8_g A N_A_c_11_p N_A_c_6_p N_A_c_7_p N_A_c_8_p VSS
+ PM_HB4XP67_ASAP7_75T_SRAM%A
x_PM_HB4XP67_ASAP7_75T_SRAM%4 N_4_M4_g N_4_c_40_n N_4_M9_g N_4_M0_s N_4_M5_s
+ N_4_c_41_n N_4_c_43_n N_4_c_46_n N_4_c_49_n N_4_c_50_n N_4_c_52_n N_4_c_55_n
+ N_4_c_58_n N_4_c_59_n N_4_c_62_n N_4_c_63_n N_4_c_65_n N_4_c_66_n N_4_c_69_n
+ N_4_c_71_n N_4_c_73_n VSS PM_HB4XP67_ASAP7_75T_SRAM%4
x_PM_HB4XP67_ASAP7_75T_SRAM%Y N_Y_M4_d N_Y_M9_d N_Y_c_79_n Y N_Y_c_81_n VSS
+ PM_HB4XP67_ASAP7_75T_SRAM%Y
x_PM_HB4XP67_ASAP7_75T_SRAM%6 N_6_M1_s N_6_M0_d VSS PM_HB4XP67_ASAP7_75T_SRAM%6
x_PM_HB4XP67_ASAP7_75T_SRAM%7 N_7_M2_s N_7_M1_d VSS PM_HB4XP67_ASAP7_75T_SRAM%7
x_PM_HB4XP67_ASAP7_75T_SRAM%8 N_8_M3_s N_8_M2_d VSS PM_HB4XP67_ASAP7_75T_SRAM%8
x_PM_HB4XP67_ASAP7_75T_SRAM%9 N_9_M6_s N_9_M5_d VSS PM_HB4XP67_ASAP7_75T_SRAM%9
x_PM_HB4XP67_ASAP7_75T_SRAM%10 N_10_M7_s N_10_M6_d VSS PM_HB4XP67_ASAP7_75T_SRAM%10
x_PM_HB4XP67_ASAP7_75T_SRAM%11 N_11_M8_s N_11_M7_d VSS PM_HB4XP67_ASAP7_75T_SRAM%11
cc_1 N_A_M2_g N_4_M4_g 2.34385e-19 $X=0.189 $Y=0.0405 $X2=0.297 $Y2=0.054
cc_2 N_A_M3_g N_4_M4_g 0.00287079f $X=0.243 $Y=0.0405 $X2=0.297 $Y2=0.054
cc_3 N_A_c_3_p N_4_c_40_n 0.00151965f $X=0.243 $Y=0.135 $X2=0.297 $Y2=0.135
cc_4 N_A_M1_g N_4_c_41_n 2.00459e-19 $X=0.135 $Y=0.0405 $X2=0.18 $Y2=0.036
cc_5 N_A_M2_g N_4_c_41_n 2.78042e-19 $X=0.189 $Y=0.0405 $X2=0.18 $Y2=0.036
cc_6 N_A_c_6_p N_4_c_43_n 3.04762e-19 $X=0.046 $Y=0.135 $X2=0.054 $Y2=0.036
cc_7 N_A_c_7_p N_4_c_43_n 3.04762e-19 $X=0.0635 $Y=0.135 $X2=0.054 $Y2=0.036
cc_8 N_A_c_8_p N_4_c_43_n 3.29221e-19 $X=0.018 $Y=0.135 $X2=0.054 $Y2=0.036
cc_9 N_A_M0_g N_4_c_46_n 4.28653e-19 $X=0.081 $Y=0.0405 $X2=0.095 $Y2=0.036
cc_10 N_A_c_3_p N_4_c_46_n 0.00132028f $X=0.243 $Y=0.135 $X2=0.095 $Y2=0.036
cc_11 N_A_c_11_p N_4_c_46_n 3.04762e-19 $X=0.081 $Y=0.135 $X2=0.095 $Y2=0.036
cc_12 N_A_M1_g N_4_c_49_n 3.45619e-19 $X=0.135 $Y=0.0405 $X2=0.1375 $Y2=0.036
cc_13 N_A_M1_g N_4_c_50_n 2.00459e-19 $X=0.135 $Y=0.0405 $X2=0.18 $Y2=0.234
cc_14 N_A_M2_g N_4_c_50_n 2.78042e-19 $X=0.189 $Y=0.0405 $X2=0.18 $Y2=0.234
cc_15 A N_4_c_52_n 5.65154e-19 $X=0.021 $Y=0.1565 $X2=0.054 $Y2=0.234
cc_16 N_A_c_6_p N_4_c_52_n 3.03951e-19 $X=0.046 $Y=0.135 $X2=0.054 $Y2=0.234
cc_17 N_A_c_7_p N_4_c_52_n 3.03951e-19 $X=0.0635 $Y=0.135 $X2=0.054 $Y2=0.234
cc_18 N_A_M0_g N_4_c_55_n 4.28653e-19 $X=0.081 $Y=0.0405 $X2=0.095 $Y2=0.234
cc_19 N_A_c_3_p N_4_c_55_n 0.00132028f $X=0.243 $Y=0.135 $X2=0.095 $Y2=0.234
cc_20 N_A_c_11_p N_4_c_55_n 3.03951e-19 $X=0.081 $Y=0.135 $X2=0.095 $Y2=0.234
cc_21 N_A_M1_g N_4_c_58_n 3.45619e-19 $X=0.135 $Y=0.0405 $X2=0.1375 $Y2=0.234
cc_22 N_A_M2_g N_4_c_59_n 4.57633e-19 $X=0.189 $Y=0.0405 $X2=0.189 $Y2=0.126
cc_23 N_A_c_3_p N_4_c_59_n 5.21939e-19 $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.126
cc_24 N_A_c_8_p N_4_c_59_n 2.85496e-19 $X=0.018 $Y=0.135 $X2=0.189 $Y2=0.126
cc_25 N_A_M2_g N_4_c_62_n 6.84745e-19 $X=0.189 $Y=0.0405 $X2=0.189 $Y2=0.081
cc_26 N_A_M2_g N_4_c_63_n 4.58544e-19 $X=0.189 $Y=0.0405 $X2=0.189 $Y2=0.099
cc_27 N_A_c_8_p N_4_c_63_n 2.85111e-19 $X=0.018 $Y=0.135 $X2=0.189 $Y2=0.099
cc_28 N_A_M2_g N_4_c_65_n 2.54412e-19 $X=0.189 $Y=0.0405 $X2=0.189 $Y2=0.225
cc_29 N_A_M2_g N_4_c_66_n 9.28674e-19 $X=0.189 $Y=0.0405 $X2=0.189 $Y2=0.189
cc_30 N_A_c_3_p N_4_c_66_n 5.21939e-19 $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.189
cc_31 A N_4_c_66_n 4.86282e-19 $X=0.021 $Y=0.1565 $X2=0.189 $Y2=0.189
cc_32 N_A_M2_g N_4_c_69_n 4.16582e-19 $X=0.189 $Y=0.0405 $X2=0.189 $Y2=0.207
cc_33 A N_4_c_69_n 2.85111e-19 $X=0.021 $Y=0.1565 $X2=0.189 $Y2=0.207
cc_34 N_A_M3_g N_4_c_71_n 8.19974e-19 $X=0.243 $Y=0.0405 $X2=0.297 $Y2=0.135
cc_35 N_A_c_3_p N_4_c_71_n 0.00489613f $X=0.243 $Y=0.135 $X2=0.297 $Y2=0.135
cc_36 N_A_c_3_p N_4_c_73_n 0.00131846f $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.135
cc_37 N_A_c_11_p N_4_c_73_n 3.02259e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_38 N_4_c_66_n N_Y_c_79_n 6.90454e-19 $X=0.189 $Y=0.189 $X2=0.135 $Y2=0.135
cc_39 N_4_c_62_n Y 6.90509e-19 $X=0.189 $Y=0.081 $X2=0.135 $Y2=0.2295
cc_40 N_4_c_40_n N_Y_c_81_n 3.15821e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_41 N_4_c_71_n N_Y_c_81_n 0.00103578f $X=0.297 $Y=0.135 $X2=0 $Y2=0

* END of "./HB4xp67_ASAP7_75t_SRAM.pex.sp.HB4XP67_ASAP7_75T_SRAM.pxi"
* 
*
.ends
*
*

