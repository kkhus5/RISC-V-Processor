************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: A2O1A1Ixp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:34 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    A2O1A1Ixp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT A2O1A1Ixp33_ASAP7_75t_L A1 A2 B C VDD VSS Y
*.PININFO A1:I A2:I B:I C:I Y:O VDD:B VSS:B
MM7 net06 B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 Y C net06 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net015 A2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net06 A1 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 Y C VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM5 Y B net2 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net2 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net2 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: A2O1A1O1Ixp25_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:35 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    A2O1A1O1Ixp25_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT A2O1A1O1Ixp25_ASAP7_75t_L A1 A2 B C D VDD VSS Y
*.PININFO A1:I A2:I B:I C:I D:I Y:O VDD:B VSS:B
MM5 net4 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net15 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net4 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 Y D net15 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net15 B net4 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 Y D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net25 A2 net12 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 Y B net12 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y A1 net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net12 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AND2x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:36 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AND2x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AND2x2_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM4 Y net10 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 net10 B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM0 net10 A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM5 Y net10 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM3 net20 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net10 B net20 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AND2x4_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:37 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AND2x4_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AND2x4_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM4 Y net9 VDD VDD pmos_lvt w=324.00n l=20n nfin=12
MM1 net9 B VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM0 net9 A VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM5 Y net9 VSS VSS nmos_lvt w=324.00n l=20n nfin=12
MM3 net19 A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 net9 B net19 VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AND2x6_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:39 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AND2x6_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AND2x6_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM4 Y net9 VDD VDD pmos_lvt w=486.00n l=20n nfin=18
MM1 net9 B VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM0 net9 A VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM5 Y net9 VSS VSS nmos_lvt w=486.00n l=20n nfin=18
MM3 net19 A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 net9 B net19 VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AND3x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:40 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AND3x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AND3x1_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM6 Y net61 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net61 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net61 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net61 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 Y net61 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net61 A net72 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net72 B net71 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net71 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AND3x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:41 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AND3x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AND3x2_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM6 Y net61 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM5 net61 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net61 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net61 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 Y net61 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 net61 A net72 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net72 B net71 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net71 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AND3x4_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:42 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AND3x4_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AND3x4_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM6 Y net83 VDD VDD pmos_lvt w=324.00n l=20n nfin=12
MM5 net83 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net83 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net83 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 Y net83 VSS VSS nmos_lvt w=324.00n l=20n nfin=12
MM0 net83 A net89 VSS nmos_lvt w=162.00n l=20n nfin=6
MM1 net89 B net90 VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 net90 C VSS VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AND4x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:43 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AND4x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AND4x1_ASAP7_75t_L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MM8 Y net12 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net12 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net12 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net12 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net12 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 Y net12 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 pd3 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 pd2 B pd3 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 pd1 C pd2 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net12 D pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AND4x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:45 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AND4x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AND4x2_ASAP7_75t_L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MM5 net33 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net33 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net33 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net33 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 Y net33 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM9 net15 D VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM8 net16 C net15 VSS nmos_lvt w=162.00n l=20n nfin=6
MM7 net17 B net16 VSS nmos_lvt w=162.00n l=20n nfin=6
MM6 net33 A net17 VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 Y net33 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AND5x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:46 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AND5x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AND5x1_ASAP7_75t_L A B C D E VDD VSS Y
*.PININFO A:I B:I C:I D:I E:I Y:O VDD:B VSS:B
MM11 Y net011 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net29 E VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net30 D net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 net024 B net023 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net011 A net024 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net023 C net30 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net011 E VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM8 net011 D VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM7 net011 C VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 net011 B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 Y net011 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net011 A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AND5x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:47 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AND5x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AND5x2_ASAP7_75t_L A B C D E VDD VSS Y
*.PININFO A:I B:I C:I D:I E:I Y:O VDD:B VSS:B
MM1 Y net14 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM9 net14 E VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net14 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net14 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net14 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net14 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 Y net14 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM6 net33 E VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM5 net34 D net33 VSS nmos_lvt w=162.00n l=20n nfin=6
MM4 net32 B net35 VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 net14 A net32 VSS nmos_lvt w=162.00n l=20n nfin=6
MM3 net35 C net34 VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO211x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:48 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO211x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO211x2_ASAP7_75t_L A1 A2 B C VDD VSS Y
*.PININFO A1:I A2:I B:I C:I Y:O VDD:B VSS:B
MM8 Y net014 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM4 net014 C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 net014 B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 net23 A2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 net014 A1 net23 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 Y net014 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 net014 C net22 VDD pmos_lvt w=162.00n l=20n nfin=6
MM5 net22 B net20 VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 net20 A2 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM25 net20 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO21x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:49 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO21x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO21x1_ASAP7_75t_L A1 A2 B VDD VSS Y
*.PININFO A1:I A2:I B:I Y:O VDD:B VSS:B
MM7 Y net16 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 net16 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net16 A1 net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net29 A2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 Y net16 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net18 A2 net16 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 VDD B net18 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net18 A1 net16 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO21x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:50 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO21x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO21x2_ASAP7_75t_L A1 A2 B VDD VSS Y
*.PININFO A1:I A2:I B:I Y:O VDD:B VSS:B
MM7 Y net16 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM4 net16 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net16 A1 net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net29 A2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 Y net16 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM5 net18 A2 net16 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 VDD B net18 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net18 A1 net16 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO221x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:52 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO221x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO221x1_ASAP7_75t_L A1 A2 B1 B2 C VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C:I Y:O VDD:B VSS:B
MM4 Y yn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM28 yn C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM27 net23 B2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM26 yn B1 net23 VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 yn A1 net24 VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 net24 A2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 Y yn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 s1 C s2 VDD pmos_lvt w=81.0n l=20n nfin=3
MM32 s2 B2 yn VDD pmos_lvt w=81.0n l=20n nfin=3
MM31 s1 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM30 s2 B1 yn VDD pmos_lvt w=81.0n l=20n nfin=3
MM29 s1 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO221x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:53 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO221x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO221x2_ASAP7_75t_L A1 A2 B1 B2 C VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C:I Y:O VDD:B VSS:B
MM4 Y yn VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM28 yn C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM27 net23 B2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM26 yn B1 net23 VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 yn A1 net24 VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 net24 A2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 Y yn VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 s1 C s2 VDD pmos_lvt w=81.0n l=20n nfin=3
MM32 s2 B2 yn VDD pmos_lvt w=81.0n l=20n nfin=3
MM31 s1 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM30 s2 B1 yn VDD pmos_lvt w=81.0n l=20n nfin=3
MM29 s1 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO222x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:54 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO222x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO222x2_ASAP7_75t_L A1 A2 B1 B2 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I Y:O VDD:B VSS:B
MM8 Y net23 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM5 net23 C2 net17 VDD pmos_lvt w=162.00n l=20n nfin=6
MM4 net17 B2 net18 VDD pmos_lvt w=162.00n l=20n nfin=6
MM3 net18 A2 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM2 net23 C1 net17 VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 net17 B1 net18 VDD pmos_lvt w=162.00n l=20n nfin=6
MM0 net18 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM14 net37 B2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 net23 B1 net37 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net36 C2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net23 C1 net36 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 Y net23 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM7 net38 A2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net23 A1 net38 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO22x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:55 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO22x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO22x1_ASAP7_75t_L A1 A2 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I Y:O VDD:B VSS:B
MM5 net18 B2 net13 VDD pmos_lvt w=54.0n l=20n nfin=2
MM4 net18 B1 net13 VDD pmos_lvt w=54.0n l=20n nfin=2
MM3 net13 A2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 Y net18 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net13 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM9 net29 B1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM8 net30 A1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM7 net18 B2 net29 VSS nmos_lvt w=54.0n l=20n nfin=2
MM6 net18 A2 net30 VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 Y net18 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO22x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:56 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO22x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO22x2_ASAP7_75t_L A1 A2 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I Y:O VDD:B VSS:B
MM5 net18 B2 net13 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net18 B1 net13 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net13 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 Y net18 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM2 net13 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 net29 B1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net30 A1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 net18 B2 net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net18 A2 net30 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y net18 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO31x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:58 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO31x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO31x2_ASAP7_75t_L A1 A2 A3 B VDD VSS Y
*.PININFO A1:I A2:I A3:I B:I Y:O VDD:B VSS:B
MM0 Y net18 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM5 net18 B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 net29 A3 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 net18 A1 net30 VSS nmos_lvt w=162.00n l=20n nfin=6
MM3 net30 A2 net29 VSS nmos_lvt w=162.00n l=20n nfin=6
MM1 Y net18 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM9 net18 B net23 VDD pmos_lvt w=162.00n l=20n nfin=6
MM10 net23 A3 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM7 net23 A2 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 net23 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO322x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:49:59 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO322x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO322x2_ASAP7_75t_L A1 A2 A3 B1 B2 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I C1:I C2:I Y:O VDD:B VSS:B
MM16 Y net25 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM6 net50 C2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 net25 C1 net50 VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 net51 B2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 net25 B1 net51 VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 net52 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net49 A2 net52 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net25 A1 net49 VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 Y net25 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM13 net27 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net25 C2 net53 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net53 B2 net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net27 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 net25 C1 net53 VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net53 B1 net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net27 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO32x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:00 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO32x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO32x1_ASAP7_75t_L A1 A2 A3 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I Y:O VDD:B VSS:B
MM21 Y net08 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net08 A1 net24 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net24 A2 net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net25 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 net26 B2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM13 net08 B1 net26 VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 Y net08 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net10 A2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM4 net10 A3 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM5 net10 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM15 net08 B2 net10 VDD pmos_lvt w=54.0n l=20n nfin=2
MM14 net08 B1 net10 VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO32x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:01 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO32x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO32x2_ASAP7_75t_L A1 A2 A3 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I Y:O VDD:B VSS:B
MM21 Y net08 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 net08 A1 net24 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net24 A2 net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net25 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 net26 B2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM13 net08 B1 net26 VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 Y net08 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 net10 A2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM4 net10 A3 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM5 net10 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM15 net08 B2 net10 VDD pmos_lvt w=54.0n l=20n nfin=2
MM14 net08 B1 net10 VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO331x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:02 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO331x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO331x1_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C:I Y:O VDD:B VSS:B
MM0 Y yb VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM23 net24 B3 net034 VDD pmos_lvt w=81.0n l=20n nfin=3
MM26 net034 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 net24 B2 net034 VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 net034 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM27 yb C net24 VDD pmos_lvt w=81.0n l=20n nfin=3
MM20 net24 B1 net034 VDD pmos_lvt w=81.0n l=20n nfin=3
MM24 net034 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 Y yb VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM22 yb C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM19 net31 B3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 net32 B2 net31 VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 yb B1 net32 VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 n2 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM15 n1 A2 n2 VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 yb A1 n1 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO331x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:04 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO331x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO331x2_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C:I Y:O VDD:B VSS:B
MM0 Y yb VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM23 net24 B3 net034 VDD pmos_lvt w=81.0n l=20n nfin=3
MM26 net034 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 net24 B2 net034 VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 net034 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM27 yb C net24 VDD pmos_lvt w=81.0n l=20n nfin=3
MM20 net24 B1 net034 VDD pmos_lvt w=81.0n l=20n nfin=3
MM24 net034 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 Y yb VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM22 yb C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM19 net31 B3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 net32 B2 net31 VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 yb B1 net32 VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 n2 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM15 n1 A2 n2 VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 yb A1 n1 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO332x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:05 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO332x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO332x1_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I Y:O VDD:B VSS:B
MM17 net018 C1 net061 VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 net061 C2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 Y net018 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net018 B1 net063 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net063 B2 net064 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net064 B3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net25 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 net018 A1 net26 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net26 A2 net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM15 Y net018 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 net031 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net031 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net031 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net030 B1 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net018 C1 net030 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net030 B2 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net030 B3 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net018 C2 net030 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO332x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:06 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO332x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO332x2_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I Y:O VDD:B VSS:B
MM17 net018 C1 net061 VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 net061 C2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 Y net018 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM12 net018 B1 net063 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net063 B2 net064 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net064 B3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net25 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 net018 A1 net26 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net26 A2 net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM15 Y net018 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM9 net031 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net031 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net031 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net030 B1 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net018 C1 net030 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net030 B2 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net030 B3 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net018 C2 net030 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO333x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:07 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO333x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO333x1_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 C3 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I C3:I Y:O VDD:B VSS:B
MM3 Y net40 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net40 C1 net55 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net55 C2 net54 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net54 C3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM19 net58 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 net59 A2 net58 VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 net40 A1 net59 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net40 B3 net56 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net56 B2 net57 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net57 B1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 net40 C1 net22 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net40 C2 net22 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net40 C3 net22 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 Y net40 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM17 net24 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM16 net24 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM15 net24 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 net22 B3 net24 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net22 B2 net24 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net22 B1 net24 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO333x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:08 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO333x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO333x2_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 C3 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I C3:I Y:O VDD:B VSS:B
MM3 Y net40 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 net40 C1 net55 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net55 C2 net54 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net54 C3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM19 net58 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 net59 A2 net58 VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 net40 A1 net59 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net40 B3 net56 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net56 B2 net57 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net57 B1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 net40 C1 net22 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net40 C2 net22 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net40 C3 net22 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 Y net40 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM17 net24 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM16 net24 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM15 net24 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 net22 B3 net24 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net22 B2 net24 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net22 B1 net24 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AO33x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:10 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AO33x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AO33x2_ASAP7_75t_L A1 A2 A3 B1 B2 B3 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I Y:O VDD:B VSS:B
MM25 Y net020 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 net020 B3 net15 VDD pmos_lvt w=54.0n l=20n nfin=2
MM5 net15 A3 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM4 net15 A2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM3 net020 B2 net15 VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 net020 B1 net15 VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 net15 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM24 Y net020 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM10 net020 B1 net39 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net022 B3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net39 B2 net022 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 net020 A1 net40 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net024 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net40 A2 net024 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI211x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:11 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI211x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI211x1_ASAP7_75t_L A1 A2 B C VDD VSS Y
*.PININFO A1:I A2:I B:I C:I Y:O VDD:B VSS:B
MM20 Y C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 Y B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 Y A2 net32 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net32 A1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM21 net17 A2 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM0 net17 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 net34 B net17 VDD pmos_lvt w=162.00n l=20n nfin=6
MM7 Y C net34 VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI211xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:12 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI211xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI211xp5_ASAP7_75t_L A1 A2 B C VDD VSS Y
*.PININFO A1:I A2:I B:I C:I Y:O VDD:B VSS:B
MM20 Y C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 Y B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 Y A2 net32 VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 net32 A1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM21 net17 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net17 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net34 B net17 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 Y C net34 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI21x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:13 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI21x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21x1_ASAP7_75t_L A1 A2 B VDD VSS Y
*.PININFO A1:I A2:I B:I Y:O VDD:B VSS:B
MM4 Y B VSS VSS nmos_lvt w=108.00n l=20n nfin=4
MM3 Y A1 net29 VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 net29 A2 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM5 net18 A2 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM0 Y B net18 VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 net18 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI21xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:14 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI21xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21xp33_ASAP7_75t_L A1 A2 B VDD VSS Y
*.PININFO A1:I A2:I B:I Y:O VDD:B VSS:B
MM4 Y B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 Y A1 net29 VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 net29 A2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 net18 A2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM0 Y B net18 VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 net18 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI21xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:15 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI21xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI21xp5_ASAP7_75t_L A1 A2 B VDD VSS Y
*.PININFO A1:I A2:I B:I Y:O VDD:B VSS:B
MM4 Y B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 Y A1 net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net29 A2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net18 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 Y B net18 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net18 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI221x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:17 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI221x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI221x1_ASAP7_75t_L A1 A2 B1 B2 C VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C:I Y:O VDD:B VSS:B
MM28 Y C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM27 net23 B2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM26 Y B1 net23 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 Y A1 net24 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net24 A2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 Y C net16 VDD pmos_lvt w=162.00n l=20n nfin=6
MM32 net16 B2 net10 VDD pmos_lvt w=162.00n l=20n nfin=6
MM31 net10 A2 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM30 net16 B1 net10 VDD pmos_lvt w=162.00n l=20n nfin=6
MM29 net10 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI221xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:18 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI221xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI221xp5_ASAP7_75t_L A1 A2 B1 B2 C VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C:I Y:O VDD:B VSS:B
MM28 Y C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM27 net23 B2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM26 Y B1 net23 VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 Y A1 net24 VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 net24 A2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 net012 C net16 VDD pmos_lvt w=81.0n l=20n nfin=3
MM32 net16 B2 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM31 net012 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM30 net16 B1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM29 net012 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI222xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:19 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI222xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI222xp33_ASAP7_75t_L A1 A2 B1 B2 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I Y:O VDD:B VSS:B
MM6 net50 C2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 Y C1 net50 VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 net51 B2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 Y B1 net51 VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 net49 A2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 Y A1 net49 VSS nmos_lvt w=54.0n l=20n nfin=2
MM12 Y A2 net53 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net53 B2 net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net27 C2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 Y A1 net53 VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net53 B1 net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net27 C1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI22x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:20 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI22x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22x1_ASAP7_75t_L A1 A2 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I Y:O VDD:B VSS:B
MM5 Y A2 net13 VDD pmos_lvt w=162.00n l=20n nfin=6
MM4 Y A1 net13 VDD pmos_lvt w=162.00n l=20n nfin=6
MM3 net13 B2 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM2 net13 B1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM9 net29 B1 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM8 net30 A1 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM7 Y B2 net29 VSS nmos_lvt w=162.00n l=20n nfin=6
MM6 Y A2 net30 VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI22xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:21 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI22xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22xp33_ASAP7_75t_L A1 A2 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I Y:O VDD:B VSS:B
MM5 Y B2 net13 VDD pmos_lvt w=54.0n l=20n nfin=2
MM4 Y B1 net13 VDD pmos_lvt w=54.0n l=20n nfin=2
MM3 net13 A2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 net13 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM9 net29 B1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM8 net30 A1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM7 Y B2 net29 VSS nmos_lvt w=54.0n l=20n nfin=2
MM6 Y A2 net30 VSS nmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI22xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:23 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI22xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI22xp5_ASAP7_75t_L A1 A2 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I Y:O VDD:B VSS:B
MM5 Y B2 net13 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 Y B1 net13 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net13 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net13 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 net29 B1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net30 A1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 Y B2 net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 Y A2 net30 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI311xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:24 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI311xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI311xp33_ASAP7_75t_L A1 A2 A3 B C VDD VSS Y
*.PININFO A1:I A2:I A3:I B:I C:I Y:O VDD:B VSS:B
MM0 Y C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 Y B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 net29 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 Y A1 net30 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net30 A2 net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 Y C net020 VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 net020 B net23 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net23 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net23 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net23 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI31xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:25 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI31xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI31xp33_ASAP7_75t_L A1 A2 A3 B VDD VSS Y
*.PININFO A1:I A2:I A3:I B:I Y:O VDD:B VSS:B
MM5 Y B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 net29 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 Y A1 net30 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net30 A2 net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 Y B net23 VDD pmos_lvt w=54.0n l=20n nfin=2
MM10 net23 A3 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM7 net23 A2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM6 net23 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI31xp67_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:26 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI31xp67_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI31xp67_ASAP7_75t_L A1 A2 A3 B VDD VSS Y
*.PININFO A1:I A2:I A3:I B:I Y:O VDD:B VSS:B
MM5 Y B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 net29 A3 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 Y A1 net30 VSS nmos_lvt w=162.00n l=20n nfin=6
MM3 net30 A2 net29 VSS nmos_lvt w=162.00n l=20n nfin=6
MM9 Y B net23 VDD pmos_lvt w=162.00n l=20n nfin=6
MM10 net23 A3 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM7 net23 A2 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 net23 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI321xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:27 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI321xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI321xp33_ASAP7_75t_L A1 A2 A3 B1 B2 C VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I C:I Y:O VDD:B VSS:B
MM11 Y B2 net026 VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 Y C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 net026 B1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 net29 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 Y A1 net30 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net30 A2 net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 Y B2 net013 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net013 C net23 VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 Y B1 net013 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net23 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net23 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net23 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI322xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:29 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI322xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI322xp5_ASAP7_75t_L A1 A2 A3 B1 B2 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I C1:I C2:I Y:O VDD:B VSS:B
MM6 net50 C2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 Y C1 net50 VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 net51 B2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 Y B1 net51 VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 net52 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net49 A2 net52 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y A1 net49 VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 net53 A3 net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 Y C2 net53 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net53 A2 net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net27 B2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 Y C1 net53 VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net53 A1 net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net27 B1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI32xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:30 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI32xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI32xp33_ASAP7_75t_L A1 A2 A3 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I Y:O VDD:B VSS:B
MM0 Y A1 net24 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net24 A2 net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net25 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 net26 B2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM13 Y B1 net26 VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 net10 A2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM4 net10 A3 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM5 net10 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM15 Y B2 net10 VDD pmos_lvt w=54.0n l=20n nfin=2
MM14 Y B1 net10 VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI331xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:31 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI331xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI331xp33_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I Y:O VDD:B VSS:B
MM17 Y C1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 Y B1 net063 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net063 B2 net064 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net064 B3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net25 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 Y A1 net26 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net26 A2 net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net031 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net031 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net031 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net030 B1 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 Y C1 net030 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net030 B2 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net030 B3 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI332xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:32 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI332xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI332xp33_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I Y:O VDD:B VSS:B
MM17 Y C1 net061 VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 net061 C2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 Y B1 net063 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net063 B2 net064 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net064 B3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net25 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 Y A1 net26 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net26 A2 net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net031 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net031 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net031 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net030 B1 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 Y C1 net030 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net030 B2 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net030 B3 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 Y C2 net030 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI333xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:33 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI333xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI333xp33_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 C3 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I C3:I Y:O VDD:B VSS:B
MM17 Y C1 net061 VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 net061 C2 net062 VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 net062 C3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 Y B1 net063 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net063 B2 net064 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net064 B3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net25 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 Y A1 net26 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net26 A2 net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net031 C1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net031 C2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net031 C3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net030 B1 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 Y A1 net030 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net030 B2 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM15 Y A3 net030 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net030 B3 net031 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 Y A2 net030 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: AOI33xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:35 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    AOI33xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT AOI33xp33_ASAP7_75t_L A1 A2 A3 B1 B2 B3 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I Y:O VDD:B VSS:B
MM44 Y B1 net52 VSS nmos_lvt w=81.0n l=20n nfin=3
MM45 net52 B2 net51 VSS nmos_lvt w=81.0n l=20n nfin=3
MM48 net51 B3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM39 Y A3 net54 VSS nmos_lvt w=81.0n l=20n nfin=3
MM46 net54 A2 net53 VSS nmos_lvt w=81.0n l=20n nfin=3
MM47 net53 A1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM33 net015 A3 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM35 Y B1 net015 VDD pmos_lvt w=54.0n l=20n nfin=2
MM32 net015 A2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM38 Y B2 net015 VDD pmos_lvt w=54.0n l=20n nfin=2
MM31 net015 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM37 Y B3 net015 VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: ASYNC_DFFHx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:36 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    ASYNC_DFFHx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT ASYNC_DFFHx1_ASAP7_75t_L CLK D QN RESET SET VDD VSS
*.PININFO CLK:I D:I RESET:I SET:I QN:O VDD:B VSS:B
MM43 pd3 SET VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 QN SH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM29 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM44 SS RESET VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM34 SH clkn pd3 VSS nmos_lvt w=54.0n l=20n nfin=2
MM48 net020 RESET VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM12 MS clkb SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM33 pd3 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb net020 VSS nmos_lvt w=54.0n l=20n nfin=2
MM8 net020 MS VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM47 MS SET VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM25 QN SH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM28 SS SH net076 VDD pmos_lvt w=54.0n l=20n nfin=2
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM45 net076 RESET VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM46 net079 SET VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM37 pd2 SS net077 VDD pmos_lvt w=54.0n l=20n nfin=2
MM35 SH clkb pd2 VDD pmos_lvt w=54.0n l=20n nfin=2
MM49 net078 RESET VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkn SH VDD pmos_lvt w=27.0n l=20n nfin=1
MM11 net051 MS net078 VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn net051 VDD pmos_lvt w=27n l=20n nfin=1
MM7 MS MH net079 VDD pmos_lvt w=54.0n l=20n nfin=2
MM42 net077 SET VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx10_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:42 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx10_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx10_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 AN A VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 Y AN VDD VDD pmos_lvt w=810.0n l=20n nfin=30
MM2 AN A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM3 Y AN VSS VSS nmos_lvt w=810.0n l=20n nfin=30
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx12_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:43 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx12_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx12_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM1 Y AN VDD VDD pmos_lvt w=972.00n l=20n nfin=36
MM0 AN A VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM3 Y AN VSS VSS nmos_lvt w=972.00n l=20n nfin=36
MM2 AN A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx12f_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:44 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx12f_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx12f_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM1 Y AN VDD VDD pmos_lvt w=972.00n l=20n nfin=36
MM0 AN A VDD VDD pmos_lvt w=324.00n l=20n nfin=12
MM3 Y AN VSS VSS nmos_lvt w=972.00n l=20n nfin=36
MM2 AN A VSS VSS nmos_lvt w=324.00n l=20n nfin=12
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx16f_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:45 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx16f_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx16f_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM1 Y AN VDD VDD pmos_lvt w=1.296u l=20n nfin=48
MM0 AN A VDD VDD pmos_lvt w=324.00n l=20n nfin=12
MM3 Y AN VSS VSS nmos_lvt w=1.296u l=20n nfin=48
MM2 AN A VSS VSS nmos_lvt w=324.00n l=20n nfin=12
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx24_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:47 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx24_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx24_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM1 Y AN VDD VDD pmos_lvt w=1.944u l=20n nfin=72
MM0 AN A VDD VDD pmos_lvt w=324.00n l=20n nfin=12
MM3 Y AN VSS VSS nmos_lvt w=1.944u l=20n nfin=72
MM2 AN A VSS VSS nmos_lvt w=324.00n l=20n nfin=12
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:48 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx2_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM3 Y AN VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 AN A VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 Y AN VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 AN A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx3_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:49 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx3_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx3_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM1 Y AN VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM0 AN A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 AN A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 Y AN VSS VSS nmos_lvt w=243.00n l=20n nfin=9
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx4_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:50 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx4_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx4_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM1 Y AN VDD VDD pmos_lvt w=324.00n l=20n nfin=12
MM0 AN A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 AN A VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 Y AN VSS VSS nmos_lvt w=324.00n l=20n nfin=12
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx4f_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:51 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx4f_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx4f_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM1 Y AN VDD VDD pmos_lvt w=324.00n l=20n nfin=12
MM0 AN A VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM3 Y AN VSS VSS nmos_lvt w=324.00n l=20n nfin=12
MM2 AN A VSS VSS nmos_lvt w=108.00n l=20n nfin=4
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:53 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx5_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM1 Y AN VDD VDD pmos_lvt w=405.00n l=20n nfin=15
MM0 AN A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 Y AN VSS VSS nmos_lvt w=405.00n l=20n nfin=15
MM2 AN A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx6f_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:54 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx6f_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx6f_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM1 Y AN VDD VDD pmos_lvt w=486.00n l=20n nfin=18
MM0 AN A VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM3 Y AN VSS VSS nmos_lvt w=486.00n l=20n nfin=18
MM2 AN A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: BUFx8_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:55 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    BUFx8_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT BUFx8_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 AN A VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM1 Y AN VDD VDD pmos_lvt w=648.00n l=20n nfin=24
MM2 AN A VSS VSS nmos_lvt w=108.00n l=20n nfin=4
MM3 Y AN VSS VSS nmos_lvt w=648.00n l=20n nfin=24
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DFFHQNx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:56 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DFFHQNx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DFFHQNx1_ASAP7_75t_L CLK D QN VDD VSS
*.PININFO CLK:I D:I QN:O VDD:B VSS:B
MM24 QN SH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM17 SH clkn pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkb SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM25 QN SH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkb pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkn SH VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DFFHQNx2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:57 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DFFHQNx2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DFFHQNx2_ASAP7_75t_L CLK D QN VDD VSS
*.PININFO CLK:I D:I QN:O VDD:B VSS:B
MM24 QN net32 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM17 net32 clkn pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 net37 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 net37 net32 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 net29 clkb net32 VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 net29 net15 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 net15 clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net29 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 net15 clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM25 QN net32 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM19 pd4 net37 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 net32 clkb pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM15 net37 net32 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 net29 clkn net32 VDD pmos_lvt w=27n l=20n nfin=1
MM7 net29 net15 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 net29 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 net15 clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 net15 clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DFFHQNx3_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:50:58 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DFFHQNx3_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DFFHQNx3_ASAP7_75t_L CLK D QN VDD VSS
*.PININFO CLK:I D:I QN:O VDD:B VSS:B
MM24 QN SH VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM17 SH clkn pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkb SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM25 QN SH VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkb pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkn SH VDD pmos_lvt w=27.0n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27.0n l=20n nfin=1
MM7 MS MH VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DFFHQx4_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:00 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DFFHQx4_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DFFHQx4_ASAP7_75t_L CLK D Q VDD VSS
*.PININFO CLK:I D:I Q:O VDD:B VSS:B
MM38 Q net049 VSS VSS nmos_lvt w=324.00n l=20n nfin=12
MM24 net049 SH VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM17 SH clkn pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkb SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM25 net049 SH VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkb pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkn SH VDD pmos_lvt w=27.0n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM37 Q net049 VDD VDD pmos_lvt w=324.00n l=20n nfin=12
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DFFLQNx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:01 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DFFLQNx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DFFLQNx1_ASAP7_75t_L CLK D QN VDD VSS
*.PININFO CLK:I D:I QN:O VDD:B VSS:B
MM24 QN SH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM17 SH clkb net0107 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 net0107 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 net029 clkn SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn net0109 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 net0109 net029 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 net029 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 net020 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb net020 VSS nmos_lvt w=81.0n l=20n nfin=3
MM25 QN SH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 net029 clkb SH VDD pmos_lvt w=27n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM19 net0108 SS VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM18 SH clkn net0108 VDD pmos_lvt w=27.0n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM11 net0110 net029 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM10 MH clkb net0110 VDD pmos_lvt w=27.0n l=20n nfin=1
MM7 net029 MH VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM1 MH clkn net06 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net06 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DFFLQNx2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:02 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DFFLQNx2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DFFLQNx2_ASAP7_75t_L CLK D QN VDD VSS
*.PININFO CLK:I D:I QN:O VDD:B VSS:B
MM24 QN SH VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM17 SH clkb pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkn SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM25 QN SH VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkn pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkb SH VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkb pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DFFLQNx3_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:03 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DFFLQNx3_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DFFLQNx3_ASAP7_75t_L CLK D QN VDD VSS
*.PININFO CLK:I D:I QN:O VDD:B VSS:B
MM27 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 QN SH VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM17 SH clkb pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkn SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM26 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM25 QN SH VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkn pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkb SH VDD pmos_lvt w=27n l=20n nfin=1
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkb pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DFFLQx4_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:04 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DFFLQx4_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DFFLQx4_ASAP7_75t_L CLK D Q VDD VSS
*.PININFO CLK:I D:I Q:O VDD:B VSS:B
MM0 Q QN VSS VSS nmos_lvt w=324.00n l=20n nfin=12
MM24 QN SH VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM17 SH clkb pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkn SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 Q QN VDD VDD pmos_lvt w=324.00n l=20n nfin=12
MM25 QN SH VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkn pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkb SH VDD pmos_lvt w=27n l=20n nfin=1
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkb pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DHLx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:06 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DHLx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DHLx1_ASAP7_75t_L CLK D Q VDD VSS
*.PININFO CLK:I D:I Q:O VDD:B VSS:B
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 Q MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net088 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net088 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM25 Q MH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM7 net088 MH VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM11 pd2 net088 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM10 MH clkb pd2 VDD pmos_lvt w=27n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DHLx2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:07 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DHLx2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DHLx2_ASAP7_75t_L CLK D Q VDD VSS
*.PININFO CLK:I D:I Q:O VDD:B VSS:B
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 Q MH VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM6 net088 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net088 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM11 pd2 net088 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM10 MH clkb pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM12 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM25 Q MH VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM7 net088 MH VDD VDD pmos_lvt w=27.0n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DHLx3_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:08 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DHLx3_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DHLx3_ASAP7_75t_L CLK D Q VDD VSS
*.PININFO CLK:I D:I Q:O VDD:B VSS:B
MM24 Q MH VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM6 net29 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net29 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM25 Q MH VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM7 net29 MH VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM11 pd2 net29 VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM10 MH clkb pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM12 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DLLx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:09 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DLLx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DLLx1_ASAP7_75t_L CLK D Q VDD VSS
*.PININFO CLK:I D:I Q:O VDD:B VSS:B
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 Q MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net085 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net085 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 Q MH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM7 net085 MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 net085 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DLLx2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:11 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DLLx2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DLLx2_ASAP7_75t_L CLK D Q VDD VSS
*.PININFO CLK:I D:I Q:O VDD:B VSS:B
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 Q MH VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM6 net085 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net085 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM11 pd2 net085 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM25 Q MH VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM7 net085 MH VDD VDD pmos_lvt w=27n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: DLLx3_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:12 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    DLLx3_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT DLLx3_ASAP7_75t_L CLK D Q VDD VSS
*.PININFO CLK:I D:I Q:O VDD:B VSS:B
MM24 Q MH VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM6 net30 MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 net30 VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 pd1 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM25 Q MH VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM7 net30 MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 net30 VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: FAx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:13 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    FAx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT FAx1_ASAP7_75t_L A B CI CON SN VDD VSS
*.PININFO A:I B:I CI:I CON:O SN:O VDD:B VSS:B
MM22 SN CI net081 VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 net081 B net082 VDD pmos_lvt w=81.0n l=20n nfin=3
MM20 net082 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM15 SN CON net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net027 CI VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 net027 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net027 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 CON A net37 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net37 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net27 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 CON CI net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net27 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 SN CI net080 VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 net080 B net079 VSS nmos_lvt w=81.0n l=20n nfin=3
MM23 net079 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM19 VSS CI net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 VSS B net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 VSS A net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 net067 CON SN VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 VSS B net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 VSS B net36 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS A net25 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net36 A CON VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 net25 CI CON VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: HAxp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:14 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    HAxp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT HAxp5_ASAP7_75t_L A B CON SN VDD VSS
*.PININFO A:I B:I CON:O SN:O VDD:B VSS:B
MM4 net015 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net015 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 SN CON net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 CON B net43 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net43 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net041 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 SN B net041 VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 SN CON VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 CON A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 CON B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: HB1xp67_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:15 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    HB1xp67_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT HB1xp67_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM23 Y net7 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 net7 A VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM22 Y net7 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 net7 A VDD VDD pmos_lvt w=27.0n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: HB2xp67_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:17 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    HB2xp67_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT HB2xp67_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM5 Y Abar VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 net17 A VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM0 Abar A net17 VSS nmos_lvt w=27.0n l=20n nfin=1
MM4 Y Abar VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM3 net16 A VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM2 Abar A net16 VDD pmos_lvt w=27.0n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: HB3xp67_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:18 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    HB3xp67_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT HB3xp67_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM3 Y net11 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 net11 A net18 VDD pmos_lvt w=27n l=20n nfin=1
MM1 net18 A net19 VDD pmos_lvt w=27n l=20n nfin=1
MM0 net19 A VDD VDD pmos_lvt w=27n l=20n nfin=1
MM7 net16 A VSS VSS nmos_lvt w=27n l=20n nfin=1
MM4 Y net11 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 net11 A net17 VSS nmos_lvt w=27n l=20n nfin=1
MM6 net17 A net16 VSS nmos_lvt w=27n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: HB4xp67_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:19 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    HB4xp67_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT HB4xp67_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM9 net16 A net17 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 net17 A VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM3 net5 A net18 VSS nmos_lvt w=27.0n l=20n nfin=1
MM0 Y net5 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM7 net18 A net16 VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 net20 A net21 VDD pmos_lvt w=27.0n l=20n nfin=1
MM5 net21 A VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM2 net5 A net19 VDD pmos_lvt w=27.0n l=20n nfin=1
MM4 net19 A net20 VDD pmos_lvt w=27.0n l=20n nfin=1
MM1 Y net5 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: ICGx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:20 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    ICGx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT ICGx1_ASAP7_75t_L CLK ENA GCLK SE VDD VSS
*.PININFO CLK:I ENA:I SE:I GCLK:O VDD:B VSS:B
MM18 nos1 SE VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM16 gclkn CLK VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH CLK pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 net0121 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 GCLK gclkn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM26 net0121 ENA nos1 VDD pmos_lvt w=54.0n l=20n nfin=2
MM0 gclkn MH VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM2 gclkn CLK net0140 VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net0141 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 net0140 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM13 gclkn CLK net0141 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 MH CLK pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM27 net0121 SE VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM19 net0121 ENA VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 GCLK gclkn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 pd1 net0121 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: ICGx2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:21 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    ICGx2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT ICGx2_ASAP7_75t_L CLK ENA GCLK SE VDD VSS
*.PININFO CLK:I ENA:I SE:I GCLK:O VDD:B VSS:B
MM18 nos1 SE VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM16 gclkn CLK VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM25 GCLK gclkn VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 MH CLK pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 net0121 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM26 net0121 ENA nos1 VDD pmos_lvt w=54.0n l=20n nfin=2
MM0 gclkn MH VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM27 net0121 SE VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM13 gclkn CLK net0141 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 net0141 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 net0140 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 gclkn CLK net0140 VSS nmos_lvt w=81.0n l=20n nfin=3
MM19 net0121 ENA VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM9 MH CLK pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 net0121 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 GCLK gclkn VSS VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: ICGx3_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:23 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    ICGx3_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT ICGx3_ASAP7_75t_L CLK ENA GCLK SE VDD VSS
*.PININFO CLK:I ENA:I SE:I GCLK:O VDD:B VSS:B
MM0 gclkn MH VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM16 gclkn CLK VDD VDD pmos_lvt w=108.00n l=20n nfin=4
MM25 GCLK gclkn VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH CLK pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 net14 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM26 net14 ENA nos1 VDD pmos_lvt w=54.0n l=20n nfin=2
MM18 nos1 SE VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM24 GCLK gclkn VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM2 gclkn CLK net056 VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net059 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH CLK pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 net14 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 net056 MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 gclkn CLK net059 VSS nmos_lvt w=81.0n l=20n nfin=3
MM27 net14 SE VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM19 net14 ENA VSS VSS nmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVx11_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:24 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVx11_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVx11_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=891.00n l=20n nfin=33
MM1 Y A VDD VDD pmos_lvt w=891.00n l=20n nfin=33
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVx13_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:25 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVx13_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVx13_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=1.053u l=20n nfin=39
MM1 Y A VDD VDD pmos_lvt w=1.053u l=20n nfin=39
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:26 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVx1_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 Y A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVx2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:27 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVx2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVx2_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM1 Y A VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVx3_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:28 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVx3_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVx3_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM1 Y A VDD VDD pmos_lvt w=243.00n l=20n nfin=9
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVx4_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:30 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVx4_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVx4_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=324.00n l=20n nfin=12
MM1 Y A VDD VDD pmos_lvt w=324.00n l=20n nfin=12
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVx5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:31 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVx5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVx5_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=405.00n l=20n nfin=15
MM1 Y A VDD VDD pmos_lvt w=405.00n l=20n nfin=15
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVx6_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:32 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVx6_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVx6_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=486.00n l=20n nfin=18
MM1 Y A VDD VDD pmos_lvt w=486.00n l=20n nfin=18
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVx8_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:33 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVx8_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVx8_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=648.00n l=20n nfin=24
MM1 Y A VDD VDD pmos_lvt w=648.00n l=20n nfin=24
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVxp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:34 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVxp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVxp33_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM1 Y A VDD VDD pmos_lvt w=27.0n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: INVxp67_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:36 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    INVxp67_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT INVxp67_ASAP7_75t_L A VDD VSS Y
*.PININFO A:I Y:O VDD:B VSS:B
MM0 Y A VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 Y A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: MAJIxp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:37 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    MAJIxp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT MAJIxp5_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM4 net17 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 Y B net17 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net1 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net1 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y A net1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net16 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 Y B net16 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net3 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net3 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 Y A net3 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: MAJx2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:38 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    MAJx2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT MAJx2_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM4 net17 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 maji B net17 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net1 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net1 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 maji A net1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 Y maji VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM9 net16 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 maji B net16 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net3 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net3 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 maji A net3 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 Y maji VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: MAJx3_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:39 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    MAJx3_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT MAJx3_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM4 net17 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 maji B net17 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net1 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net1 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 maji A net1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 Y maji VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM9 net16 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 maji B net16 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net3 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net3 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 maji A net3 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 Y maji VDD VDD pmos_lvt w=243.00n l=20n nfin=9
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND2x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:40 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND2x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2x1_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM3 net16 A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 Y B net16 VSS nmos_lvt w=162.00n l=20n nfin=6
MM1 Y B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 Y A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND2x1p5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:41 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND2x1p5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2x1p5_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM3 net16 A VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM2 Y B net16 VSS nmos_lvt w=243.00n l=20n nfin=9
MM1 Y B VDD VDD pmos_lvt w=135.00n l=20n nfin=5
MM0 Y A VDD VDD pmos_lvt w=135.00n l=20n nfin=5
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND2x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:43 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND2x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2x2_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM3 net16 A VSS VSS nmos_lvt w=324.00n l=20n nfin=12
MM2 Y B net16 VSS nmos_lvt w=324.00n l=20n nfin=12
MM1 Y B VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM0 Y A VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND2xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:44 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND2xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2xp33_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM3 net16 A VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 Y B net16 VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 Y B VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM0 Y A VDD VDD pmos_lvt w=27.0n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND2xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:45 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND2xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2xp5_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM3 net16 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 Y B net16 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 Y B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM0 Y A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND2xp67_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:46 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND2xp67_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND2xp67_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM4 net15 A VSS VSS nmos_lvt w=108.00n l=20n nfin=4
MM3 Y B net15 VSS nmos_lvt w=108.00n l=20n nfin=4
MM5 Y B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 Y A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND3x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:47 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND3x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3x1_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM0 Y A net22 VSS nmos_lvt w=243.00n l=20n nfin=9
MM1 net22 B net21 VSS nmos_lvt w=243.00n l=20n nfin=9
MM2 net21 C VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM3 Y A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 Y B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 Y C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND3x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:49 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND3x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3x2_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM0 Y A net22 VSS nmos_lvt w=486.00n l=20n nfin=18
MM1 net22 B net21 VSS nmos_lvt w=486.00n l=20n nfin=18
MM2 net21 C VSS VSS nmos_lvt w=486.00n l=20n nfin=18
MM3 Y A VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM4 Y B VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM5 Y C VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND3xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:50 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND3xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND3xp33_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM0 Y A net22 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net22 B net21 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net21 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 Y A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM4 Y B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM5 Y C VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND4xp25_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:51 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND4xp25_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4xp25_ASAP7_75t_L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MM5 pd3 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 pd2 C pd3 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 pd1 B pd2 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y A pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 Y D VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM6 Y C VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 Y B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 Y A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND4xp75_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:53 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND4xp75_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND4xp75_ASAP7_75t_L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MM5 pd3 D VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM3 pd2 C pd3 VSS nmos_lvt w=243.00n l=20n nfin=9
MM4 pd1 B pd2 VSS nmos_lvt w=243.00n l=20n nfin=9
MM0 Y A pd1 VSS nmos_lvt w=243.00n l=20n nfin=9
MM7 Y D VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 Y C VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM2 Y B VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 Y A VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NAND5xp2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:54 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NAND5xp2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NAND5xp2_ASAP7_75t_L A B C D E VDD VSS Y
*.PININFO A:I B:I C:I D:I E:I Y:O VDD:B VSS:B
MM6 net29 E VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net30 D net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 net024 B net023 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y A net024 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net023 C net30 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 Y E VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM8 Y D VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM7 Y C VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 Y B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM10 Y A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR2x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:55 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR2x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2x1_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM2 VSS A Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 VSS B Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 net16 B Y VDD pmos_lvt w=162.00n l=20n nfin=6
MM3 VDD A net16 VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR2x1p5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:56 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR2x1p5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2x1p5_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM2 VSS A Y VSS nmos_lvt w=135.00n l=20n nfin=5
MM1 VSS B Y VSS nmos_lvt w=135.00n l=20n nfin=5
MM4 net16 B Y VDD pmos_lvt w=243.00n l=20n nfin=9
MM3 VDD A net16 VDD pmos_lvt w=243.00n l=20n nfin=9
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR2x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:57 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR2x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2x2_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM2 VSS A Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM1 VSS B Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM4 net16 B Y VDD pmos_lvt w=324.00n l=20n nfin=12
MM3 VDD A net16 VDD pmos_lvt w=324.00n l=20n nfin=12
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR2xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:51:58 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR2xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2xp33_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM2 VSS A Y VSS nmos_lvt w=27.0n l=20n nfin=1
MM1 VSS B Y VSS nmos_lvt w=27.0n l=20n nfin=1
MM4 net16 B Y VDD pmos_lvt w=54.0n l=20n nfin=2
MM3 VDD A net16 VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR2xp67_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:00 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR2xp67_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR2xp67_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM2 VSS A Y VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 VSS B Y VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 net16 B Y VDD pmos_lvt w=108.00n l=20n nfin=4
MM3 VDD A net16 VDD pmos_lvt w=108.00n l=20n nfin=4
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR3x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:01 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR3x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3x1_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM14 Y C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 Y B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 Y A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net21 C VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM10 net22 B net21 VDD pmos_lvt w=243.00n l=20n nfin=9
MM11 Y A net22 VDD pmos_lvt w=243.00n l=20n nfin=9
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR3x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:02 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR3x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3x2_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM14 Y C VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM13 Y B VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM12 Y A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM8 net21 C VDD VDD pmos_lvt w=486.00n l=20n nfin=18
MM10 net22 B net21 VDD pmos_lvt w=486.00n l=20n nfin=18
MM11 Y A net22 VDD pmos_lvt w=486.00n l=20n nfin=18
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR3xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:03 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR3xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR3xp33_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM14 Y C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM13 Y B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM12 Y A VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM8 net21 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net22 B net21 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 Y A net22 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR4xp25_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:04 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR4xp25_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4xp25_ASAP7_75t_L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MM7 Y A pd1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 pd1 B pd2 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 pd2 C pd3 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 pd3 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 Y D VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 Y C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 Y B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 Y A VSS VSS nmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR4xp75_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:06 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR4xp75_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR4xp75_ASAP7_75t_L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MM7 Y A pd1 VDD pmos_lvt w=243.00n l=20n nfin=9
MM6 pd1 B pd2 VDD pmos_lvt w=243.00n l=20n nfin=9
MM5 pd2 C pd3 VDD pmos_lvt w=243.00n l=20n nfin=9
MM4 pd3 D VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM3 Y D VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 Y C VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM1 Y B VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 Y A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: NOR5xp2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:07 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    NOR5xp2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT NOR5xp2_ASAP7_75t_L A B C D E VDD VSS Y
*.PININFO A:I B:I C:I D:I E:I Y:O VDD:B VSS:B
MM9 Y A net024 VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net024 B net023 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net30 D net29 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net29 E VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net023 C net30 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 Y E VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM3 Y D VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 Y C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 Y B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 Y A VSS VSS nmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: O2A1O1Ixp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:08 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    O2A1O1Ixp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT O2A1O1Ixp33_ASAP7_75t_L A1 A2 B C VDD VSS Y
*.PININFO A1:I A2:I B:I C:I Y:O VDD:B VSS:B
MM7 net010 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 Y C net010 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net010 A2 net019 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net019 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 Y C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 net022 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 Y A2 net022 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y A1 net022 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: O2A1O1Ixp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:09 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    O2A1O1Ixp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT O2A1O1Ixp5_ASAP7_75t_L A1 A2 B C VDD VSS Y
*.PININFO A1:I A2:I B:I C:I Y:O VDD:B VSS:B
MM9 Y B net011 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 Y C VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 net011 A2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net011 A1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net03 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net010 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 net03 A2 net010 VDD pmos_lvt w=162.00n l=20n nfin=6
MM5 Y C net03 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA211x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:10 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA211x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA211x2_ASAP7_75t_L A1 A2 B C VDD VSS Y
*.PININFO A1:I A2:I B:I C:I Y:O VDD:B VSS:B
MM0 Y net019 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM39 net019 C VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM38 net019 B VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM37 net019 A2 net20 VDD pmos_lvt w=54.0n l=20n nfin=2
MM36 net20 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 Y net019 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM41 net019 A2 net10 VSS nmos_lvt w=81.0n l=20n nfin=3
MM43 net19 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM40 net019 A1 net10 VSS nmos_lvt w=81.0n l=20n nfin=3
MM42 net10 B net19 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA21x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:12 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA21x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA21x2_ASAP7_75t_L A1 A2 B VDD VSS Y
*.PININFO A1:I A2:I B:I Y:O VDD:B VSS:B
MM3 Y net25 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM2 net25 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net25 A2 net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net27 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 Y net25 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM6 net11 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net25 A2 net11 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 net25 A1 net11 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA221x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:13 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA221x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA221x2_ASAP7_75t_L A1 A2 B1 B2 C VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C:I Y:O VDD:B VSS:B
MM11 net15 B2 net29 VSS nmos_lvt w=162.00n l=20n nfin=6
MM10 net29 A2 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM9 net29 A1 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM6 net15 B1 net29 VSS nmos_lvt w=162.00n l=20n nfin=6
MM12 net014 C net15 VSS nmos_lvt w=162.00n l=20n nfin=6
MM24 Y net014 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM4 net014 C VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM3 net014 B2 net32 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net32 B1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net014 A2 net30 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net30 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 Y net014 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA222x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:14 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA222x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA222x2_ASAP7_75t_L A1 A2 B1 B2 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I Y:O VDD:B VSS:B
MM7 net28 C2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net014 C1 net28 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net014 B1 net29 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net29 B2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net014 A1 net30 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net30 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 Y net014 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM13 net010 C2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net011 B2 net010 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net014 A2 net011 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net010 C1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net011 B1 net010 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net014 A1 net011 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y net014 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA22x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:15 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA22x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA22x2_ASAP7_75t_L A1 A2 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I Y:O VDD:B VSS:B
MM9 Y net033 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM3 net3 B2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net033 A2 net3 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net3 B1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net033 A1 net3 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net13 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net033 A2 net13 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net14 B1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 Y net033 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM10 net033 B2 net14 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA31x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:16 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA31x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA31x2_ASAP7_75t_L A1 A2 A3 B1 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I Y:O VDD:B VSS:B
MM9 Y net20 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM4 net17 B1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net20 A3 net17 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net20 A2 net17 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net20 A1 net17 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 Y net20 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM7 net20 B1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM6 net20 A3 net36 VDD pmos_lvt w=162.00n l=20n nfin=6
MM5 net36 A2 net37 VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 net37 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA331x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:18 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA331x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA331x1_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I Y:O VDD:B VSS:B
MM4 net012 B3 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 VSS net027 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS A1 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS A2 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 VSS A3 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net012 B1 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net031 C1 net027 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net012 B2 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 VDD C1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net033 B1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net063 B2 net033 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 VDD B3 net063 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A3 net26 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net037 A1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net26 A2 net037 VDD pmos_lvt w=81.0n l=20n nfin=3
MM19 VDD net027 Y VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA331x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:19 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA331x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA331x2_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I Y:O VDD:B VSS:B
MM4 net012 B3 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 VSS net027 Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM9 VSS A1 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS A2 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 VSS A3 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net012 B1 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net031 C1 net027 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net012 B2 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 VDD C1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net033 B1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net063 B2 net033 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 VDD B3 net063 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A3 net26 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net037 A1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net26 A2 net037 VDD pmos_lvt w=81.0n l=20n nfin=3
MM19 VDD net027 Y VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA332x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:20 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA332x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA332x1_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I Y:O VDD:B VSS:B
MM4 net059 B3 net060 VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 VSS net027 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS A1 net059 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS A2 net059 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 VSS A3 net059 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net059 B1 net060 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net060 C2 net027 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net060 C1 net027 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net059 B2 net060 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 VDD B3 net080 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A3 net079 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net081 B1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net080 B2 net081 VDD pmos_lvt w=81.0n l=20n nfin=3
MM16 VDD C2 net082 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net079 A2 net078 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net078 A1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM17 net082 C1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM19 VDD net027 Y VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA332x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:21 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA332x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA332x2_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I Y:O VDD:B VSS:B
MM4 net059 B3 net060 VSS nmos_lvt w=81.0n l=20n nfin=3
MM18 VSS net027 Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM9 VSS A1 net059 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS A2 net059 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 VSS A3 net059 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net059 B1 net060 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net060 C2 net027 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net060 C1 net027 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net059 B2 net060 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 VDD B3 net080 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A3 net079 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net081 B1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net080 B2 net081 VDD pmos_lvt w=81.0n l=20n nfin=3
MM16 VDD C2 net082 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net079 A2 net078 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net078 A1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM17 net082 C1 net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM19 VDD net027 Y VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA333x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:22 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA333x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA333x1_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 C3 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I C3:I Y:O VDD:B VSS:B
MM19 VDD net020 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 VDD C3 net040 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net084 A1 net020 VDD pmos_lvt w=81.0n l=20n nfin=3
MM16 net040 C2 net086 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net087 B1 net020 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net041 B2 net087 VDD pmos_lvt w=81.0n l=20n nfin=3
MM17 net086 C1 net020 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A3 net038 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 VDD B3 net041 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net038 A2 net084 VDD pmos_lvt w=81.0n l=20n nfin=3
MM18 VSS net020 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 net068 B3 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net015 A1 net020 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS C2 net068 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS C1 net068 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net068 B1 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 VSS C3 net068 VSS nmos_lvt w=81.0n l=20n nfin=3
MM15 net015 A3 net020 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net068 B2 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net015 A2 net020 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA333x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:24 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA333x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA333x2_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 C3 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I C3:I Y:O VDD:B VSS:B
MM19 VDD net020 Y VDD pmos_lvt w=162.00n l=20n nfin=6
MM13 VDD C3 net040 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net084 A1 net020 VDD pmos_lvt w=81.0n l=20n nfin=3
MM16 net040 C2 net086 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net087 B1 net020 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net041 B2 net087 VDD pmos_lvt w=81.0n l=20n nfin=3
MM17 net086 C1 net020 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A3 net038 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 VDD B3 net041 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net038 A2 net084 VDD pmos_lvt w=81.0n l=20n nfin=3
MM18 VSS net020 Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM4 net068 B3 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net015 A1 net020 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS C2 net068 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS C1 net068 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net068 B1 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 VSS C3 net068 VSS nmos_lvt w=81.0n l=20n nfin=3
MM15 net015 A3 net020 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net068 B2 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net015 A2 net020 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OA33x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:25 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OA33x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OA33x2_ASAP7_75t_L A1 A2 A3 B1 B2 B3 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I Y:O VDD:B VSS:B
MM7 Y net015 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM5 net21 A3 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net015 B3 net21 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 net21 A2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net015 B2 net21 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net21 A1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net015 B1 net21 VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 Y net015 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM13 net34 B1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net33 B2 net34 VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net015 B3 net33 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net35 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 net36 A2 net35 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net015 A3 net36 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI211xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:26 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI211xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI211xp5_ASAP7_75t_L A1 A2 B C VDD VSS Y
*.PININFO A1:I A2:I B:I C:I Y:O VDD:B VSS:B
MM39 Y C VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM38 Y B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM37 Y A2 net20 VDD pmos_lvt w=54.0n l=20n nfin=2
MM36 net20 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM41 Y A2 net10 VSS nmos_lvt w=81.0n l=20n nfin=3
MM43 net19 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM40 Y A1 net10 VSS nmos_lvt w=81.0n l=20n nfin=3
MM42 net10 B net19 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI21x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:27 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI21x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21x1_ASAP7_75t_L A1 A2 B VDD VSS Y
*.PININFO A1:I A2:I B:I Y:O VDD:B VSS:B
MM2 Y B VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM1 Y A2 net27 VDD pmos_lvt w=162.00n l=20n nfin=6
MM0 net27 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 net11 B VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM5 Y A2 net11 VSS nmos_lvt w=162.00n l=20n nfin=6
MM4 Y A1 net11 VSS nmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI21xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:28 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI21xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21xp33_ASAP7_75t_L A1 A2 B VDD VSS Y
*.PININFO A1:I A2:I B:I Y:O VDD:B VSS:B
MM2 Y B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 Y A2 net27 VDD pmos_lvt w=54.0n l=20n nfin=2
MM0 net27 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM6 net11 B VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 Y A2 net11 VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 Y A1 net11 VSS nmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI21xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:30 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI21xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI21xp5_ASAP7_75t_L A1 A2 B VDD VSS Y
*.PININFO A1:I A2:I B:I Y:O VDD:B VSS:B
MM2 Y B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 Y A2 net27 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net27 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net11 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 Y A2 net11 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 Y A1 net11 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI221xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:31 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI221xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI221xp5_ASAP7_75t_L A1 A2 B1 B2 C VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C:I Y:O VDD:B VSS:B
MM11 net15 B2 net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net29 A2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net29 A1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net15 B1 net29 VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 Y C net15 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 Y C VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM3 Y B2 net32 VDD pmos_lvt w=54.0n l=20n nfin=2
MM2 net32 B1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 Y A2 net30 VDD pmos_lvt w=54.0n l=20n nfin=2
MM0 net30 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI222xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:32 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI222xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI222xp33_ASAP7_75t_L A1 A2 B1 B2 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I Y:O VDD:B VSS:B
MM7 net28 C2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 Y C1 net28 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 Y B1 net29 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net29 B2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 Y A1 net30 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net30 A2 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 net010 C2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net011 B2 net010 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 Y A2 net011 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net010 C1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net011 B1 net010 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 Y A1 net011 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI22x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:33 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI22x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22x1_ASAP7_75t_L A1 A2 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I Y:O VDD:B VSS:B
MM3 net3 B2 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 Y A2 net3 VSS nmos_lvt w=162.00n l=20n nfin=6
MM1 net3 B1 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 Y A1 net3 VSS nmos_lvt w=162.00n l=20n nfin=6
MM8 net13 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM11 Y A2 net13 VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 net14 B1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM10 Y B2 net14 VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI22xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:34 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI22xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22xp33_ASAP7_75t_L A1 A2 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I Y:O VDD:B VSS:B
MM3 net3 B2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 Y A2 net3 VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 net3 B1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 Y A1 net3 VSS nmos_lvt w=54.0n l=20n nfin=2
MM8 net13 A1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM11 Y A2 net13 VDD pmos_lvt w=54.0n l=20n nfin=2
MM6 net14 B1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM10 Y B2 net14 VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI22xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:36 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI22xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI22xp5_ASAP7_75t_L A1 A2 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I B1:I B2:I Y:O VDD:B VSS:B
MM3 net3 B2 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 Y A2 net3 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net3 B1 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y A1 net3 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 net13 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 Y A2 net13 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net14 B1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 Y B2 net14 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI311xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:37 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI311xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI311xp33_ASAP7_75t_L A1 A2 A3 B1 C1 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I C1:I Y:O VDD:B VSS:B
MM16 net037 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 Y C1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM5 Y B1 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM3 Y A1 net30 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net30 A2 net037 VDD pmos_lvt w=81.0n l=20n nfin=3
MM22 VSS A3 net011 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 VSS A1 net011 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net022 C1 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net011 B1 net022 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS A2 net011 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI31xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:38 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI31xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI31xp33_ASAP7_75t_L A1 A2 A3 B VDD VSS Y
*.PININFO A1:I A2:I A3:I B:I Y:O VDD:B VSS:B
MM1 net039 A2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM11 Y B net039 VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 net039 A1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM8 net039 A3 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM15 Y B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM14 net047 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 net048 A2 net047 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 Y A3 net048 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI31xp67_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:39 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI31xp67_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI31xp67_ASAP7_75t_L A1 A2 A3 B VDD VSS Y
*.PININFO A1:I A2:I A3:I B:I Y:O VDD:B VSS:B
MM1 net17 A2 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM11 Y B net17 VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 net17 A1 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM8 net17 A3 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM15 Y B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM14 net22 A1 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM13 net23 A2 net22 VDD pmos_lvt w=162.00n l=20n nfin=6
MM12 Y A3 net23 VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI321xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:40 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI321xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI321xp33_ASAP7_75t_L A1 A2 A3 B1 B2 C VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I C:I Y:O VDD:B VSS:B
MM8 net013 B2 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net012 C net013 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net013 B1 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 VSS A3 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 VSS A2 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 VSS A1 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net031 B2 Y VDD pmos_lvt w=54.0n l=20n nfin=2
MM0 VDD C Y VDD pmos_lvt w=54.0n l=20n nfin=2
MM5 VDD B1 net031 VDD pmos_lvt w=54.0n l=20n nfin=2
MM4 VDD A3 net032 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net29 A1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net032 A2 net29 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI322xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:41 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI322xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI322xp33_ASAP7_75t_L A1 A2 A3 B1 B2 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I C1:I C2:I Y:O VDD:B VSS:B
MM16 net037 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net28 C2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM6 Y C1 net28 VDD pmos_lvt w=54.0n l=20n nfin=2
MM5 Y B1 net29 VDD pmos_lvt w=54.0n l=20n nfin=2
MM4 net29 B2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM3 Y A3 net30 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net30 A2 net037 VDD pmos_lvt w=81.0n l=20n nfin=3
MM22 net026 A3 net022 VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 net022 C1 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net026 A2 net022 VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 VSS B2 net026 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net022 C2 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 net026 A1 net022 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS B1 net026 VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI32xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:43 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI32xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI32xp33_ASAP7_75t_L A1 A2 A3 B1 B2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I Y:O VDD:B VSS:B
MM21 net019 A3 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 Y B2 net019 VSS nmos_lvt w=54.0n l=20n nfin=2
MM5 Y B1 net019 VSS nmos_lvt w=54.0n l=20n nfin=2
MM15 net019 A2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM14 net019 A1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 net025 A3 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net24 A2 net025 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 Y A1 net24 VDD pmos_lvt w=81.0n l=20n nfin=3
MM18 Y B1 net027 VDD pmos_lvt w=54.0n l=20n nfin=2
MM13 net027 B2 VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI331xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:44 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI331xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI331xp33_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I Y:O VDD:B VSS:B
MM4 net012 B3 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS A1 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS A2 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 VSS A3 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net012 B1 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net031 C1 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net012 B2 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 VDD C1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net033 B1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net063 B2 net033 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 VDD B3 net063 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A3 net26 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net037 A1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net26 A2 net037 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI332xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:45 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI332xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI332xp33_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I Y:O VDD:B VSS:B
MM9 VSS A1 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS A2 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 VSS A3 net012 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net012 B1 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net031 C1 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net012 B2 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 net012 B3 net031 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net031 C2 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 net035 C1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM16 VDD C2 net035 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net033 B1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net063 B2 net033 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 VDD B3 net063 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A3 net26 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net037 A1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net26 A2 net037 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI333xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:46 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI333xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI333xp33_ASAP7_75t_L A1 A2 A3 B1 B2 B3 C1 C2 C3 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I C1:I C2:I C3:I Y:O VDD:B VSS:B
MM13 VDD C3 net040 VDD pmos_lvt w=81.0n l=20n nfin=3
MM14 net084 A1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM16 net040 C2 net086 VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 net087 B1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net041 B2 net087 VDD pmos_lvt w=81.0n l=20n nfin=3
MM17 net086 C1 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A3 net038 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 VDD B3 net041 VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net038 A2 net084 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net068 B3 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net015 A1 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 VSS C2 net068 VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS C1 net068 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 net068 B1 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 VSS C3 net068 VSS nmos_lvt w=81.0n l=20n nfin=3
MM15 net015 A3 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net068 B2 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net015 A2 Y VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OAI33xp33_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:47 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OAI33xp33_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OAI33xp33_ASAP7_75t_L A1 A2 A3 B1 B2 B3 VDD VSS Y
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I Y:O VDD:B VSS:B
MM33 Y B1 net028 VSS nmos_lvt w=54.0n l=20n nfin=2
MM35 net028 A3 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM32 Y B2 net028 VSS nmos_lvt w=54.0n l=20n nfin=2
MM38 net028 A2 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM31 Y B3 net028 VSS nmos_lvt w=54.0n l=20n nfin=2
MM37 net028 A1 VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM44 net052 B1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM45 net050 B2 net052 VDD pmos_lvt w=81.0n l=20n nfin=3
MM48 Y B3 net050 VDD pmos_lvt w=81.0n l=20n nfin=3
MM39 net018 A1 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM46 net54 A2 net018 VDD pmos_lvt w=81.0n l=20n nfin=3
MM47 Y A3 net54 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OR2x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:49 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OR2x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OR2x2_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM5 VSS net7 Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM1 VSS B net7 VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 VSS A net7 VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 VDD net7 Y VDD pmos_lvt w=162.00n l=20n nfin=6
MM4 net15 B net7 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A net15 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OR2x4_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:50 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OR2x4_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OR2x4_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM5 VSS net7 Y VSS nmos_lvt w=324.00n l=20n nfin=12
MM1 VSS B net7 VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 VSS A net7 VSS nmos_lvt w=54.0n l=20n nfin=2
MM0 VDD net7 Y VDD pmos_lvt w=324.00n l=20n nfin=12
MM4 net15 B net7 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A net15 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OR2x6_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:51 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OR2x6_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OR2x6_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM5 VSS net7 Y VSS nmos_lvt w=486.00n l=20n nfin=18
MM1 VSS B net7 VSS nmos_lvt w=108.00n l=20n nfin=4
MM2 VSS A net7 VSS nmos_lvt w=108.00n l=20n nfin=4
MM0 VDD net7 Y VDD pmos_lvt w=486.00n l=20n nfin=18
MM4 net15 B net7 VDD pmos_lvt w=162.00n l=20n nfin=6
MM3 VDD A net15 VDD pmos_lvt w=162.00n l=20n nfin=6
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OR3x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:53 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OR3x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OR3x1_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM1 Y net61 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 net61 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 net61 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net61 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y net61 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM8 net66 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net67 B net66 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net61 A net67 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OR3x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:54 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OR3x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OR3x2_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM1 Y net61 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM14 net61 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 net61 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net61 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y net61 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM8 net66 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net67 B net66 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net61 A net67 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OR3x4_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:55 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OR3x4_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OR3x4_ASAP7_75t_L A B C VDD VSS Y
*.PININFO A:I B:I C:I Y:O VDD:B VSS:B
MM1 Y net61 VSS VSS nmos_lvt w=324.00n l=20n nfin=12
MM14 net61 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 net61 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 net61 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 Y net61 VDD VDD pmos_lvt w=324.00n l=20n nfin=12
MM8 net66 C VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 net67 B net66 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 net61 A net67 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OR4x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:56 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OR4x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OR4x1_ASAP7_75t_L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MM9 Y net12 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net12 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net12 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net12 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net12 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 Y net12 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 net12 A pd1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 pd1 B pd2 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 pd2 C pd3 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 pd3 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OR4x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:57 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OR4x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OR4x2_ASAP7_75t_L A B C D VDD VSS Y
*.PININFO A:I B:I C:I D:I Y:O VDD:B VSS:B
MM9 Y net12 VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM3 net12 D VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net12 C VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 net12 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net12 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 Y net12 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM7 net12 A pd1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 pd1 B pd2 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 pd2 C pd3 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 pd3 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OR5x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:52:59 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OR5x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OR5x1_ASAP7_75t_L A B C D E VDD VSS Y
*.PININFO A:I B:I C:I D:I E:I Y:O VDD:B VSS:B
MM9 VSS E net024 VSS nmos_lvt w=54.0n l=20n nfin=2
MM8 VSS D net024 VSS nmos_lvt w=54.0n l=20n nfin=2
MM7 VSS C net024 VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 VSS B net024 VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 VSS net024 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 VSS A net024 VSS nmos_lvt w=54.0n l=20n nfin=2
MM11 VDD net024 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 VDD E net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net027 D net29 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net30 B net023 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net023 A net024 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net29 C net30 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: OR5x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:00 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    OR5x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT OR5x2_ASAP7_75t_L A B C D E VDD VSS Y
*.PININFO A:I B:I C:I D:I E:I Y:O VDD:B VSS:B
MM9 VSS E net024 VSS nmos_lvt w=54.0n l=20n nfin=2
MM8 VSS D net024 VSS nmos_lvt w=54.0n l=20n nfin=2
MM7 VSS C net024 VSS nmos_lvt w=54.0n l=20n nfin=2
MM2 VSS B net024 VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 VSS net024 Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM10 VSS A net024 VSS nmos_lvt w=54.0n l=20n nfin=2
MM11 VDD net024 Y VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 VDD E net027 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 net027 D net29 VDD pmos_lvt w=81.0n l=20n nfin=3
MM4 net30 B net023 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net023 A net024 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net29 C net30 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: SDFHx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:01 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    SDFHx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT SDFHx1_ASAP7_75t_L CLK D QN SE SI VDD VSS
*.PININFO CLK:I D:I SE:I SI:I QN:O VDD:B VSS:B
MM28 net0166 SEn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 net0167 SE VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM29 net0118 D net0166 VSS nmos_lvt w=81.0n l=20n nfin=3
MM30 SEn SE VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkb SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM17 SH clkn pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 QN SH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn net0118 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net0118 SI net0167 VSS nmos_lvt w=81.0n l=20n nfin=3
MM27 net0120 SI net0141 VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM3 net0120 SE net0141 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 MH clkb net0120 VDD pmos_lvt w=81.0n l=20n nfin=3
MM31 SEn SE VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM2 net0141 SEn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkn SH VDD pmos_lvt w=27n l=20n nfin=1
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkb pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM25 QN SH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM26 net0141 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: SDFHx2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:02 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    SDFHx2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT SDFHx2_ASAP7_75t_L CLK D QN SE SI VDD VSS
*.PININFO CLK:I D:I SE:I SI:I QN:O VDD:B VSS:B
MM5 net0118 SI net0166 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn net0118 VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 QN SH VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM17 SH clkn pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkb SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM30 SEn SE VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM29 net0118 D net0167 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM0 net0166 SE VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM28 net0167 SEn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkb pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM26 net0141 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 QN SH VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkn SH VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM2 net0141 SEn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM31 SEn SE VDD VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH clkb net0120 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net0120 SE net0141 VDD pmos_lvt w=81.0n l=20n nfin=3
MM27 net0120 SI net0141 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: SDFHx3_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:03 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    SDFHx3_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT SDFHx3_ASAP7_75t_L CLK D QN SE SI VDD VSS
*.PININFO CLK:I D:I SE:I SI:I QN:O VDD:B VSS:B
MM5 net13 SI net134 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn net13 VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 QN SH VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM17 SH clkn pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkb SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkb pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM30 SEn SE VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM29 net13 D net137 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM0 net134 SE VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM28 net137 SEn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM2 net62 SEn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM31 SEn SE VDD VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH clkb net15 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 net15 SE net62 VDD pmos_lvt w=81.0n l=20n nfin=3
MM27 net15 SI net62 VDD pmos_lvt w=81.0n l=20n nfin=3
MM26 net62 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 QN SH VDD VDD pmos_lvt w=243.00n l=20n nfin=9
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkb pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkn SH VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkn pd2 VDD pmos_lvt w=27n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: SDFHx4_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:05 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    SDFHx4_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT SDFHx4_ASAP7_75t_L CLK D QN SE SI VDD VSS
*.PININFO CLK:I D:I SE:I SI:I QN:O VDD:B VSS:B
MM30 SEn SE VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM29 pd1 D net066 VSS nmos_lvt w=81.0n l=20n nfin=3
MM28 net066 SEn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM27 net067 SE VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkn pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 pd1 SI net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 pd3 MS VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 MH clkb pd3 VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 MS clkb SH VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 SS SH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 pd5 SS VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 SH clkn pd5 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM23 clkb clkn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 QN SH VSS VSS nmos_lvt w=324.00n l=20n nfin=12
MM31 SEn SE VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM26 net54 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 pu1 SI net54 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net54 SEn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 SE net54 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 MH clkb pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 MS MH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 MH clkn pd2 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 pd2 MS VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 MS clkn SH VDD pmos_lvt w=81.0n l=20n nfin=3
MM15 SS SH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM18 SH clkb pd4 VDD pmos_lvt w=81.0n l=20n nfin=3
MM19 pd4 SS VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM22 clkb clkn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 QN SH VDD VDD pmos_lvt w=324.00n l=20n nfin=12
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: SDFLx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:06 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    SDFLx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT SDFLx1_ASAP7_75t_L CLK D QN SE SI VDD VSS
*.PININFO CLK:I D:I SE:I SI:I QN:O VDD:B VSS:B
MM24 QN SH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM17 SH clkb pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkn SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM5 pd1 SE net0168 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 SEn SE VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM26 net0168 SI VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM32 pd1 D net0167 VSS nmos_lvt w=81.0n l=20n nfin=3
MM29 net0167 SEn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 MS clkb SH VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 SI net0144 VDD pmos_lvt w=81.0n l=20n nfin=3
MM31 pu1 SE net0144 VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 MH clkb pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM2 SEn SE VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM27 net0144 SEn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM30 net0144 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM25 QN SH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkn pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: SDFLx2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:07 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    SDFLx2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT SDFLx2_ASAP7_75t_L CLK D QN SE SI VDD VSS
*.PININFO CLK:I D:I SE:I SI:I QN:O VDD:B VSS:B
MM29 net0168 SEn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM32 pd1 D net0168 VSS nmos_lvt w=81.0n l=20n nfin=3
MM26 net0167 SI VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 SEn SE VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 pd1 SE net0167 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkn SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM17 SH clkb pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 QN SH VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkb pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkn pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM25 QN SH VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM13 MS clkb SH VDD pmos_lvt w=27n l=20n nfin=1
MM30 net0144 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM27 net0144 SEn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 SEn SE VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM31 pu1 SE net0144 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 SI net0144 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: SDFLx3_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:08 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    SDFLx3_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT SDFLx3_ASAP7_75t_L CLK D QN SE SI VDD VSS
*.PININFO CLK:I D:I SE:I SI:I QN:O VDD:B VSS:B
MM29 net061 SEn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM32 pd1 D net061 VSS nmos_lvt w=81.0n l=20n nfin=3
MM26 net062 SI VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 SEn SE VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 pd1 SE net062 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM8 pd3 MS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM9 MH clkn pd3 VSS nmos_lvt w=27.0n l=20n nfin=1
MM12 MS clkn SH VSS nmos_lvt w=27.0n l=20n nfin=1
MM14 SS SH VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM16 pd5 SS VSS VSS nmos_lvt w=27.0n l=20n nfin=1
MM17 SH clkb pd5 VSS nmos_lvt w=27.0n l=20n nfin=1
MM20 clkn CLK VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM23 clkb clkn VSS VSS nmos_lvt w=54.0n l=20n nfin=2
MM24 QN SH VSS VSS nmos_lvt w=243.00n l=20n nfin=9
MM30 net063 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM27 net063 SEn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 SEn SE VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM31 pu1 SE net063 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 SI net063 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 MS MH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM10 MH clkb pd2 VDD pmos_lvt w=27n l=20n nfin=1
MM11 pd2 MS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM13 MS clkb SH VDD pmos_lvt w=27n l=20n nfin=1
MM15 SS SH VDD VDD pmos_lvt w=27n l=20n nfin=1
MM18 SH clkn pd4 VDD pmos_lvt w=27n l=20n nfin=1
MM19 pd4 SS VDD VDD pmos_lvt w=27n l=20n nfin=1
MM21 clkn CLK VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM22 clkb clkn VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM25 QN SH VDD VDD pmos_lvt w=243.00n l=20n nfin=9
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: SDFLx4_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:09 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    SDFLx4_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT SDFLx4_ASAP7_75t_L CLK D QN SE SI VDD VSS
*.PININFO CLK:I D:I SE:I SI:I QN:O VDD:B VSS:B
MM30 SEn SE VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM29 pd1 D net066 VSS nmos_lvt w=81.0n l=20n nfin=3
MM28 net066 SEn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM27 net067 SE VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 MH clkb pd1 VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 pd1 SI net067 VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 MS MH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM8 pd3 MS VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 MH clkn pd3 VSS nmos_lvt w=81.0n l=20n nfin=3
MM12 MS clkn SH VSS nmos_lvt w=81.0n l=20n nfin=3
MM14 SS SH VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM16 pd5 SS VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM17 SH clkb pd5 VSS nmos_lvt w=81.0n l=20n nfin=3
MM20 clkn CLK VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM23 clkb clkn VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM24 QN SH VSS VSS nmos_lvt w=324.00n l=20n nfin=12
MM31 SEn SE VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM26 net54 D VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 pu1 SI net54 VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net54 SEn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 pu1 SE net54 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 MH clkn pu1 VDD pmos_lvt w=81.0n l=20n nfin=3
MM7 MS MH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 MH clkb pd2 VDD pmos_lvt w=81.0n l=20n nfin=3
MM11 pd2 MS VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM13 MS clkb SH VDD pmos_lvt w=81.0n l=20n nfin=3
MM15 SS SH VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM18 SH clkn pd4 VDD pmos_lvt w=81.0n l=20n nfin=3
MM19 pd4 SS VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM21 clkn CLK VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM22 clkb clkn VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM25 QN SH VDD VDD pmos_lvt w=324.00n l=20n nfin=12
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: TIEHIx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:10 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    TIEHIx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT TIEHIx1_ASAP7_75t_L H VDD VSS
*.PININFO H:O VDD:B VSS:B
MM1 H net7 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net7 H VSS VSS nmos_lvt w=27.0n l=20n nfin=1
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: TIELOx1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:12 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    TIELOx1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT TIELOx1_ASAP7_75t_L L VDD VSS
*.PININFO L:O VDD:B VSS:B
MM1 net9 L VDD VDD pmos_lvt w=27.0n l=20n nfin=1
MM2 L net9 VSS VSS nmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: XNOR2x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:13 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    XNOR2x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2x1_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM4 net015 A VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM5 net015 B VSS VSS nmos_lvt w=162.00n l=20n nfin=6
MM6 Y net29 net015 VSS nmos_lvt w=162.00n l=20n nfin=6
MM2 net29 B net43 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net43 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net041 A VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM10 Y B net041 VDD pmos_lvt w=162.00n l=20n nfin=6
MM9 Y net29 VDD VDD pmos_lvt w=162.00n l=20n nfin=6
MM0 net29 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net29 B VDD VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: XNOR2x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:14 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    XNOR2x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2x2_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM11 VSS A net047 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net047 B xor VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS net036 xor VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 VSS xor Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 VSS A net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 VSS B net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 VDD A net019 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 VDD B net019 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net019 net036 xor VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 VDD xor Y VDD pmos_lvt w=162.00n l=20n nfin=6
MM2 net048 B net036 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A net048 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: XNOR2xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:15 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    XNOR2xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT XNOR2xp5_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM4 net015 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net015 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM6 Y net29 net015 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net29 B net43 VSS nmos_lvt w=81.0n l=20n nfin=3
MM3 net43 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net041 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM10 Y B net041 VDD pmos_lvt w=81.0n l=20n nfin=3
MM9 Y net29 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net29 A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM1 net29 B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: XOR2x1_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:16 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    XOR2x1_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2x1_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM11 VSS A net047 VSS nmos_lvt w=162.00n l=20n nfin=6
MM10 net047 B Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM9 VSS net036 Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM0 VSS A net036 VSS nmos_lvt w=81.0n l=20n nfin=3
MM1 VSS B net036 VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 VDD A net019 VDD pmos_lvt w=162.00n l=20n nfin=6
MM5 VDD B net019 VDD pmos_lvt w=162.00n l=20n nfin=6
MM6 net019 net036 Y VDD pmos_lvt w=162.00n l=20n nfin=6
MM2 net048 B net036 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A net048 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: XOR2x2_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:18 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    XOR2x2_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2x2_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM6 xor net045 net049 VSS nmos_lvt w=81.0n l=20n nfin=3
MM2 net045 B net060 VSS nmos_lvt w=81.0n l=20n nfin=3
MM13 VSS xor Y VSS nmos_lvt w=162.00n l=20n nfin=6
MM3 net060 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM4 net049 A VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM5 net049 B VSS VSS nmos_lvt w=81.0n l=20n nfin=3
MM11 net059 A VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM0 net045 A VDD VDD pmos_lvt w=54.0n l=20n nfin=2
MM9 xor net045 VDD VDD pmos_lvt w=81.0n l=20n nfin=3
MM12 VDD xor Y VDD pmos_lvt w=162.00n l=20n nfin=6
MM10 xor B net059 VDD pmos_lvt w=81.0n l=20n nfin=3
MM1 net045 B VDD VDD pmos_lvt w=54.0n l=20n nfin=2
.ENDS

************************************************************************
* auCdl Netlist:
* 
* Library Name:  asap7sc7p5t_24_L
* Top Cell Name: XOR2xp5_ASAP7_75t_L
* View Name:     schematic
* Netlisted on:  Sep  8 16:53:19 2017
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: asap7sc7p5t_24_L
* Cell Name:    XOR2xp5_ASAP7_75t_L
* View Name:    schematic
************************************************************************

.SUBCKT XOR2xp5_ASAP7_75t_L A B VDD VSS Y
*.PININFO A:I B:I Y:O VDD:B VSS:B
MM11 VSS A net047 VSS nmos_lvt w=81.0n l=20n nfin=3
MM10 net047 B Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM9 VSS net036 Y VSS nmos_lvt w=81.0n l=20n nfin=3
MM0 VSS A net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MM1 VSS B net036 VSS nmos_lvt w=54.0n l=20n nfin=2
MM4 VDD A net019 VDD pmos_lvt w=81.0n l=20n nfin=3
MM5 VDD B net019 VDD pmos_lvt w=81.0n l=20n nfin=3
MM6 net019 net036 Y VDD pmos_lvt w=81.0n l=20n nfin=3
MM2 net048 B net036 VDD pmos_lvt w=81.0n l=20n nfin=3
MM3 VDD A net048 VDD pmos_lvt w=81.0n l=20n nfin=3
.ENDS

