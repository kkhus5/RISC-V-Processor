`include "const.vh"

module Riscv151(
    input clk,
    input reset,

    // Memory system ports
    output [31:0] dcache_addr,
    output [31:0] icache_addr,
    output [3:0] dcache_we,
    output dcache_re,
    output icache_re,
    output [31:0] dcache_din,
    input [31:0] dcache_dout,
    input [31:0] icache_dout,
    input stall,
    output [31:0] csr

);

    // TODO: Your code
    // Please use REGFILE_1W2R for your register file
    // (two async read ports, 1 sync write port)
    // Please use REGISTER* modules for all sequential logic


endmodule
