* File: NAND2x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:37:58 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND2x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND2x1_ASAP7_75t_R.pex.sp.pex"
* File: NAND2x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:37:58 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND2X1_ASAP7_75T_R%A 2 8 11 13 29 VSS
c15 29 VSS 0.0177504f $X=0.07 $Y=0.136
c16 11 VSS 0.00986222f $X=0.135 $Y=0.1345
c17 8 VSS 0.0631368f $X=0.135 $Y=0.0675
c18 2 VSS 0.0689981f $X=0.081 $Y=0.0675
r19 26 29 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.07 $Y=0.135 $X2=0.07
+ $Y2=0.135
r20 11 13 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1345 $X2=0.135 $Y2=0.2025
r21 8 11 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1345
r22 5 11 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1345 $X2=0.135 $Y2=0.1345
r23 5 26 9.56522 $w=2.3e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1345 $X2=0.07 $Y2=0.1345
r24 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.1345
.ends

.subckt PM_NAND2X1_ASAP7_75T_R%B 2 7 10 13 18 23 VSS
c21 25 VSS 5.59368e-20 $X=0.243 $Y=0.148
c22 23 VSS 0.00121422f $X=0.24 $Y=0.152
c23 18 VSS 9.98653e-19 $X=0.243 $Y=0.135
c24 13 VSS 0.00433435f $X=0.243 $Y=0.135
c25 10 VSS 0.0680685f $X=0.243 $Y=0.0675
c26 2 VSS 0.0623886f $X=0.189 $Y=0.0675
r27 24 25 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.144 $X2=0.243 $Y2=0.148
r28 23 25 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.152 $X2=0.243 $Y2=0.148
r29 18 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.144
r30 13 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r31 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r32 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r33 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r34 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_NAND2X1_ASAP7_75T_R%5 1 6 7 11 14 17 18 24 25 28 29 30 31 VSS
c21 31 VSS 0.00263922f $X=0.236 $Y=0.036
c22 30 VSS 0.0123864f $X=0.202 $Y=0.036
c23 29 VSS 0.00289079f $X=0.27 $Y=0.036
c24 28 VSS 0.0049699f $X=0.27 $Y=0.036
c25 26 VSS 9.61037e-19 $X=0.094 $Y=0.036
c26 25 VSS 0.00270713f $X=0.084 $Y=0.036
c27 24 VSS 0.00659293f $X=0.162 $Y=0.036
c28 18 VSS 0.00651324f $X=0.054 $Y=0.036
c29 17 VSS 0.00190113f $X=0.054 $Y=0.036
c30 14 VSS 3.4551e-19 $X=0.268 $Y=0.0675
c31 6 VSS 6.15054e-19 $X=0.179 $Y=0.0675
c32 1 VSS 4.64427e-19 $X=0.071 $Y=0.0675
r33 30 31 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.036 $X2=0.236 $Y2=0.036
r34 28 31 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.236 $Y2=0.036
r35 28 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r36 25 26 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.084
+ $Y=0.036 $X2=0.094 $Y2=0.036
r37 23 30 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.202 $Y2=0.036
r38 23 26 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.094 $Y2=0.036
r39 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r40 17 25 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.084 $Y2=0.036
r41 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r42 14 29 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r43 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.268 $Y2=0.0675
r44 10 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r45 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r46 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r47 4 18 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r48 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends

.subckt PM_NAND2X1_ASAP7_75T_R%Y 1 2 5 6 9 11 14 24 26 27 30 35 36 40 42 VSS
c29 44 VSS 5.3979e-19 $X=0.297 $Y=0.216
c30 42 VSS 9.39445e-19 $X=0.297 $Y=0.122
c31 41 VSS 8.85605e-19 $X=0.297 $Y=0.099
c32 40 VSS 0.00369303f $X=0.298 $Y=0.145
c33 38 VSS 5.09802e-19 $X=0.297 $Y=0.225
c34 36 VSS 3.28196e-19 $X=0.284 $Y=0.072
c35 35 VSS 8.46035e-21 $X=0.252 $Y=0.072
c36 30 VSS 3.5796e-19 $X=0.216 $Y=0.072
c37 28 VSS 0.00199089f $X=0.288 $Y=0.072
c38 27 VSS 0.00187504f $X=0.27 $Y=0.234
c39 26 VSS 0.0029456f $X=0.252 $Y=0.234
c40 25 VSS 0.00110824f $X=0.215 $Y=0.234
c41 24 VSS 0.0128273f $X=0.202 $Y=0.234
c42 16 VSS 0.00522611f $X=0.288 $Y=0.234
c43 14 VSS 0.00739362f $X=0.214 $Y=0.2025
c44 9 VSS 0.00719461f $X=0.11 $Y=0.2025
c45 6 VSS 4.6121e-19 $X=0.125 $Y=0.2025
c46 5 VSS 0.00299094f $X=0.216 $Y=0.0675
c47 1 VSS 6.09911e-19 $X=0.233 $Y=0.0675
r48 43 44 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.207 $X2=0.297 $Y2=0.216
r49 41 42 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.099 $X2=0.297 $Y2=0.122
r50 40 43 4.20988 $w=1.8e-08 $l=6.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.145 $X2=0.297 $Y2=0.207
r51 40 42 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.145 $X2=0.297 $Y2=0.122
r52 38 44 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.216
r53 37 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.081 $X2=0.297 $Y2=0.099
r54 35 36 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.072 $X2=0.284 $Y2=0.072
r55 30 35 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.072 $X2=0.252 $Y2=0.072
r56 28 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.072 $X2=0.297 $Y2=0.081
r57 28 36 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.284 $Y2=0.072
r58 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.27 $Y2=0.234
r59 24 25 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.234 $X2=0.215 $Y2=0.234
r60 22 26 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.252 $Y2=0.234
r61 22 25 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.215 $Y2=0.234
r62 18 24 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.202 $Y2=0.234
r63 16 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.234 $X2=0.297 $Y2=0.225
r64 16 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.27 $Y2=0.234
r65 14 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r66 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.214 $Y2=0.2025
r67 9 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r68 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.11 $Y2=0.2025
r69 5 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072 $X2=0.216
+ $Y2=0.072
r70 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r71 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./NAND2x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND2x1_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 VSS N_A_M0_g N_5_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 VSS N_A_M1_g N_5_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_B_M2_g N_5_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_Y_M3_d N_B_M3_g N_5_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 VDD N_A_M4_g N_Y_M4_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M5 N_Y_M5_d N_B_M5_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
*
* 
* .include "NAND2x1_ASAP7_75t_R.pex.sp.NAND2X1_ASAP7_75T_R.pxi"
* BEGIN of "./NAND2x1_ASAP7_75t_R.pex.sp.NAND2X1_ASAP7_75T_R.pxi"
* File: NAND2x1_ASAP7_75t_R.pex.sp.NAND2X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:37:58 2017
* 
x_PM_NAND2X1_ASAP7_75T_R%A N_A_M0_g N_A_M1_g N_A_c_4_p N_A_M4_g A VSS
+ PM_NAND2X1_ASAP7_75T_R%A
x_PM_NAND2X1_ASAP7_75T_R%B N_B_M2_g N_B_M5_g N_B_M3_g N_B_c_19_n N_B_c_21_p B
+ VSS PM_NAND2X1_ASAP7_75T_R%B
x_PM_NAND2X1_ASAP7_75T_R%5 N_5_M0_s N_5_M2_s N_5_M1_s N_5_M3_s N_5_c_55_p
+ N_5_c_37_n N_5_c_38_n N_5_c_47_p N_5_c_39_n N_5_c_43_n N_5_c_44_n N_5_c_42_n
+ N_5_c_49_p VSS PM_NAND2X1_ASAP7_75T_R%5
x_PM_NAND2X1_ASAP7_75T_R%Y N_Y_M3_d N_Y_M2_d N_Y_c_64_n N_Y_M4_s N_Y_c_58_n
+ N_Y_M5_d N_Y_c_66_n N_Y_c_60_n N_Y_c_70_n N_Y_c_80_n N_Y_c_81_n N_Y_c_72_n
+ N_Y_c_84_n Y N_Y_c_75_n VSS PM_NAND2X1_ASAP7_75T_R%Y
cc_1 N_A_M0_g N_B_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_A_M1_g N_B_M2_g 0.0032073f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A_M1_g N_B_M3_g 2.66145e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_4 N_A_c_4_p N_B_c_19_n 0.00220839f $X=0.135 $Y=0.1345 $X2=0.243 $Y2=0.135
cc_5 A N_5_c_37_n 0.00116786f $X=0.07 $Y=0.136 $X2=0.243 $Y2=0.135
cc_6 A N_5_c_38_n 0.00222573f $X=0.07 $Y=0.136 $X2=0.243 $Y2=0.135
cc_7 N_A_M0_g N_5_c_39_n 2.7229e-19 $X=0.081 $Y=0.0675 $X2=0.243 $Y2=0.148
cc_8 N_A_c_4_p N_5_c_39_n 0.0010215f $X=0.135 $Y=0.1345 $X2=0.243 $Y2=0.148
cc_9 A N_5_c_39_n 2.11212e-19 $X=0.07 $Y=0.136 $X2=0.243 $Y2=0.148
cc_10 N_A_M1_g N_5_c_42_n 4.56095e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_11 N_A_c_4_p N_Y_c_58_n 8.01479e-19 $X=0.135 $Y=0.1345 $X2=0.243 $Y2=0.0675
cc_12 A N_Y_c_58_n 0.00166117f $X=0.07 $Y=0.136 $X2=0.243 $Y2=0.0675
cc_13 N_A_M1_g N_Y_c_60_n 4.58656e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.144
cc_14 N_A_c_4_p N_Y_c_60_n 5.29557e-19 $X=0.135 $Y=0.1345 $X2=0.243 $Y2=0.144
cc_15 A N_Y_c_60_n 8.40589e-19 $X=0.07 $Y=0.136 $X2=0.243 $Y2=0.144
cc_16 N_B_M3_g N_5_c_43_n 2.08515e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_17 N_B_c_21_p N_5_c_44_n 2.73699e-19 $X=0.243 $Y=0.135 $X2=0.07 $Y2=0.136
cc_18 N_B_M2_g N_5_c_42_n 4.58656e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_19 N_B_c_19_n N_5_c_42_n 2.67739e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_20 N_B_c_19_n N_Y_M3_d 3.78404e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_21 N_B_c_19_n N_Y_c_64_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.1345
cc_22 N_B_c_21_p N_Y_c_64_n 8.82763e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.1345
cc_23 N_B_c_19_n N_Y_c_66_n 8.00061e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_24 B N_Y_c_66_n 0.00319197f $X=0.24 $Y=0.152 $X2=0 $Y2=0
cc_25 N_B_M2_g N_Y_c_60_n 4.58656e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_B_c_19_n N_Y_c_60_n 3.87029e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_27 N_B_M3_g N_Y_c_70_n 2.34993e-19 $X=0.243 $Y=0.0675 $X2=0.07 $Y2=0.135
cc_28 B N_Y_c_70_n 0.00371828f $X=0.24 $Y=0.152 $X2=0.07 $Y2=0.135
cc_29 N_B_M3_g N_Y_c_72_n 2.52885e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_B_c_21_p N_Y_c_72_n 0.00371264f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 N_B_c_21_p Y 0.00257364f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_32 N_B_c_21_p N_Y_c_75_n 0.00257364f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_33 N_5_c_47_p N_Y_c_64_n 0.00339108f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.1345
cc_34 N_5_c_44_n N_Y_c_64_n 0.00384465f $X=0.27 $Y=0.036 $X2=0.081 $Y2=0.1345
cc_35 N_5_c_49_p N_Y_c_64_n 0.00253713f $X=0.236 $Y=0.036 $X2=0.081 $Y2=0.1345
cc_36 N_5_c_42_n N_Y_c_60_n 2.48138e-19 $X=0.202 $Y=0.036 $X2=0 $Y2=0
cc_37 N_5_c_43_n N_Y_c_80_n 2.48138e-19 $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_38 N_5_c_47_p N_Y_c_81_n 5.19937e-19 $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_39 N_5_c_49_p N_Y_c_81_n 0.00351928f $X=0.236 $Y=0.036 $X2=0 $Y2=0
cc_40 N_5_c_43_n N_Y_c_72_n 0.00351928f $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_41 N_5_c_55_p N_Y_c_84_n 2.53396e-19 $X=0.268 $Y=0.0675 $X2=0.07 $Y2=0.1345
cc_42 N_5_c_44_n N_Y_c_84_n 0.00260156f $X=0.27 $Y=0.036 $X2=0.07 $Y2=0.1345
cc_43 N_5_c_44_n N_Y_c_75_n 2.86097e-19 $X=0.27 $Y=0.036 $X2=0 $Y2=0

* END of "./NAND2x1_ASAP7_75t_R.pex.sp.NAND2X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND2x1p5_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:38:20 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND2x1p5_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND2x1p5_ASAP7_75t_R.pex.sp.pex"
* File: NAND2x1p5_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:38:20 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND2X1P5_ASAP7_75T_R%A 2 8 13 16 19 21 37 VSS
c22 37 VSS 0.0246493f $X=0.07 $Y=0.136
c23 19 VSS 0.012275f $X=0.189 $Y=0.1345
c24 16 VSS 0.0622543f $X=0.189 $Y=0.0675
c25 8 VSS 0.0638575f $X=0.135 $Y=0.0675
c26 2 VSS 0.067082f $X=0.081 $Y=0.0675
r27 34 37 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.07 $Y=0.135 $X2=0.07
+ $Y2=0.135
r28 19 21 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1345 $X2=0.189 $Y2=0.216
r29 16 19 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.1345
r30 11 19 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.1345 $X2=0.189 $Y2=0.1345
r31 11 13 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1345 $X2=0.135 $Y2=0.2025
r32 8 11 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1345
r33 5 11 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1345 $X2=0.135 $Y2=0.1345
r34 5 34 9.56522 $w=2.3e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1345 $X2=0.07 $Y2=0.1345
r35 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.1345
.ends

.subckt PM_NAND2X1P5_ASAP7_75T_R%B 2 7 10 15 18 21 29 31 32 37 VSS
c34 37 VSS 0.00657098f $X=0.135 $Y=0.136
c35 32 VSS 1.63059e-19 $X=0.202 $Y=0.135
c36 31 VSS 1.06681e-21 $X=0.163 $Y=0.135
c37 29 VSS 6.5551e-19 $X=0.243 $Y=0.135
c38 21 VSS 0.00869806f $X=0.351 $Y=0.135
c39 18 VSS 0.0683897f $X=0.351 $Y=0.0675
c40 10 VSS 0.0645037f $X=0.297 $Y=0.0675
c41 2 VSS 0.0621762f $X=0.243 $Y=0.0675
r42 31 32 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.163
+ $Y=0.135 $X2=0.202 $Y2=0.135
r43 29 32 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.202 $Y2=0.135
r44 27 37 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.135 $Y2=0.135
r45 27 31 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.163 $Y2=0.135
r46 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r47 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r48 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r49 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r50 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r51 5 29 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r52 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r53 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_NAND2X1P5_ASAP7_75T_R%5 1 2 6 7 11 12 15 17 18 23 24 25 26 33 35 36
+ 37 38 VSS
c29 38 VSS 5.12412e-19 $X=0.2925 $Y=0.072
c30 37 VSS 2.79488e-19 $X=0.261 $Y=0.072
c31 36 VSS 9.73694e-19 $X=0.257 $Y=0.072
c32 35 VSS 4.97766e-19 $X=0.225 $Y=0.072
c33 33 VSS 2.92324e-19 $X=0.324 $Y=0.072
c34 26 VSS 0.0074475f $X=0.202 $Y=0.036
c35 25 VSS 0.00286574f $X=0.144 $Y=0.036
c36 24 VSS 0.00603836f $X=0.216 $Y=0.036
c37 23 VSS 0.0022696f $X=0.216 $Y=0.036
c38 18 VSS 0.0105454f $X=0.108 $Y=0.036
c39 17 VSS 0.0021938f $X=0.108 $Y=0.036
c40 15 VSS 0.0026225f $X=0.324 $Y=0.0675
c41 11 VSS 5.75221e-19 $X=0.341 $Y=0.0675
c42 6 VSS 7.04766e-19 $X=0.233 $Y=0.0675
c43 1 VSS 6.18024e-19 $X=0.125 $Y=0.0675
r44 37 38 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.072 $X2=0.2925 $Y2=0.072
r45 36 37 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.257
+ $Y=0.072 $X2=0.261 $Y2=0.072
r46 35 36 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.072 $X2=0.257 $Y2=0.072
r47 33 38 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.072 $X2=0.2925 $Y2=0.072
r48 29 35 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.072 $X2=0.225 $Y2=0.072
r49 25 26 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.202 $Y2=0.036
r50 23 26 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.202 $Y2=0.036
r51 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r52 17 25 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.144 $Y2=0.036
r53 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r54 15 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.072 $X2=0.324
+ $Y2=0.072
r55 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r56 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r57 10 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r58 10 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072 $X2=0.216
+ $Y2=0.072
r59 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r60 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r61 5 18 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r62 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r63 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends

.subckt PM_NAND2X1P5_ASAP7_75T_R%Y 1 2 6 11 14 16 17 20 21 24 28 37 41 43 44 48
+ 52 53 54 58 60 61 VSS
c33 64 VSS 7.83596e-19 $X=0.405 $Y=0.207
c34 62 VSS 9.22213e-19 $X=0.405 $Y=0.144
c35 61 VSS 0.00237618f $X=0.405 $Y=0.126
c36 60 VSS 6.86417e-19 $X=0.405 $Y=0.081
c37 59 VSS 8.85605e-19 $X=0.405 $Y=0.063
c38 58 VSS 0.00243102f $X=0.405 $Y=0.145
c39 56 VSS 0.00104959f $X=0.405 $Y=0.225
c40 54 VSS 0.00175149f $X=0.358 $Y=0.036
c41 53 VSS 0.00657771f $X=0.338 $Y=0.036
c42 52 VSS 0.00281049f $X=0.378 $Y=0.036
c43 48 VSS 0.00488081f $X=0.27 $Y=0.036
c44 45 VSS 0.00707768f $X=0.396 $Y=0.036
c45 44 VSS 0.00266146f $X=0.367 $Y=0.234
c46 43 VSS 0.00425376f $X=0.338 $Y=0.234
c47 42 VSS 0.00567501f $X=0.2905 $Y=0.234
c48 41 VSS 0.0089446f $X=0.257 $Y=0.234
c49 37 VSS 0.00429709f $X=0.163 $Y=0.234
c50 36 VSS 0.00163196f $X=0.126 $Y=0.234
c51 28 VSS 0.00187319f $X=0.108 $Y=0.234
c52 26 VSS 0.00634021f $X=0.396 $Y=0.234
c53 24 VSS 0.0067281f $X=0.322 $Y=0.2025
c54 20 VSS 0.00783498f $X=0.216 $Y=0.216
c55 16 VSS 5.3314e-19 $X=0.233 $Y=0.216
c56 14 VSS 0.00671331f $X=0.11 $Y=0.2025
c57 11 VSS 4.6121e-19 $X=0.125 $Y=0.2025
c58 9 VSS 2.69461e-19 $X=0.376 $Y=0.0675
c59 1 VSS 6.56704e-19 $X=0.287 $Y=0.0675
r60 63 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.207
r61 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.126 $X2=0.405 $Y2=0.144
r62 60 61 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.081 $X2=0.405 $Y2=0.126
r63 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.063 $X2=0.405 $Y2=0.081
r64 58 63 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.145 $X2=0.405 $Y2=0.189
r65 58 62 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.145 $X2=0.405 $Y2=0.144
r66 56 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.207
r67 55 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.063
r68 53 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.036 $X2=0.358 $Y2=0.036
r69 51 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.358 $Y2=0.036
r70 51 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r71 47 53 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.338 $Y2=0.036
r72 47 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r73 45 55 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r74 45 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.378 $Y2=0.036
r75 43 44 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.234 $X2=0.367 $Y2=0.234
r76 41 42 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.257
+ $Y=0.234 $X2=0.2905 $Y2=0.234
r77 39 43 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.338 $Y2=0.234
r78 39 42 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.2905 $Y2=0.234
r79 36 37 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.163 $Y2=0.234
r80 34 41 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.257 $Y2=0.234
r81 34 37 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.163 $Y2=0.234
r82 28 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r83 26 56 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r84 26 44 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.367 $Y2=0.234
r85 24 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r86 21 24 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.322 $Y2=0.2025
r87 20 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r88 17 20 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.216 $X2=0.216 $Y2=0.216
r89 16 20 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.216 $X2=0.216 $Y2=0.216
r90 14 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r91 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.11 $Y2=0.2025
r92 9 52 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r93 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.0675 $X2=0.376 $Y2=0.0675
r94 5 48 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r95 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
r96 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends


* END of "./NAND2x1p5_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND2x1p5_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 N_5_M0_d N_A_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_5_M1_d N_A_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_5_M2_d N_A_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_B_M3_g N_5_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_B_M4_g N_5_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 N_Y_M5_d N_B_M5_g N_5_M5_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 VDD N_A_M6_g N_Y_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M7 VDD N_A_M7_g N_Y_M7_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.189
M8 VDD N_B_M8_g N_Y_M8_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.189
M9 VDD N_B_M9_g N_Y_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
*
* 
* .include "NAND2x1p5_ASAP7_75t_R.pex.sp.NAND2X1P5_ASAP7_75T_R.pxi"
* BEGIN of "./NAND2x1p5_ASAP7_75t_R.pex.sp.NAND2X1P5_ASAP7_75T_R.pxi"
* File: NAND2x1p5_ASAP7_75t_R.pex.sp.NAND2X1P5_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:38:20 2017
* 
x_PM_NAND2X1P5_ASAP7_75T_R%A N_A_M0_g N_A_M1_g N_A_M6_g N_A_M2_g N_A_c_4_p
+ N_A_M7_g A VSS PM_NAND2X1P5_ASAP7_75T_R%A
x_PM_NAND2X1P5_ASAP7_75T_R%B N_B_M3_g N_B_M8_g N_B_M4_g N_B_M9_g N_B_M5_g
+ N_B_c_26_n N_B_c_39_p N_B_c_27_n N_B_c_28_n B VSS PM_NAND2X1P5_ASAP7_75T_R%B
x_PM_NAND2X1P5_ASAP7_75T_R%5 N_5_M1_d N_5_M0_d N_5_M3_s N_5_M2_d N_5_M5_s
+ N_5_M4_s N_5_c_64_n N_5_c_58_n N_5_c_59_n N_5_c_83_p N_5_c_74_p N_5_c_60_n
+ N_5_c_61_n N_5_c_68_n N_5_c_69_n N_5_c_71_n N_5_c_78_p N_5_c_79_p VSS
+ PM_NAND2X1P5_ASAP7_75T_R%5
x_PM_NAND2X1P5_ASAP7_75T_R%Y N_Y_M4_d N_Y_M3_d N_Y_M5_d N_Y_M6_s N_Y_c_86_n
+ N_Y_M8_s N_Y_M7_s N_Y_c_107_n N_Y_M9_s N_Y_c_94_n N_Y_c_88_n N_Y_c_90_n
+ N_Y_c_91_n N_Y_c_99_n N_Y_c_100_n N_Y_c_101_n N_Y_c_113_n N_Y_c_102_n
+ N_Y_c_103_n Y N_Y_c_118_n N_Y_c_105_n VSS PM_NAND2X1P5_ASAP7_75T_R%Y
cc_1 N_A_M1_g N_B_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_2 N_A_M2_g N_B_M3_g 0.00344695f $X=0.189 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_3 N_A_M2_g N_B_M4_g 2.66145e-19 $X=0.189 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_4 N_A_c_4_p N_B_c_26_n 0.0020914f $X=0.189 $Y=0.1345 $X2=0.351 $Y2=0.135
cc_5 N_A_c_4_p N_B_c_27_n 0.00109734f $X=0.189 $Y=0.1345 $X2=0.163 $Y2=0.135
cc_6 N_A_M2_g N_B_c_28_n 7.24562e-19 $X=0.189 $Y=0.0675 $X2=0.202 $Y2=0.135
cc_7 N_A_c_4_p N_B_c_28_n 0.00297492f $X=0.189 $Y=0.1345 $X2=0.202 $Y2=0.135
cc_8 N_A_M1_g B 6.18619e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.136
cc_9 N_A_c_4_p B 0.00239456f $X=0.189 $Y=0.1345 $X2=0.135 $Y2=0.136
cc_10 A B 0.00188432f $X=0.07 $Y=0.136 $X2=0.135 $Y2=0.136
cc_11 N_A_c_4_p N_5_M1_d 3.8991e-19 $X=0.189 $Y=0.1345 $X2=0.243 $Y2=0.0675
cc_12 A N_5_c_58_n 5.26979e-19 $X=0.07 $Y=0.136 $X2=0.351 $Y2=0.0675
cc_13 N_A_c_4_p N_5_c_59_n 8.45347e-19 $X=0.189 $Y=0.1345 $X2=0.351 $Y2=0.0675
cc_14 N_A_M1_g N_5_c_60_n 2.34767e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 N_A_M2_g N_5_c_61_n 4.27122e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_16 N_A_c_4_p N_5_c_61_n 2.13568e-19 $X=0.189 $Y=0.1345 $X2=0 $Y2=0
cc_17 N_A_c_4_p N_Y_c_86_n 8.01479e-19 $X=0.189 $Y=0.1345 $X2=0.297 $Y2=0.2025
cc_18 A N_Y_c_86_n 0.0013808f $X=0.07 $Y=0.136 $X2=0.297 $Y2=0.2025
cc_19 N_A_c_4_p N_Y_c_88_n 3.08716e-19 $X=0.189 $Y=0.1345 $X2=0.243 $Y2=0.135
cc_20 A N_Y_c_88_n 8.43259e-19 $X=0.07 $Y=0.136 $X2=0.243 $Y2=0.135
cc_21 N_A_M1_g N_Y_c_90_n 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.136
cc_22 N_A_M2_g N_Y_c_91_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_23 N_B_c_26_n N_5_M5_s 3.80371e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.1345
cc_24 N_B_c_26_n N_5_c_64_n 8.0006e-19 $X=0.351 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_25 B N_5_c_59_n 0.00216211f $X=0.135 $Y=0.136 $X2=0.189 $Y2=0.1345
cc_26 B N_5_c_60_n 0.00372796f $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_27 N_B_c_27_n N_5_c_61_n 8.54443e-19 $X=0.163 $Y=0.135 $X2=0 $Y2=0
cc_28 N_B_M4_g N_5_c_68_n 2.83374e-19 $X=0.297 $Y=0.0675 $X2=0.07 $Y2=0.135
cc_29 N_B_c_39_p N_5_c_69_n 0.00189395f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_30 B N_5_c_69_n 3.68725e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_31 N_B_M3_g N_5_c_71_n 4.27107e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_32 N_B_c_26_n N_5_c_71_n 0.00133835f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_33 N_B_c_26_n N_Y_M4_d 3.80413e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_34 B N_Y_c_86_n 0.00157124f $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_35 N_B_c_26_n N_Y_c_94_n 8.0006e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_36 B N_Y_c_90_n 0.00377179f $X=0.135 $Y=0.136 $X2=0.07 $Y2=0.136
cc_37 N_B_M3_g N_Y_c_91_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_38 N_B_c_26_n N_Y_c_91_n 0.00129524f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_39 N_B_c_28_n N_Y_c_91_n 0.00157481f $X=0.202 $Y=0.135 $X2=0 $Y2=0
cc_40 N_B_M4_g N_Y_c_99_n 3.58606e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_41 N_B_M5_g N_Y_c_100_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.07 $Y2=0.1345
cc_42 N_B_c_26_n N_Y_c_101_n 8.0006e-19 $X=0.351 $Y=0.135 $X2=0.189 $Y2=0.1345
cc_43 N_B_M4_g N_Y_c_102_n 2.64781e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_B_M5_g N_Y_c_103_n 3.90391e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_45 N_B_c_26_n N_Y_c_103_n 2.53248e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_46 N_B_c_26_n N_Y_c_105_n 3.35167e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_47 N_5_c_59_n N_Y_c_86_n 0.00122007f $X=0.108 $Y=0.036 $X2=0 $Y2=0
cc_48 N_5_c_74_p N_Y_c_107_n 0.00103326f $X=0.216 $Y=0.036 $X2=0.189 $Y2=0.216
cc_49 N_5_c_64_n N_Y_c_94_n 0.00137166f $X=0.324 $Y=0.0675 $X2=0 $Y2=0
cc_50 N_5_c_64_n N_Y_c_101_n 0.00350506f $X=0.324 $Y=0.0675 $X2=0.189 $Y2=0.1345
cc_51 N_5_c_74_p N_Y_c_101_n 0.00328977f $X=0.216 $Y=0.036 $X2=0.189 $Y2=0.1345
cc_52 N_5_c_78_p N_Y_c_101_n 5.59832e-19 $X=0.261 $Y=0.072 $X2=0.189 $Y2=0.1345
cc_53 N_5_c_79_p N_Y_c_101_n 0.00175493f $X=0.2925 $Y=0.072 $X2=0.189 $Y2=0.1345
cc_54 N_5_c_64_n N_Y_c_113_n 0.00374846f $X=0.324 $Y=0.0675 $X2=0 $Y2=0
cc_55 N_5_c_68_n N_Y_c_113_n 3.97701e-19 $X=0.324 $Y=0.072 $X2=0 $Y2=0
cc_56 N_5_c_64_n N_Y_c_102_n 0.0025091f $X=0.324 $Y=0.0675 $X2=0 $Y2=0
cc_57 N_5_c_83_p N_Y_c_102_n 6.95286e-19 $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_58 N_5_c_79_p N_Y_c_102_n 0.00640856f $X=0.2925 $Y=0.072 $X2=0 $Y2=0
cc_59 N_5_c_68_n N_Y_c_118_n 3.4706e-19 $X=0.324 $Y=0.072 $X2=0 $Y2=0

* END of "./NAND2x1p5_ASAP7_75t_R.pex.sp.NAND2X1P5_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND2x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:38:43 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND2x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND2x2_ASAP7_75t_R.pex.sp.pex"
* File: NAND2x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:38:43 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND2X2_ASAP7_75T_R%B 2 8 11 13 16 21 24 27 32 35 36 37 38 39 42 43
+ 44 45 46 47 50 51 52 53 54 VSS
c75 54 VSS 5.56748e-19 $X=0.459 $Y=0.117
c76 53 VSS 2.64552e-19 $X=0.434 $Y=0.108
c77 52 VSS 0.00120695f $X=0.418 $Y=0.108
c78 51 VSS 0.00127853f $X=0.34 $Y=0.108
c79 50 VSS 2.97889e-19 $X=0.45 $Y=0.108
c80 49 VSS 6.6029e-19 $X=0.331 $Y=0.099
c81 47 VSS 3.12831e-19 $X=0.3005 $Y=0.072
c82 46 VSS 8.46035e-21 $X=0.279 $Y=0.072
c83 45 VSS 3.14008e-19 $X=0.261 $Y=0.072
c84 44 VSS 0.00152288f $X=0.242 $Y=0.072
c85 43 VSS 7.41509e-19 $X=0.218 $Y=0.072
c86 42 VSS 0.0022087f $X=0.322 $Y=0.072
c87 41 VSS 6.6029e-19 $X=0.209 $Y=0.099
c88 39 VSS 2.13186e-19 $X=0.122 $Y=0.108
c89 38 VSS 9.36999e-20 $X=0.109 $Y=0.108
c90 37 VSS 6.87104e-20 $X=0.09 $Y=0.108
c91 36 VSS 0.00248547f $X=0.2 $Y=0.108
c92 35 VSS 6.60211e-19 $X=0.084 $Y=0.152
c93 32 VSS 6.01798e-19 $X=0.081 $Y=0.135
c94 27 VSS 0.00390182f $X=0.459 $Y=0.135
c95 24 VSS 0.0679058f $X=0.459 $Y=0.0675
c96 16 VSS 0.0623886f $X=0.405 $Y=0.0675
c97 11 VSS 0.00381026f $X=0.135 $Y=0.135
c98 8 VSS 0.0623954f $X=0.135 $Y=0.0675
c99 2 VSS 0.0680685f $X=0.081 $Y=0.0675
r100 54 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.117 $X2=0.459 $Y2=0.135
r101 52 53 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.108 $X2=0.434 $Y2=0.108
r102 51 52 5.2963 $w=1.8e-08 $l=7.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.34
+ $Y=0.108 $X2=0.418 $Y2=0.108
r103 50 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.108 $X2=0.459 $Y2=0.117
r104 50 53 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.108 $X2=0.434 $Y2=0.108
r105 49 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.331 $Y=0.099 $X2=0.34 $Y2=0.108
r106 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.331
+ $Y=0.081 $X2=0.331 $Y2=0.099
r107 46 47 1.45988 $w=1.8e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.072 $X2=0.3005 $Y2=0.072
r108 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.072 $X2=0.279 $Y2=0.072
r109 44 45 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.242
+ $Y=0.072 $X2=0.261 $Y2=0.072
r110 43 44 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.218
+ $Y=0.072 $X2=0.242 $Y2=0.072
r111 42 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.322 $Y=0.072 $X2=0.331 $Y2=0.081
r112 42 47 1.45988 $w=1.8e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.322
+ $Y=0.072 $X2=0.3005 $Y2=0.072
r113 40 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.209 $Y=0.081 $X2=0.218 $Y2=0.072
r114 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.209
+ $Y=0.081 $X2=0.209 $Y2=0.099
r115 38 39 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.108 $X2=0.122 $Y2=0.108
r116 37 38 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.108 $X2=0.109 $Y2=0.108
r117 36 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2 $Y=0.108 $X2=0.209 $Y2=0.099
r118 36 39 5.2963 $w=1.8e-08 $l=7.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2
+ $Y=0.108 $X2=0.122 $Y2=0.108
r119 32 35 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.152
r120 29 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.117 $X2=0.09 $Y2=0.108
r121 29 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.117 $X2=0.081 $Y2=0.135
r122 27 56 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r123 24 27 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r124 19 27 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r125 19 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r126 16 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r127 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r128 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r129 5 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r130 5 32 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r131 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NAND2X2_ASAP7_75T_R%A 2 7 10 16 22 25 27 36 VSS
c39 36 VSS 0.00226203f $X=0.272 $Y=0.136
c40 25 VSS 0.0123218f $X=0.351 $Y=0.1345
c41 22 VSS 0.062303f $X=0.351 $Y=0.0675
c42 16 VSS 0.0643897f $X=0.297 $Y=0.0675
c43 10 VSS 0.0645813f $X=0.243 $Y=0.0675
c44 2 VSS 0.0622987f $X=0.189 $Y=0.0675
r45 32 36 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.27 $Y=0.135 $X2=0.27
+ $Y2=0.135
r46 25 27 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.1345 $X2=0.351 $Y2=0.2025
r47 22 25 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.1345
r48 19 25 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.1345 $X2=0.351 $Y2=0.1345
r49 19 32 23.4783 $w=2.3e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.1345 $X2=0.27 $Y2=0.1345
r50 16 19 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.1345
r51 13 32 23.4783 $w=2.3e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.1345 $X2=0.27 $Y2=0.1345
r52 10 13 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.1345
r53 5 13 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.1345 $X2=0.243 $Y2=0.1345
r54 5 7 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1345 $X2=0.189 $Y2=0.2025
r55 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.1345
.ends

.subckt PM_NAND2X2_ASAP7_75T_R%5 1 6 7 11 12 16 17 21 24 28 32 33 34 37 38 39 42
+ 43 44 46 47 48 49 VSS
c41 49 VSS 0.00261806f $X=0.452 $Y=0.036
c42 48 VSS 0.00456882f $X=0.418 $Y=0.036
c43 47 VSS 0.00228092f $X=0.486 $Y=0.036
c44 46 VSS 0.00500247f $X=0.486 $Y=0.036
c45 44 VSS 0.0015425f $X=0.359 $Y=0.036
c46 43 VSS 0.0107131f $X=0.34 $Y=0.036
c47 42 VSS 0.00713099f $X=0.378 $Y=0.036
c48 39 VSS 0.00520575f $X=0.235 $Y=0.036
c49 38 VSS 0.0044884f $X=0.2 $Y=0.036
c50 37 VSS 0.0100322f $X=0.27 $Y=0.036
c51 34 VSS 0.00162279f $X=0.142 $Y=0.036
c52 33 VSS 0.00762831f $X=0.122 $Y=0.036
c53 32 VSS 0.00713099f $X=0.162 $Y=0.036
c54 28 VSS 0.00228092f $X=0.054 $Y=0.036
c55 24 VSS 3.4551e-19 $X=0.484 $Y=0.0675
c56 16 VSS 7.6997e-19 $X=0.395 $Y=0.0675
c57 11 VSS 6.26354e-19 $X=0.287 $Y=0.0675
c58 6 VSS 7.6997e-19 $X=0.179 $Y=0.0675
c59 1 VSS 3.4551e-19 $X=0.071 $Y=0.0675
r60 48 49 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.036 $X2=0.452 $Y2=0.036
r61 46 49 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.452 $Y2=0.036
r62 46 47 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036 $X2=0.486
+ $Y2=0.036
r63 43 44 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.34
+ $Y=0.036 $X2=0.359 $Y2=0.036
r64 41 48 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.418 $Y2=0.036
r65 41 44 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.359 $Y2=0.036
r66 41 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r67 38 39 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2
+ $Y=0.036 $X2=0.235 $Y2=0.036
r68 36 43 4.75309 $w=1.8e-08 $l=7e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.34 $Y2=0.036
r69 36 39 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.235 $Y2=0.036
r70 36 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r71 33 34 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.122
+ $Y=0.036 $X2=0.142 $Y2=0.036
r72 31 38 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.2 $Y2=0.036
r73 31 34 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.142 $Y2=0.036
r74 31 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r75 27 33 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.122 $Y2=0.036
r76 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r77 24 47 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0675 $X2=0.486 $Y2=0.036
r78 21 24 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.484 $Y2=0.0675
r79 20 42 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r80 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.378 $Y2=0.0675
r81 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.0675 $X2=0.378 $Y2=0.0675
r82 15 37 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r83 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r84 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r85 10 32 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r86 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r87 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r88 4 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r89 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends

.subckt PM_NAND2X2_ASAP7_75T_R%Y 1 2 5 6 7 10 11 14 16 19 21 24 26 29 34 37 40
+ 48 52 53 57 58 59 60 64 65 71 72 76 78 VSS
c65 80 VSS 0.00130599f $X=0.513 $Y=0.207
c66 78 VSS 9.39445e-19 $X=0.513 $Y=0.122
c67 77 VSS 7.39581e-19 $X=0.513 $Y=0.099
c68 76 VSS 0.0023804f $X=0.514 $Y=0.145
c69 74 VSS 9.03568e-19 $X=0.513 $Y=0.225
c70 72 VSS 4.78169e-19 $X=0.5 $Y=0.072
c71 71 VSS 8.46035e-21 $X=0.468 $Y=0.072
c72 66 VSS 0.00220485f $X=0.504 $Y=0.072
c73 65 VSS 0.00146362f $X=0.468 $Y=0.234
c74 64 VSS 0.0137555f $X=0.45 $Y=0.234
c75 60 VSS 0.00395819f $X=0.322 $Y=0.234
c76 59 VSS 0.00324847f $X=0.279 $Y=0.234
c77 58 VSS 0.00226617f $X=0.242 $Y=0.234
c78 57 VSS 0.00608839f $X=0.218 $Y=0.234
c79 53 VSS 0.00606865f $X=0.1625 $Y=0.234
c80 52 VSS 0.00142953f $X=0.109 $Y=0.234
c81 48 VSS 0.00146362f $X=0.09 $Y=0.234
c82 47 VSS 0.00346625f $X=0.072 $Y=0.234
c83 43 VSS 0.00350046f $X=0.036 $Y=0.234
c84 42 VSS 0.00696671f $X=0.504 $Y=0.234
c85 40 VSS 4.78169e-19 $X=0.072 $Y=0.072
c86 39 VSS 2.76758e-19 $X=0.04 $Y=0.072
c87 37 VSS 8.46035e-21 $X=0.108 $Y=0.072
c88 35 VSS 0.00192809f $X=0.036 $Y=0.072
c89 34 VSS 0.00462133f $X=0.027 $Y=0.207
c90 33 VSS 7.39581e-19 $X=0.027 $Y=0.099
c91 32 VSS 9.03568e-19 $X=0.027 $Y=0.225
c92 29 VSS 0.0069163f $X=0.43 $Y=0.2025
c93 24 VSS 0.0071986f $X=0.326 $Y=0.2025
c94 21 VSS 4.6121e-19 $X=0.341 $Y=0.2025
c95 19 VSS 0.00765911f $X=0.214 $Y=0.2025
c96 14 VSS 0.0069473f $X=0.11 $Y=0.2025
c97 11 VSS 4.59792e-19 $X=0.125 $Y=0.2025
c98 10 VSS 0.00283195f $X=0.432 $Y=0.0675
c99 6 VSS 6.19444e-19 $X=0.449 $Y=0.0675
c100 5 VSS 0.00283195f $X=0.108 $Y=0.0675
c101 1 VSS 6.18143e-19 $X=0.125 $Y=0.0675
r102 79 80 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.177 $X2=0.513 $Y2=0.207
r103 77 78 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.099 $X2=0.513 $Y2=0.122
r104 76 79 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.145 $X2=0.513 $Y2=0.177
r105 76 78 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.145 $X2=0.513 $Y2=0.122
r106 74 80 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.207
r107 73 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.081 $X2=0.513 $Y2=0.099
r108 71 72 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.072 $X2=0.5 $Y2=0.072
r109 68 71 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.072 $X2=0.468 $Y2=0.072
r110 66 73 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.072 $X2=0.513 $Y2=0.081
r111 66 72 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.072 $X2=0.5 $Y2=0.072
r112 64 65 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r113 62 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.45 $Y2=0.234
r114 59 60 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.234 $X2=0.322 $Y2=0.234
r115 58 59 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.242
+ $Y=0.234 $X2=0.279 $Y2=0.234
r116 57 58 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.218
+ $Y=0.234 $X2=0.242 $Y2=0.234
r117 55 62 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r118 55 60 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.322 $Y2=0.234
r119 52 53 3.63272 $w=1.8e-08 $l=5.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.234 $X2=0.1625 $Y2=0.234
r120 50 57 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.218 $Y2=0.234
r121 50 53 3.63272 $w=1.8e-08 $l=5.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.1625 $Y2=0.234
r122 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r123 45 52 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.109 $Y2=0.234
r124 45 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.09 $Y2=0.234
r125 43 47 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.072 $Y2=0.234
r126 42 74 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.234 $X2=0.513 $Y2=0.225
r127 42 65 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.468 $Y2=0.234
r128 39 40 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.072 $X2=0.072 $Y2=0.072
r129 37 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.072 $Y2=0.072
r130 35 39 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.072 $X2=0.04 $Y2=0.072
r131 33 34 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.099 $X2=0.027 $Y2=0.207
r132 32 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.225 $X2=0.036 $Y2=0.234
r133 32 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.207
r134 31 35 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.081 $X2=0.036 $Y2=0.072
r135 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.081 $X2=0.027 $Y2=0.099
r136 29 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r137 26 29 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.43 $Y2=0.2025
r138 24 55 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r139 21 24 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.326 $Y2=0.2025
r140 19 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r141 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.214 $Y2=0.2025
r142 14 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r143 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.11 $Y2=0.2025
r144 10 68 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.072
+ $X2=0.432 $Y2=0.072
r145 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r146 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r147 5 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072 $X2=0.108
+ $Y2=0.072
r148 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r149 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends


* END of "./NAND2x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND2x2_ASAP7_75t_R  VSS VDD B A Y
* 
* Y	Y
* A	A
* B	B
M0 N_Y_M0_d N_B_M0_g N_5_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_Y_M1_d N_B_M1_g N_5_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_A_M2_g N_5_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 VSS N_A_M3_g N_5_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 VSS N_A_M4_g N_5_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 VSS N_A_M5_g N_5_M5_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_B_M6_g N_5_M6_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_Y_M7_d N_B_M7_g N_5_M7_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 VDD N_B_M8_g N_Y_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M9 N_Y_M9_d N_A_M9_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M10 N_Y_M10_d N_A_M10_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M11 VDD N_B_M11_g N_Y_M11_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
*
* 
* .include "NAND2x2_ASAP7_75t_R.pex.sp.NAND2X2_ASAP7_75T_R.pxi"
* BEGIN of "./NAND2x2_ASAP7_75t_R.pex.sp.NAND2X2_ASAP7_75T_R.pxi"
* File: NAND2x2_ASAP7_75t_R.pex.sp.NAND2X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:38:43 2017
* 
x_PM_NAND2X2_ASAP7_75T_R%B N_B_M0_g N_B_M1_g N_B_c_11_p N_B_M8_g N_B_M6_g
+ N_B_M11_g N_B_M7_g N_B_c_12_p N_B_c_17_p B N_B_c_3_p N_B_c_22_p N_B_c_41_p
+ N_B_c_42_p N_B_c_32_p N_B_c_24_p N_B_c_14_p N_B_c_5_p N_B_c_19_p N_B_c_7_p
+ N_B_c_37_p N_B_c_16_p N_B_c_10_p N_B_c_46_p N_B_c_21_p VSS
+ PM_NAND2X2_ASAP7_75T_R%B
x_PM_NAND2X2_ASAP7_75T_R%A N_A_M2_g N_A_M9_g N_A_M3_g N_A_M4_g N_A_M5_g
+ N_A_c_86_n N_A_M10_g A VSS PM_NAND2X2_ASAP7_75T_R%A
x_PM_NAND2X2_ASAP7_75T_R%5 N_5_M0_s N_5_M2_s N_5_M1_s N_5_M4_s N_5_M3_s N_5_M6_s
+ N_5_M5_s N_5_M7_s N_5_c_152_p N_5_c_115_n N_5_c_116_n N_5_c_118_n N_5_c_119_n
+ N_5_c_121_n N_5_c_135_n N_5_c_124_n N_5_c_125_n N_5_c_127_n N_5_c_128_n
+ N_5_c_129_n N_5_c_130_n N_5_c_131_n N_5_c_144_p VSS PM_NAND2X2_ASAP7_75T_R%5
x_PM_NAND2X2_ASAP7_75T_R%Y N_Y_M1_d N_Y_M0_d N_Y_c_157_n N_Y_M7_d N_Y_M6_d
+ N_Y_c_161_n N_Y_M8_s N_Y_c_165_n N_Y_M9_d N_Y_c_193_n N_Y_M10_d N_Y_c_195_n
+ N_Y_M11_s N_Y_c_168_n N_Y_c_170_n N_Y_c_172_n N_Y_c_212_n N_Y_c_175_n
+ N_Y_c_177_n N_Y_c_178_n N_Y_c_181_n N_Y_c_199_n N_Y_c_200_n N_Y_c_201_n
+ N_Y_c_182_n N_Y_c_185_n N_Y_c_187_n N_Y_c_217_n Y N_Y_c_192_n VSS
+ PM_NAND2X2_ASAP7_75T_R%Y
cc_1 N_B_M0_g N_A_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_B_M1_g N_A_M2_g 0.0032073f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_B_c_3_p N_A_M2_g 4.19577e-19 $X=0.2 $Y=0.108 $X2=0.189 $Y2=0.0675
cc_4 N_B_M1_g N_A_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_5 N_B_c_5_p N_A_M3_g 2.1804e-19 $X=0.261 $Y=0.072 $X2=0.243 $Y2=0.0675
cc_6 N_B_M6_g N_A_M4_g 2.31381e-19 $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_7 N_B_c_7_p N_A_M4_g 2.66132e-19 $X=0.3005 $Y=0.072 $X2=0.297 $Y2=0.0675
cc_8 N_B_M6_g N_A_M5_g 0.0032073f $X=0.405 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_9 N_B_M7_g N_A_M5_g 2.66145e-19 $X=0.459 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_10 N_B_c_10_p N_A_M5_g 4.19577e-19 $X=0.418 $Y=0.108 $X2=0.351 $Y2=0.0675
cc_11 N_B_c_11_p N_A_c_86_n 0.00227362f $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.1345
cc_12 N_B_c_12_p N_A_c_86_n 0.00227362f $X=0.459 $Y=0.135 $X2=0.351 $Y2=0.1345
cc_13 N_B_c_3_p N_A_c_86_n 0.00124067f $X=0.2 $Y=0.108 $X2=0.351 $Y2=0.1345
cc_14 N_B_c_14_p N_A_c_86_n 8.12001e-19 $X=0.242 $Y=0.072 $X2=0.351 $Y2=0.1345
cc_15 N_B_c_7_p N_A_c_86_n 8.41977e-19 $X=0.3005 $Y=0.072 $X2=0.351 $Y2=0.1345
cc_16 N_B_c_16_p N_A_c_86_n 0.00124067f $X=0.34 $Y=0.108 $X2=0.351 $Y2=0.1345
cc_17 N_B_c_17_p A 5.14434e-19 $X=0.081 $Y=0.135 $X2=0.272 $Y2=0.136
cc_18 N_B_c_3_p A 4.72303e-19 $X=0.2 $Y=0.108 $X2=0.272 $Y2=0.136
cc_19 N_B_c_19_p A 0.00101457f $X=0.279 $Y=0.072 $X2=0.272 $Y2=0.136
cc_20 N_B_c_16_p A 6.2809e-19 $X=0.34 $Y=0.108 $X2=0.272 $Y2=0.136
cc_21 N_B_c_21_p A 4.36649e-19 $X=0.459 $Y=0.117 $X2=0.272 $Y2=0.136
cc_22 N_B_c_22_p N_5_c_115_n 2.78572e-19 $X=0.09 $Y=0.108 $X2=0 $Y2=0
cc_23 N_B_c_3_p N_5_c_116_n 0.00201076f $X=0.2 $Y=0.108 $X2=0.27 $Y2=0.135
cc_24 N_B_c_24_p N_5_c_116_n 7.67394e-19 $X=0.218 $Y=0.072 $X2=0.27 $Y2=0.135
cc_25 N_B_M0_g N_5_c_118_n 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_B_M1_g N_5_c_119_n 3.24635e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_B_c_3_p N_5_c_119_n 0.00230303f $X=0.2 $Y=0.108 $X2=0 $Y2=0
cc_28 N_B_c_5_p N_5_c_121_n 5.61323e-19 $X=0.261 $Y=0.072 $X2=0 $Y2=0
cc_29 N_B_c_19_p N_5_c_121_n 0.00124096f $X=0.279 $Y=0.072 $X2=0 $Y2=0
cc_30 N_B_c_7_p N_5_c_121_n 5.58359e-19 $X=0.3005 $Y=0.072 $X2=0 $Y2=0
cc_31 N_B_c_24_p N_5_c_124_n 0.0059448f $X=0.218 $Y=0.072 $X2=0 $Y2=0
cc_32 N_B_c_32_p N_5_c_125_n 7.67394e-19 $X=0.322 $Y=0.072 $X2=0 $Y2=0
cc_33 N_B_c_10_p N_5_c_125_n 0.00201076f $X=0.418 $Y=0.108 $X2=0 $Y2=0
cc_34 N_B_c_19_p N_5_c_127_n 0.0059448f $X=0.279 $Y=0.072 $X2=0.243 $Y2=0.1345
cc_35 N_B_c_10_p N_5_c_128_n 0.00230302f $X=0.418 $Y=0.108 $X2=0.27 $Y2=0.1345
cc_36 N_B_M7_g N_5_c_129_n 2.08515e-19 $X=0.459 $Y=0.0675 $X2=0.351 $Y2=0.1345
cc_37 N_B_c_37_p N_5_c_130_n 2.78572e-19 $X=0.45 $Y=0.108 $X2=0 $Y2=0
cc_38 N_B_M6_g N_5_c_131_n 3.81924e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_B_c_11_p N_Y_M1_d 3.70143e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_40 N_B_c_11_p N_Y_c_157_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.1345
cc_41 N_B_c_41_p N_Y_c_157_n 7.62637e-19 $X=0.109 $Y=0.108 $X2=0.189 $Y2=0.1345
cc_42 N_B_c_42_p N_Y_c_157_n 8.29904e-19 $X=0.122 $Y=0.108 $X2=0.189 $Y2=0.1345
cc_43 N_B_c_12_p N_Y_M7_d 3.70143e-19 $X=0.459 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_44 N_B_c_12_p N_Y_c_161_n 8.0006e-19 $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_45 N_B_c_37_p N_Y_c_161_n 6.01614e-19 $X=0.45 $Y=0.108 $X2=0.243 $Y2=0.0675
cc_46 N_B_c_46_p N_Y_c_161_n 9.90927e-19 $X=0.434 $Y=0.108 $X2=0.243 $Y2=0.0675
cc_47 B N_Y_M8_s 2.0764e-19 $X=0.084 $Y=0.152 $X2=0 $Y2=0
cc_48 N_B_c_11_p N_Y_c_165_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_49 N_B_c_17_p N_Y_c_165_n 9.47875e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_50 B N_Y_c_165_n 0.00166646f $X=0.084 $Y=0.152 $X2=0 $Y2=0
cc_51 N_B_c_12_p N_Y_c_168_n 8.0006e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_52 N_B_c_21_p N_Y_c_168_n 5.27536e-19 $X=0.459 $Y=0.117 $X2=0 $Y2=0
cc_53 N_B_c_11_p N_Y_c_170_n 3.39417e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_54 N_B_c_22_p N_Y_c_170_n 0.00519692f $X=0.09 $Y=0.108 $X2=0 $Y2=0
cc_55 N_B_M0_g N_Y_c_172_n 2.52885e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_56 N_B_c_22_p N_Y_c_172_n 0.00408818f $X=0.09 $Y=0.108 $X2=0 $Y2=0
cc_57 N_B_c_24_p N_Y_c_172_n 2.95701e-19 $X=0.218 $Y=0.072 $X2=0 $Y2=0
cc_58 N_B_M0_g N_Y_c_175_n 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_59 B N_Y_c_175_n 0.00371886f $X=0.084 $Y=0.152 $X2=0 $Y2=0
cc_60 N_B_c_41_p N_Y_c_177_n 4.64167e-19 $X=0.109 $Y=0.108 $X2=0 $Y2=0
cc_61 N_B_M1_g N_Y_c_178_n 4.52603e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_62 N_B_c_11_p N_Y_c_178_n 3.30932e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_63 N_B_c_42_p N_Y_c_178_n 4.64167e-19 $X=0.122 $Y=0.108 $X2=0 $Y2=0
cc_64 N_B_c_3_p N_Y_c_181_n 4.64167e-19 $X=0.2 $Y=0.108 $X2=0 $Y2=0
cc_65 N_B_M6_g N_Y_c_182_n 4.52603e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_66 N_B_c_12_p N_Y_c_182_n 4.74833e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_67 N_B_c_16_p N_Y_c_182_n 0.00160573f $X=0.34 $Y=0.108 $X2=0 $Y2=0
cc_68 N_B_M7_g N_Y_c_185_n 3.30638e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_69 N_B_c_21_p N_Y_c_185_n 6.86694e-19 $X=0.459 $Y=0.117 $X2=0 $Y2=0
cc_70 N_B_M7_g N_Y_c_187_n 2.52885e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_71 N_B_c_32_p N_Y_c_187_n 2.95701e-19 $X=0.322 $Y=0.072 $X2=0 $Y2=0
cc_72 N_B_c_46_p N_Y_c_187_n 0.00407975f $X=0.434 $Y=0.108 $X2=0 $Y2=0
cc_73 N_B_c_12_p Y 3.39417e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_74 N_B_c_21_p Y 0.00186387f $X=0.459 $Y=0.117 $X2=0 $Y2=0
cc_75 N_B_c_37_p N_Y_c_192_n 0.00186387f $X=0.45 $Y=0.108 $X2=0 $Y2=0
cc_76 N_A_c_86_n N_5_M4_s 3.89915e-19 $X=0.351 $Y=0.1345 $X2=0.135 $Y2=0.135
cc_77 N_A_c_86_n N_5_c_121_n 0.00227427f $X=0.351 $Y=0.1345 $X2=0.09 $Y2=0.108
cc_78 A N_5_c_121_n 0.0438982f $X=0.272 $Y=0.136 $X2=0.09 $Y2=0.108
cc_79 N_A_M2_g N_5_c_135_n 3.80935e-19 $X=0.189 $Y=0.0675 $X2=0.109 $Y2=0.108
cc_80 N_A_M3_g N_5_c_127_n 2.34767e-19 $X=0.243 $Y=0.0675 $X2=0.218 $Y2=0.072
cc_81 N_A_M4_g N_5_c_127_n 2.64526e-19 $X=0.297 $Y=0.0675 $X2=0.218 $Y2=0.072
cc_82 N_A_M5_g N_5_c_128_n 3.42841e-19 $X=0.351 $Y=0.0675 $X2=0.242 $Y2=0.072
cc_83 N_A_c_86_n N_Y_c_193_n 8.01479e-19 $X=0.351 $Y=0.1345 $X2=0.405 $Y2=0.135
cc_84 A N_Y_c_193_n 0.00105831f $X=0.272 $Y=0.136 $X2=0.405 $Y2=0.135
cc_85 N_A_c_86_n N_Y_c_195_n 8.01479e-19 $X=0.351 $Y=0.1345 $X2=0.459 $Y2=0.0675
cc_86 A N_Y_c_195_n 0.00105316f $X=0.272 $Y=0.136 $X2=0.459 $Y2=0.0675
cc_87 N_A_M2_g N_Y_c_181_n 4.52603e-19 $X=0.189 $Y=0.0675 $X2=0.459 $Y2=0.135
cc_88 N_A_c_86_n N_Y_c_181_n 5.47817e-19 $X=0.351 $Y=0.1345 $X2=0.459 $Y2=0.135
cc_89 N_A_M3_g N_Y_c_199_n 2.08223e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_90 A N_Y_c_200_n 0.0035884f $X=0.272 $Y=0.136 $X2=0 $Y2=0
cc_91 N_A_M4_g N_Y_c_201_n 4.62717e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_92 N_A_c_86_n N_Y_c_201_n 7.12009e-19 $X=0.351 $Y=0.1345 $X2=0.081 $Y2=0.135
cc_93 N_A_M5_g N_Y_c_182_n 4.52603e-19 $X=0.351 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_94 N_5_c_115_n N_Y_c_157_n 0.00384463f $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.135
cc_95 N_5_c_116_n N_Y_c_157_n 0.00363853f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.135
cc_96 N_5_c_118_n N_Y_c_157_n 0.0025091f $X=0.122 $Y=0.036 $X2=0.081 $Y2=0.135
cc_97 N_5_c_125_n N_Y_c_161_n 0.00363853f $X=0.378 $Y=0.036 $X2=0.135 $Y2=0.135
cc_98 N_5_c_130_n N_Y_c_161_n 0.00384463f $X=0.486 $Y=0.036 $X2=0.135 $Y2=0.135
cc_99 N_5_c_144_p N_Y_c_161_n 0.0025091f $X=0.452 $Y=0.036 $X2=0.135 $Y2=0.135
cc_100 N_5_c_115_n N_Y_c_170_n 2.86097e-19 $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.152
cc_101 N_5_c_116_n N_Y_c_172_n 4.45525e-19 $X=0.162 $Y=0.036 $X2=0.09 $Y2=0.108
cc_102 N_5_M0_s N_Y_c_212_n 2.53396e-19 $X=0.071 $Y=0.0675 $X2=0.209 $Y2=0.081
cc_103 N_5_c_115_n N_Y_c_212_n 0.00263302f $X=0.054 $Y=0.036 $X2=0.209 $Y2=0.081
cc_104 N_5_c_118_n N_Y_c_212_n 0.00709175f $X=0.122 $Y=0.036 $X2=0.209 $Y2=0.081
cc_105 N_5_c_125_n N_Y_c_187_n 4.45525e-19 $X=0.378 $Y=0.036 $X2=0 $Y2=0
cc_106 N_5_c_144_p N_Y_c_187_n 0.00354594f $X=0.452 $Y=0.036 $X2=0 $Y2=0
cc_107 N_5_c_152_p N_Y_c_217_n 2.53396e-19 $X=0.484 $Y=0.0675 $X2=0 $Y2=0
cc_108 N_5_c_129_n N_Y_c_217_n 0.00354594f $X=0.486 $Y=0.036 $X2=0 $Y2=0
cc_109 N_5_c_130_n N_Y_c_217_n 0.00263302f $X=0.486 $Y=0.036 $X2=0 $Y2=0
cc_110 N_5_c_130_n N_Y_c_192_n 2.86097e-19 $X=0.486 $Y=0.036 $X2=0 $Y2=0

* END of "./NAND2x2_ASAP7_75t_R.pex.sp.NAND2X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND2xp33_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:39:05 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND2xp33_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND2xp33_ASAP7_75t_R.pex.sp.pex"
* File: NAND2xp33_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:39:05 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND2XP33_ASAP7_75T_R%A 2 5 7 19 VSS
c5 19 VSS 0.0263471f $X=0.06 $Y=0.135
c6 5 VSS 0.00582264f $X=0.081 $Y=0.135
c7 2 VSS 0.0643819f $X=0.081 $Y=0.054
r8 19 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r9 5 23 18.8889 $w=1.8e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r10 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2295
r11 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NAND2XP33_ASAP7_75T_R%B 2 5 7 12 VSS
c10 12 VSS 0.00423739f $X=0.135 $Y=0.135
c11 5 VSS 0.00156845f $X=0.135 $Y=0.135
c12 2 VSS 0.0638285f $X=0.135 $Y=0.054
r13 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r14 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2295
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_NAND2XP33_ASAP7_75T_R%Y 1 4 6 7 13 18 22 30 32 VSS
c8 34 VSS 4.55454e-19 $X=0.189 $Y=0.216
c9 32 VSS 0.00150666f $X=0.189 $Y=0.099
c10 31 VSS 8.85605e-19 $X=0.189 $Y=0.063
c11 30 VSS 0.00490677f $X=0.19 $Y=0.135
c12 28 VSS 4.30151e-19 $X=0.189 $Y=0.225
c13 22 VSS 0.00166239f $X=0.162 $Y=0.036
c14 20 VSS 0.00607663f $X=0.18 $Y=0.036
c15 19 VSS 0.00303662f $X=0.162 $Y=0.234
c16 18 VSS 0.00288209f $X=0.144 $Y=0.234
c17 13 VSS 0.0023094f $X=0.108 $Y=0.234
c18 11 VSS 0.00621531f $X=0.18 $Y=0.234
c19 10 VSS 0.00562504f $X=0.108 $Y=0.2295
c20 6 VSS 6.15566e-19 $X=0.125 $Y=0.2295
c21 4 VSS 0.0041197f $X=0.16 $Y=0.054
r22 33 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.207 $X2=0.189 $Y2=0.216
r23 31 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.063 $X2=0.189 $Y2=0.099
r24 30 33 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.207
r25 30 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.099
r26 28 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.216
r27 27 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r28 20 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r29 20 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.162 $Y2=0.036
r30 18 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.162 $Y2=0.234
r31 13 18 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.144 $Y2=0.234
r32 11 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.234 $X2=0.189 $Y2=0.225
r33 11 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.162 $Y2=0.234
r34 10 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r35 7 10 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2295 $X2=0.108 $Y2=0.2295
r36 6 10 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2295 $X2=0.108 $Y2=0.2295
r37 4 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r38 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.054 $X2=0.16 $Y2=0.054
.ends

.subckt PM_NAND2XP33_ASAP7_75T_R%6 1 2 VSS
c1 1 VSS 0.00221012f $X=0.125 $Y=0.054
r2 1 2 25.1852 $w=5.4e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.054 $X2=0.091 $Y2=0.054
.ends


* END of "./NAND2xp33_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND2xp33_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 N_6_M0_d N_A_M0_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_B_M1_g N_6_M1_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_A_M2_g VDD VDD PMOS_RVT L=2e-08 W=2.7e-08 NFIN=1 $X=0.071 $Y=0.216
M3 VDD N_B_M3_g N_Y_M3_s VDD PMOS_RVT L=2e-08 W=2.7e-08 NFIN=1 $X=0.125 $Y=0.216
*
* 
* .include "NAND2xp33_ASAP7_75t_R.pex.sp.NAND2XP33_ASAP7_75T_R.pxi"
* BEGIN of "./NAND2xp33_ASAP7_75t_R.pex.sp.NAND2XP33_ASAP7_75T_R.pxi"
* File: NAND2xp33_ASAP7_75t_R.pex.sp.NAND2XP33_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:39:05 2017
* 
x_PM_NAND2XP33_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M2_g A VSS
+ PM_NAND2XP33_ASAP7_75T_R%A
x_PM_NAND2XP33_ASAP7_75T_R%B N_B_M1_g N_B_c_7_n N_B_M3_g B VSS
+ PM_NAND2XP33_ASAP7_75T_R%B
x_PM_NAND2XP33_ASAP7_75T_R%Y N_Y_M1_d N_Y_c_18_n N_Y_M3_s N_Y_M2_d N_Y_c_16_n
+ N_Y_c_19_n N_Y_c_17_n Y N_Y_c_23_n VSS PM_NAND2XP33_ASAP7_75T_R%Y
x_PM_NAND2XP33_ASAP7_75T_R%6 N_6_M1_s N_6_M0_d VSS PM_NAND2XP33_ASAP7_75T_R%6
cc_1 N_A_M0_g N_B_M1_g 0.00344695f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A_c_2_p N_B_c_7_n 8.71247e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A B 0.0027917f $X=0.06 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 A N_Y_c_16_n 5.24213e-19 $X=0.06 $Y=0.135 $X2=0 $Y2=0
cc_5 A N_Y_c_17_n 2.61367e-19 $X=0.06 $Y=0.135 $X2=0 $Y2=0
cc_6 B N_Y_c_18_n 6.42527e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_7 N_B_M1_g N_Y_c_19_n 2.25474e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_8 B N_Y_c_19_n 0.0036051f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_9 N_B_M1_g N_Y_c_17_n 3.14377e-19 $X=0.135 $Y=0.054 $X2=0.064 $Y2=0.135
cc_10 B Y 0.00340582f $X=0.135 $Y=0.135 $X2=0.064 $Y2=0.135
cc_11 B N_Y_c_23_n 0.00340582f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_12 B N_6_M1_s 2.75518e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.054

* END of "./NAND2xp33_ASAP7_75t_R.pex.sp.NAND2XP33_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND2xp5_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:39:28 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND2xp5_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND2xp5_ASAP7_75t_R.pex.sp.pex"
* File: NAND2xp5_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:39:28 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND2XP5_ASAP7_75T_R%A 2 5 7 19 VSS
c6 19 VSS 0.0261022f $X=0.06 $Y=0.135
c7 5 VSS 0.00677211f $X=0.081 $Y=0.135
c8 2 VSS 0.0643819f $X=0.081 $Y=0.0675
r9 19 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r10 5 23 18.8889 $w=1.8e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r11 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r12 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NAND2XP5_ASAP7_75T_R%B 2 5 7 12 17 19 VSS
c12 19 VSS 3.77561e-20 $X=0.135 $Y=0.148
c13 17 VSS 0.00163815f $X=0.135 $Y=0.152
c14 12 VSS 0.00315936f $X=0.135 $Y=0.135
c15 5 VSS 0.00156845f $X=0.135 $Y=0.135
c16 2 VSS 0.0638285f $X=0.135 $Y=0.0675
r17 18 19 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.148
r18 17 19 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.152 $X2=0.135 $Y2=0.148
r19 12 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r20 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r21 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_NAND2XP5_ASAP7_75T_R%Y 1 6 7 10 13 18 22 23 30 32 VSS
c9 34 VSS 4.55454e-19 $X=0.189 $Y=0.216
c10 32 VSS 3.29451e-19 $X=0.189 $Y=0.073
c11 31 VSS 8.85605e-19 $X=0.189 $Y=0.063
c12 30 VSS 0.00599446f $X=0.19 $Y=0.083
c13 28 VSS 4.30151e-19 $X=0.189 $Y=0.225
c14 23 VSS 0.00465482f $X=0.162 $Y=0.036
c15 22 VSS 0.00165544f $X=0.162 $Y=0.036
c16 20 VSS 0.00604756f $X=0.18 $Y=0.036
c17 19 VSS 0.00280896f $X=0.162 $Y=0.234
c18 18 VSS 0.00287092f $X=0.144 $Y=0.234
c19 13 VSS 0.00225637f $X=0.108 $Y=0.234
c20 11 VSS 0.00599224f $X=0.18 $Y=0.234
c21 10 VSS 0.00801905f $X=0.108 $Y=0.216
c22 6 VSS 6.05457e-19 $X=0.125 $Y=0.216
c23 4 VSS 2.69461e-19 $X=0.16 $Y=0.0675
r24 33 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.207 $X2=0.189 $Y2=0.216
r25 31 32 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.063 $X2=0.189 $Y2=0.073
r26 30 33 8.41975 $w=1.8e-08 $l=1.24e-07 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.083 $X2=0.189 $Y2=0.207
r27 30 32 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.083 $X2=0.189 $Y2=0.073
r28 28 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.216
r29 27 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r30 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r31 20 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r32 20 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.162 $Y2=0.036
r33 18 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.162 $Y2=0.234
r34 13 18 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.144 $Y2=0.234
r35 11 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.234 $X2=0.189 $Y2=0.225
r36 11 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.162 $Y2=0.234
r37 10 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r38 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.216 $X2=0.108 $Y2=0.216
r39 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.216 $X2=0.108 $Y2=0.216
r40 4 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r41 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.0675 $X2=0.16 $Y2=0.0675
.ends

.subckt PM_NAND2XP5_ASAP7_75T_R%6 1 2 VSS
c1 1 VSS 0.00224788f $X=0.125 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends


* END of "./NAND2xp5_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND2xp5_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 N_6_M0_d N_A_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_B_M1_g N_6_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_A_M2_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M3 VDD N_B_M3_g N_Y_M3_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
*
* 
* .include "NAND2xp5_ASAP7_75t_R.pex.sp.NAND2XP5_ASAP7_75T_R.pxi"
* BEGIN of "./NAND2xp5_ASAP7_75t_R.pex.sp.NAND2XP5_ASAP7_75T_R.pxi"
* File: NAND2xp5_ASAP7_75t_R.pex.sp.NAND2XP5_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:39:28 2017
* 
x_PM_NAND2XP5_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M2_g A VSS
+ PM_NAND2XP5_ASAP7_75T_R%A
x_PM_NAND2XP5_ASAP7_75T_R%B N_B_M1_g N_B_c_8_n N_B_M3_g N_B_c_9_n B N_B_c_10_n
+ VSS PM_NAND2XP5_ASAP7_75T_R%B
x_PM_NAND2XP5_ASAP7_75T_R%Y N_Y_M1_d N_Y_M3_s N_Y_M2_d N_Y_c_21_n N_Y_c_19_n
+ N_Y_c_22_n N_Y_c_20_n N_Y_c_25_n Y N_Y_c_27_n VSS PM_NAND2XP5_ASAP7_75T_R%Y
x_PM_NAND2XP5_ASAP7_75T_R%6 N_6_M1_s N_6_M0_d VSS PM_NAND2XP5_ASAP7_75T_R%6
cc_1 N_A_M0_g N_B_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_8_n 8.71247e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A N_B_c_9_n 0.00123389f $X=0.06 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 A N_B_c_10_n 8.2966e-19 $X=0.06 $Y=0.135 $X2=0.135 $Y2=0.148
cc_5 A N_Y_c_19_n 5.24213e-19 $X=0.06 $Y=0.135 $X2=0.135 $Y2=0.135
cc_6 A N_Y_c_20_n 2.61367e-19 $X=0.06 $Y=0.135 $X2=0 $Y2=0
cc_7 B N_Y_c_21_n 0.00184579f $X=0.135 $Y=0.152 $X2=0 $Y2=0
cc_8 N_B_M1_g N_Y_c_22_n 2.25474e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_9 B N_Y_c_22_n 0.00374774f $X=0.135 $Y=0.152 $X2=0 $Y2=0
cc_10 N_B_M1_g N_Y_c_20_n 3.14377e-19 $X=0.135 $Y=0.0675 $X2=0.064 $Y2=0.135
cc_11 N_B_c_9_n N_Y_c_25_n 0.00158333f $X=0.135 $Y=0.135 $X2=0.064 $Y2=0.135
cc_12 N_B_c_9_n Y 0.0029629f $X=0.135 $Y=0.135 $X2=0.064 $Y2=0.135
cc_13 N_B_c_9_n N_Y_c_27_n 0.0029629f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 N_B_c_9_n N_6_M1_s 2.67285e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.0675

* END of "./NAND2xp5_ASAP7_75t_R.pex.sp.NAND2XP5_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND2xp67_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:39:50 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND2xp67_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND2xp67_ASAP7_75t_R.pex.sp.pex"
* File: NAND2xp67_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:39:50 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND2XP67_ASAP7_75T_R%A 2 7 10 13 29 VSS
c13 29 VSS 0.0214717f $X=0.081 $Y=0.135
c14 13 VSS 0.00825442f $X=0.135 $Y=0.134
c15 10 VSS 0.0641083f $X=0.135 $Y=0.054
c16 2 VSS 0.067081f $X=0.081 $Y=0.054
r17 10 13 299.72 $w=2e-08 $l=8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.134
r18 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.134 $X2=0.135 $Y2=0.134
r19 5 29 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.134 $X2=0.081
+ $Y2=0.134
r20 5 7 307.213 $w=2e-08 $l=8.2e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.134 $X2=0.081 $Y2=0.216
r21 2 5 299.72 $w=2e-08 $l=8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.134
.ends

.subckt PM_NAND2XP67_ASAP7_75T_R%B 2 7 10 13 22 27 VSS
c23 29 VSS 1.25858e-19 $X=0.243 $Y=0.1495
c24 27 VSS 0.00309799f $X=0.243 $Y=0.156
c25 22 VSS 0.00169371f $X=0.243 $Y=0.135
c26 13 VSS 0.00450327f $X=0.243 $Y=0.134
c27 10 VSS 0.0680265f $X=0.243 $Y=0.054
c28 2 VSS 0.0631829f $X=0.189 $Y=0.054
r29 28 29 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.143 $X2=0.243 $Y2=0.1495
r30 27 29 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.156 $X2=0.243 $Y2=0.1495
r31 22 28 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.143
r32 13 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r33 10 13 299.72 $w=2e-08 $l=8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.134
r34 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.134 $X2=0.243 $Y2=0.134
r35 5 7 307.213 $w=2e-08 $l=8.2e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.134 $X2=0.189 $Y2=0.216
r36 2 5 299.72 $w=2e-08 $l=8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.134
.ends

.subckt PM_NAND2XP67_ASAP7_75T_R%5 1 4 6 7 10 11 14 17 25 26 28 30 32 33 VSS
c18 33 VSS 0.00261791f $X=0.236 $Y=0.036
c19 32 VSS 0.00328455f $X=0.202 $Y=0.036
c20 30 VSS 0.00496337f $X=0.27 $Y=0.036
c21 28 VSS 1.16009e-19 $X=0.1605 $Y=0.036
c22 27 VSS 0.00107916f $X=0.159 $Y=0.036
c23 26 VSS 0.0076767f $X=0.148 $Y=0.036
c24 25 VSS 0.00361761f $X=0.095 $Y=0.036
c25 17 VSS 0.00190391f $X=0.054 $Y=0.036
c26 14 VSS 0.00248078f $X=0.268 $Y=0.054
c27 10 VSS 0.00478875f $X=0.162 $Y=0.054
c28 6 VSS 5.74992e-19 $X=0.179 $Y=0.054
c29 4 VSS 0.0059531f $X=0.056 $Y=0.054
c30 1 VSS 2.6657e-19 $X=0.071 $Y=0.054
r31 32 33 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.036 $X2=0.236 $Y2=0.036
r32 30 33 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.236 $Y2=0.036
r33 27 28 0.101852 $w=1.8e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.159
+ $Y=0.036 $X2=0.1605 $Y2=0.036
r34 26 27 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.036 $X2=0.159 $Y2=0.036
r35 25 26 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.036 $X2=0.148 $Y2=0.036
r36 23 32 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.202 $Y2=0.036
r37 23 28 0.101852 $w=1.8e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.1605 $Y2=0.036
r38 17 25 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.095 $Y2=0.036
r39 14 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r40 11 14 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.054 $X2=0.268 $Y2=0.054
r41 10 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r42 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.162 $Y2=0.054
r43 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.054 $X2=0.162 $Y2=0.054
r44 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r45 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.054 $X2=0.056 $Y2=0.054
.ends

.subckt PM_NAND2XP67_ASAP7_75T_R%Y 1 2 5 6 11 14 18 23 24 30 31 35 37 VSS
c24 39 VSS 5.3979e-19 $X=0.297 $Y=0.216
c25 37 VSS 1.3028e-19 $X=0.297 $Y=0.1025
c26 36 VSS 8.85605e-19 $X=0.297 $Y=0.099
c27 35 VSS 0.00467429f $X=0.298 $Y=0.106
c28 33 VSS 5.09802e-19 $X=0.297 $Y=0.225
c29 31 VSS 4.19287e-19 $X=0.284 $Y=0.072
c30 30 VSS 1.45192e-19 $X=0.252 $Y=0.072
c31 25 VSS 0.00215853f $X=0.288 $Y=0.072
c32 24 VSS 0.0048568f $X=0.252 $Y=0.234
c33 23 VSS 0.00593438f $X=0.215 $Y=0.234
c34 18 VSS 0.00213478f $X=0.162 $Y=0.234
c35 16 VSS 0.00749146f $X=0.288 $Y=0.234
c36 14 VSS 0.0242364f $X=0.164 $Y=0.216
c37 11 VSS 2.6657e-19 $X=0.179 $Y=0.216
c38 9 VSS 3.19801e-19 $X=0.106 $Y=0.216
c39 5 VSS 0.00327684f $X=0.216 $Y=0.054
c40 1 VSS 6.1827e-19 $X=0.233 $Y=0.054
r41 38 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.207 $X2=0.297 $Y2=0.216
r42 36 37 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.099 $X2=0.297 $Y2=0.1025
r43 35 38 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.207
r44 35 37 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.106 $X2=0.297 $Y2=0.1025
r45 33 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.216
r46 32 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.081 $X2=0.297 $Y2=0.099
r47 30 31 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.072 $X2=0.284 $Y2=0.072
r48 27 30 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.072 $X2=0.252 $Y2=0.072
r49 25 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.072 $X2=0.297 $Y2=0.081
r50 25 31 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.284 $Y2=0.072
r51 23 24 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.215
+ $Y=0.234 $X2=0.252 $Y2=0.234
r52 18 23 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.215 $Y2=0.234
r53 16 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.234 $X2=0.297 $Y2=0.225
r54 16 24 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.252 $Y2=0.234
r55 14 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r56 11 14 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.216 $X2=0.164 $Y2=0.216
r57 9 14 21.4815 $w=5.4e-08 $l=5.6e-08 $layer=LISD $thickness=2.8e-08 $X=0.106
+ $Y=0.216 $X2=0.162 $Y2=0.216
r58 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.216 $X2=0.106 $Y2=0.216
r59 5 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072 $X2=0.216
+ $Y2=0.072
r60 2 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.054 $X2=0.216 $Y2=0.054
r61 1 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.054 $X2=0.216 $Y2=0.054
.ends


* END of "./NAND2xp67_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND2xp67_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 VSS N_A_M0_g N_5_M0_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 VSS N_A_M1_g N_5_M1_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_B_M2_g N_5_M2_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.027
M3 N_Y_M3_d N_B_M3_g N_5_M3_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_A_M4_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M5 VDD N_B_M5_g N_Y_M5_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.189
*
* 
* .include "NAND2xp67_ASAP7_75t_R.pex.sp.NAND2XP67_ASAP7_75T_R.pxi"
* BEGIN of "./NAND2xp67_ASAP7_75t_R.pex.sp.NAND2XP67_ASAP7_75T_R.pxi"
* File: NAND2xp67_ASAP7_75t_R.pex.sp.NAND2XP67_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:39:50 2017
* 
x_PM_NAND2XP67_ASAP7_75T_R%A N_A_M0_g N_A_M4_g N_A_M1_g N_A_c_4_p A VSS
+ PM_NAND2XP67_ASAP7_75T_R%A
x_PM_NAND2XP67_ASAP7_75T_R%B N_B_M2_g N_B_M5_g N_B_M3_g N_B_c_17_n N_B_c_18_n B
+ VSS PM_NAND2XP67_ASAP7_75T_R%B
x_PM_NAND2XP67_ASAP7_75T_R%5 N_5_M0_s N_5_c_37_n N_5_M2_s N_5_M1_s N_5_c_47_p
+ N_5_M3_s N_5_c_48_p N_5_c_38_n N_5_c_39_n N_5_c_42_n N_5_c_43_n N_5_c_44_n
+ N_5_c_45_n N_5_c_49_p VSS PM_NAND2XP67_ASAP7_75T_R%5
x_PM_NAND2XP67_ASAP7_75T_R%Y N_Y_M3_d N_Y_M2_d N_Y_c_57_n N_Y_M4_d N_Y_M5_s
+ N_Y_c_55_n N_Y_c_59_n N_Y_c_60_n N_Y_c_63_n N_Y_c_66_n N_Y_c_77_n Y N_Y_c_70_n
+ VSS PM_NAND2XP67_ASAP7_75T_R%Y
cc_1 N_A_M0_g N_B_M2_g 2.60402e-19 $X=0.081 $Y=0.054 $X2=0.189 $Y2=0.054
cc_2 N_A_M1_g N_B_M2_g 0.0035196f $X=0.135 $Y=0.054 $X2=0.189 $Y2=0.054
cc_3 N_A_M1_g N_B_M3_g 2.66145e-19 $X=0.135 $Y=0.054 $X2=0.243 $Y2=0.054
cc_4 N_A_c_4_p N_B_c_17_n 0.00166687f $X=0.135 $Y=0.134 $X2=0.243 $Y2=0.134
cc_5 A N_B_c_18_n 2.96242e-19 $X=0.081 $Y=0.135 $X2=0.243 $Y2=0.135
cc_6 A N_5_c_37_n 0.00127611f $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.134
cc_7 A N_5_c_38_n 0.0013084f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_8 N_A_M0_g N_5_c_39_n 3.94108e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_9 N_A_c_4_p N_5_c_39_n 0.0012051f $X=0.135 $Y=0.134 $X2=0 $Y2=0
cc_10 A N_5_c_39_n 2.8148e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 N_A_M1_g N_5_c_42_n 2.64594e-19 $X=0.135 $Y=0.054 $X2=0.243 $Y2=0.156
cc_12 N_A_M1_g N_Y_c_55_n 0.00417587f $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_13 N_A_c_4_p N_Y_c_55_n 0.00112995f $X=0.135 $Y=0.134 $X2=0 $Y2=0
cc_14 N_B_c_18_n N_5_c_43_n 7.67449e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_15 N_B_M3_g N_5_c_44_n 2.08314e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_16 N_B_M2_g N_5_c_45_n 3.80935e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_17 N_B_c_18_n N_5_c_45_n 7.67449e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_18 N_B_c_17_n N_Y_c_57_n 2.22621e-19 $X=0.243 $Y=0.134 $X2=0.081 $Y2=0.134
cc_19 N_B_c_18_n N_Y_c_57_n 3.67635e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.134
cc_20 N_B_c_18_n N_Y_c_59_n 2.39189e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_21 N_B_M2_g N_Y_c_60_n 4.54533e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_22 N_B_c_17_n N_Y_c_60_n 4.57463e-19 $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_23 N_B_c_18_n N_Y_c_60_n 2.39189e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_24 N_B_M3_g N_Y_c_63_n 2.38524e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_25 N_B_c_18_n N_Y_c_63_n 2.39189e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_26 B N_Y_c_63_n 0.00374293f $X=0.243 $Y=0.156 $X2=0 $Y2=0
cc_27 N_B_M3_g N_Y_c_66_n 2.52075e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_28 N_B_c_18_n N_Y_c_66_n 0.00435317f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_29 N_B_c_17_n Y 3.53802e-19 $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_30 N_B_c_18_n Y 0.00270826f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 N_B_c_18_n N_Y_c_70_n 0.00270826f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_32 N_5_c_47_p N_Y_c_57_n 0.00268053f $X=0.162 $Y=0.054 $X2=0.081 $Y2=0.134
cc_33 N_5_c_48_p N_Y_c_57_n 0.00302498f $X=0.268 $Y=0.054 $X2=0.081 $Y2=0.134
cc_34 N_5_c_49_p N_Y_c_57_n 0.00250906f $X=0.236 $Y=0.036 $X2=0.081 $Y2=0.134
cc_35 N_5_c_47_p N_Y_c_55_n 6.10379e-19 $X=0.162 $Y=0.054 $X2=0 $Y2=0
cc_36 N_5_c_47_p N_Y_c_66_n 5.19937e-19 $X=0.162 $Y=0.054 $X2=0 $Y2=0
cc_37 N_5_c_49_p N_Y_c_66_n 0.00353851f $X=0.236 $Y=0.036 $X2=0 $Y2=0
cc_38 N_5_c_48_p N_Y_c_77_n 0.00418478f $X=0.268 $Y=0.054 $X2=0 $Y2=0
cc_39 N_5_c_44_n N_Y_c_77_n 0.00353851f $X=0.27 $Y=0.036 $X2=0 $Y2=0

* END of "./NAND2xp67_ASAP7_75t_R.pex.sp.NAND2XP67_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND3x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:40:12 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND3x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND3x1_ASAP7_75t_R.pex.sp.pex"
* File: NAND3x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:40:12 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND3X1_ASAP7_75T_R%C 2 8 14 17 19 27 VSS
c9 27 VSS 0.00530818f $X=0.069 $Y=0.137
c10 17 VSS 0.0135792f $X=0.189 $Y=0.135
c11 14 VSS 0.0633654f $X=0.189 $Y=0.0675
c12 8 VSS 0.0651217f $X=0.135 $Y=0.0675
c13 2 VSS 0.0678661f $X=0.081 $Y=0.0675
r14 23 27 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.07 $Y=0.135 $X2=0.07
+ $Y2=0.135
r15 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r16 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r17 11 17 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135 $Y=0.135
+ $X2=0.189 $Y2=0.135
r18 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r19 5 11 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081 $Y=0.135
+ $X2=0.135 $Y2=0.135
r20 5 23 11 $w=2e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.081 $Y=0.135
+ $X2=0.07 $Y2=0.135
r21 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NAND3X1_ASAP7_75T_R%B 2 7 10 16 19 32 VSS
c26 32 VSS 0.00451624f $X=0.296 $Y=0.137
c27 19 VSS 0.00872156f $X=0.351 $Y=0.135
c28 16 VSS 0.0622709f $X=0.351 $Y=0.0675
c29 10 VSS 0.0637068f $X=0.297 $Y=0.0675
c30 2 VSS 0.0632372f $X=0.243 $Y=0.0675
r31 16 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r32 13 19 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297 $Y=0.135
+ $X2=0.351 $Y2=0.135
r33 13 32 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r34 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r35 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243 $Y=0.135
+ $X2=0.297 $Y2=0.135
r36 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r37 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_NAND3X1_ASAP7_75T_R%A 2 7 10 16 19 32 VSS
c25 32 VSS 0.00187217f $X=0.459 $Y=0.137
c26 19 VSS 0.00643044f $X=0.513 $Y=0.135
c27 16 VSS 0.0684308f $X=0.513 $Y=0.0675
c28 10 VSS 0.0645812f $X=0.459 $Y=0.0675
c29 2 VSS 0.0626082f $X=0.405 $Y=0.0675
r30 16 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
r31 13 19 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459 $Y=0.135
+ $X2=0.513 $Y2=0.135
r32 13 32 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r33 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r34 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405 $Y=0.135
+ $X2=0.459 $Y2=0.135
r35 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r36 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_NAND3X1_ASAP7_75T_R%6 1 2 5 6 7 10 11 12 15 23 24 26 28 30 31 VSS
c23 31 VSS 1.29789e-19 $X=0.306 $Y=0.072
c24 30 VSS 4.27727e-19 $X=0.256 $Y=0.072
c25 29 VSS 2.16375e-19 $X=0.246 $Y=0.072
c26 28 VSS 0.00189039f $X=0.243 $Y=0.072
c27 26 VSS 2.61023e-19 $X=0.324 $Y=0.072
c28 24 VSS 0.00103795f $X=0.202 $Y=0.072
c29 23 VSS 0.0109894f $X=0.176 $Y=0.072
c30 15 VSS 0.00275624f $X=0.324 $Y=0.0675
c31 11 VSS 5.7545e-19 $X=0.341 $Y=0.0675
c32 10 VSS 0.00416712f $X=0.216 $Y=0.0675
c33 6 VSS 6.69874e-19 $X=0.233 $Y=0.0675
c34 5 VSS 0.0124244f $X=0.108 $Y=0.0675
c35 1 VSS 6.89902e-19 $X=0.125 $Y=0.0675
r36 30 31 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.072 $X2=0.306 $Y2=0.072
r37 29 30 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.246
+ $Y=0.072 $X2=0.256 $Y2=0.072
r38 28 29 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.072 $X2=0.246 $Y2=0.072
r39 26 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.072 $X2=0.306 $Y2=0.072
r40 23 24 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.072 $X2=0.202 $Y2=0.072
r41 21 28 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.072 $X2=0.243 $Y2=0.072
r42 21 24 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.072 $X2=0.202 $Y2=0.072
r43 17 23 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.176 $Y2=0.072
r44 15 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.072 $X2=0.324
+ $Y2=0.072
r45 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r46 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r47 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072 $X2=0.216
+ $Y2=0.072
r48 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r49 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r50 5 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072 $X2=0.108
+ $Y2=0.072
r51 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r52 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends

.subckt PM_NAND3X1_ASAP7_75T_R%7 1 2 6 7 11 12 18 22 23 24 26 27 29 VSS
c26 29 VSS 0.00146166f $X=0.418 $Y=0.036
c27 28 VSS 0.00440359f $X=0.4 $Y=0.036
c28 27 VSS 0.00269882f $X=0.486 $Y=0.036
c29 26 VSS 0.00696613f $X=0.486 $Y=0.036
c30 24 VSS 0.00193338f $X=0.358 $Y=0.036
c31 23 VSS 0.00716859f $X=0.338 $Y=0.036
c32 22 VSS 0.00329808f $X=0.378 $Y=0.036
c33 18 VSS 0.00452674f $X=0.27 $Y=0.036
c34 11 VSS 6.4978e-19 $X=0.503 $Y=0.0675
c35 6 VSS 5.38922e-19 $X=0.395 $Y=0.0675
c36 1 VSS 7.48473e-19 $X=0.287 $Y=0.0675
r37 28 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.4
+ $Y=0.036 $X2=0.418 $Y2=0.036
r38 26 29 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.418 $Y2=0.036
r39 26 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036 $X2=0.486
+ $Y2=0.036
r40 23 24 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.036 $X2=0.358 $Y2=0.036
r41 21 28 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.4 $Y2=0.036
r42 21 24 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.358 $Y2=0.036
r43 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r44 17 23 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.338 $Y2=0.036
r45 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r46 15 27 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0675 $X2=0.486 $Y2=0.036
r47 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.486 $Y2=0.0675
r48 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.0675 $X2=0.486 $Y2=0.0675
r49 10 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r50 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.378 $Y2=0.0675
r51 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.0675 $X2=0.378 $Y2=0.0675
r52 5 18 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r53 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
r54 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends

.subckt PM_NAND3X1_ASAP7_75T_R%Y 1 2 5 6 9 11 12 15 16 19 21 29 30 31 32 34 35
+ 36 37 45 46 50 52 VSS
c33 54 VSS 6.71881e-19 $X=0.567 $Y=0.2115
c34 52 VSS 0.00103607f $X=0.567 $Y=0.1255
c35 51 VSS 0.00118799f $X=0.567 $Y=0.108
c36 50 VSS 0.00346075f $X=0.566 $Y=0.143
c37 48 VSS 7.79697e-19 $X=0.567 $Y=0.225
c38 46 VSS 2.77631e-19 $X=0.5 $Y=0.072
c39 45 VSS 8.6783e-20 $X=0.468 $Y=0.072
c40 37 VSS 0.00420063f $X=0.558 $Y=0.072
c41 36 VSS 0.00414532f $X=0.513 $Y=0.234
c42 35 VSS 0.00397796f $X=0.468 $Y=0.234
c43 34 VSS 0.00141093f $X=0.417 $Y=0.234
c44 33 VSS 2.01672e-19 $X=0.402 $Y=0.234
c45 32 VSS 0.00915231f $X=0.4 $Y=0.234
c46 31 VSS 0.00312606f $X=0.338 $Y=0.234
c47 30 VSS 0.0083386f $X=0.306 $Y=0.234
c48 29 VSS 0.0052167f $X=0.243 $Y=0.234
c49 21 VSS 0.00782805f $X=0.558 $Y=0.234
c50 19 VSS 0.00719327f $X=0.43 $Y=0.2025
c51 15 VSS 0.00963529f $X=0.216 $Y=0.2025
c52 11 VSS 5.72268e-19 $X=0.233 $Y=0.2025
c53 9 VSS 0.00107488f $X=0.538 $Y=0.0675
c54 5 VSS 0.00286008f $X=0.432 $Y=0.0675
c55 1 VSS 6.95637e-19 $X=0.449 $Y=0.0675
r56 53 54 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.198 $X2=0.567 $Y2=0.2115
r57 51 52 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.108 $X2=0.567 $Y2=0.1255
r58 50 53 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.143 $X2=0.567 $Y2=0.198
r59 50 52 1.18827 $w=1.8e-08 $l=1.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.143 $X2=0.567 $Y2=0.1255
r60 48 54 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.225 $X2=0.567 $Y2=0.2115
r61 47 51 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.567 $Y2=0.108
r62 45 46 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.072 $X2=0.5 $Y2=0.072
r63 43 46 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.072 $X2=0.5 $Y2=0.072
r64 39 45 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.072 $X2=0.468 $Y2=0.072
r65 37 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.072 $X2=0.567 $Y2=0.081
r66 37 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.072 $X2=0.54 $Y2=0.072
r67 35 36 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.513 $Y2=0.234
r68 33 34 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.402
+ $Y=0.234 $X2=0.417 $Y2=0.234
r69 32 33 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.4
+ $Y=0.234 $X2=0.402 $Y2=0.234
r70 31 32 4.20988 $w=1.8e-08 $l=6.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.234 $X2=0.4 $Y2=0.234
r71 30 31 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.338 $Y2=0.234
r72 29 30 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.234 $X2=0.306 $Y2=0.234
r73 27 35 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.468 $Y2=0.234
r74 27 34 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.417 $Y2=0.234
r75 23 29 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.243 $Y2=0.234
r76 21 48 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.234 $X2=0.567 $Y2=0.225
r77 21 36 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.513 $Y2=0.234
r78 19 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r79 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.43 $Y2=0.2025
r80 15 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r81 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r82 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r83 9 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.072 $X2=0.54
+ $Y2=0.072
r84 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.523
+ $Y=0.0675 $X2=0.538 $Y2=0.0675
r85 5 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.072 $X2=0.432
+ $Y2=0.072
r86 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.432 $Y2=0.0675
r87 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.449
+ $Y=0.0675 $X2=0.432 $Y2=0.0675
.ends


* END of "./NAND3x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND3x1_ASAP7_75t_R  VSS VDD C B A Y
* 
* Y	Y
* A	A
* B	B
* C	C
M0 N_6_M0_d N_C_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_6_M1_d N_C_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_6_M2_d N_C_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_7_M3_d N_B_M3_g N_6_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_7_M4_d N_B_M4_g N_6_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 N_7_M5_d N_B_M5_g N_6_M5_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 N_Y_M6_d N_A_M6_g N_7_M6_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_Y_M7_d N_A_M7_g N_7_M7_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_Y_M8_d N_A_M8_g N_7_M8_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 N_Y_M9_d N_C_M9_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M10 VDD N_B_M10_g N_Y_M10_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M11 N_Y_M11_d N_A_M11_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
*
* 
* .include "NAND3x1_ASAP7_75t_R.pex.sp.NAND3X1_ASAP7_75T_R.pxi"
* BEGIN of "./NAND3x1_ASAP7_75t_R.pex.sp.NAND3X1_ASAP7_75T_R.pxi"
* File: NAND3x1_ASAP7_75t_R.pex.sp.NAND3X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:40:12 2017
* 
x_PM_NAND3X1_ASAP7_75T_R%C N_C_M0_g N_C_M1_g N_C_M2_g N_C_c_4_p N_C_M9_g C VSS
+ PM_NAND3X1_ASAP7_75T_R%C
x_PM_NAND3X1_ASAP7_75T_R%B N_B_M3_g N_B_M10_g N_B_M4_g N_B_M5_g N_B_c_13_n B VSS
+ PM_NAND3X1_ASAP7_75T_R%B
x_PM_NAND3X1_ASAP7_75T_R%A N_A_M6_g N_A_M11_g N_A_M7_g N_A_M8_g N_A_c_39_n A VSS
+ PM_NAND3X1_ASAP7_75T_R%A
x_PM_NAND3X1_ASAP7_75T_R%6 N_6_M1_d N_6_M0_d N_6_c_62_n N_6_M3_s N_6_M2_d
+ N_6_c_72_p N_6_M5_s N_6_M4_s N_6_c_67_n N_6_c_63_n N_6_c_65_n N_6_c_68_n
+ N_6_c_69_n N_6_c_70_n N_6_c_71_n VSS PM_NAND3X1_ASAP7_75T_R%6
x_PM_NAND3X1_ASAP7_75T_R%7 N_7_M4_d N_7_M3_d N_7_M6_s N_7_M5_d N_7_M8_s N_7_M7_s
+ N_7_c_85_n N_7_c_97_n N_7_c_86_n N_7_c_87_n N_7_c_90_n N_7_c_91_n N_7_c_92_n
+ VSS PM_NAND3X1_ASAP7_75T_R%7
x_PM_NAND3X1_ASAP7_75T_R%Y N_Y_M7_d N_Y_M6_d N_Y_c_117_n N_Y_M8_d N_Y_c_138_n
+ N_Y_M10_s N_Y_M9_d N_Y_c_110_n N_Y_M11_d N_Y_c_118_n N_Y_c_120_n N_Y_c_111_n
+ N_Y_c_112_n N_Y_c_114_n N_Y_c_115_n N_Y_c_121_n N_Y_c_122_n N_Y_c_123_n
+ N_Y_c_125_n N_Y_c_126_n N_Y_c_128_n Y N_Y_c_130_n VSS PM_NAND3X1_ASAP7_75T_R%Y
cc_1 N_C_M1_g N_B_M3_g 2.71887e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_2 N_C_M2_g N_B_M3_g 0.00357042f $X=0.189 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_3 N_C_M2_g N_B_M4_g 2.71887e-19 $X=0.189 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_4 N_C_c_4_p N_B_c_13_n 0.00175803f $X=0.189 $Y=0.135 $X2=0.351 $Y2=0.135
cc_5 N_C_c_4_p N_6_M1_d 3.67575e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_6 N_C_c_4_p N_6_c_62_n 0.00203185f $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.135
cc_7 N_C_M1_g N_6_c_63_n 3.91767e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_8 N_C_c_4_p N_6_c_63_n 0.00173937f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_9 N_C_M2_g N_6_c_65_n 4.87149e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_10 N_B_M4_g N_A_M6_g 2.71887e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_11 N_B_M5_g N_A_M6_g 0.00333077f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_12 N_B_M5_g N_A_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_13 N_B_c_13_n N_A_c_39_n 0.00160961f $X=0.351 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_14 B A 9.49045e-19 $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_15 N_B_c_13_n N_6_M5_s 3.67575e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_16 N_B_c_13_n N_6_c_67_n 0.00203185f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_17 N_B_c_13_n N_6_c_68_n 4.94606e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_18 N_B_M3_g N_6_c_69_n 2.42055e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_19 B N_6_c_70_n 0.00387635f $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_20 N_B_M4_g N_6_c_71_n 2.82354e-19 $X=0.297 $Y=0.0675 $X2=0.07 $Y2=0.135
cc_21 N_B_c_13_n N_7_M4_d 3.1125e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_22 N_B_c_13_n N_7_c_85_n 7.57503e-19 $X=0.351 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_23 N_B_M4_g N_7_c_86_n 2.38524e-19 $X=0.297 $Y=0.0675 $X2=0.07 $Y2=0.135
cc_24 N_B_M5_g N_7_c_87_n 3.92012e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_25 N_B_c_13_n N_7_c_87_n 2.49103e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_26 B N_Y_c_110_n 5.84163e-19 $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_27 N_B_M3_g N_Y_c_111_n 2.26704e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_28 N_B_M4_g N_Y_c_112_n 2.71534e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_29 B N_Y_c_112_n 0.00407548f $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_30 N_B_c_13_n N_Y_c_114_n 4.93209e-19 $X=0.351 $Y=0.135 $X2=0.07 $Y2=0.135
cc_31 N_B_M5_g N_Y_c_115_n 4.61191e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_32 N_A_c_39_n N_7_M8_s 3.67193e-19 $X=0.513 $Y=0.135 $X2=0.135 $Y2=0.135
cc_33 N_A_M7_g N_7_c_90_n 2.38524e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_34 N_A_c_39_n N_7_c_91_n 0.00203185f $X=0.513 $Y=0.135 $X2=0.069 $Y2=0.137
cc_35 N_A_M6_g N_7_c_92_n 3.01362e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_36 A N_7_c_92_n 5.94322e-19 $X=0.459 $Y=0.137 $X2=0 $Y2=0
cc_37 N_A_c_39_n N_Y_M7_d 3.03469e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_38 N_A_c_39_n N_Y_c_117_n 7.57503e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.135
cc_39 N_A_c_39_n N_Y_c_118_n 7.57503e-19 $X=0.513 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_40 A N_Y_c_118_n 0.00236517f $X=0.459 $Y=0.137 $X2=0.189 $Y2=0.2025
cc_41 N_A_M8_g N_Y_c_120_n 2.70934e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_42 A N_Y_c_121_n 0.0042539f $X=0.459 $Y=0.137 $X2=0.135 $Y2=0.135
cc_43 N_A_M7_g N_Y_c_122_n 2.67763e-19 $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.135
cc_44 N_A_M8_g N_Y_c_123_n 2.77881e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_45 N_A_c_39_n N_Y_c_123_n 4.7342e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_46 N_A_M8_g N_Y_c_125_n 4.944e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_A_M7_g N_Y_c_126_n 2.78432e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_48 A N_Y_c_126_n 0.0030377f $X=0.459 $Y=0.137 $X2=0 $Y2=0
cc_49 N_A_c_39_n N_Y_c_128_n 8.63627e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_50 A Y 9.2038e-19 $X=0.459 $Y=0.137 $X2=0 $Y2=0
cc_51 A N_Y_c_130_n 9.2038e-19 $X=0.459 $Y=0.137 $X2=0 $Y2=0
cc_52 N_6_c_72_p N_7_c_85_n 0.00318646f $X=0.216 $Y=0.0675 $X2=0.189 $Y2=0.2025
cc_53 N_6_c_67_n N_7_c_85_n 0.00350522f $X=0.324 $Y=0.0675 $X2=0.189 $Y2=0.2025
cc_54 N_6_c_71_n N_7_c_85_n 0.00206264f $X=0.306 $Y=0.072 $X2=0.189 $Y2=0.2025
cc_55 N_6_c_67_n N_7_c_97_n 0.00328789f $X=0.324 $Y=0.0675 $X2=0.07 $Y2=0.135
cc_56 N_6_c_68_n N_7_c_97_n 4.49606e-19 $X=0.324 $Y=0.072 $X2=0.07 $Y2=0.135
cc_57 N_6_c_72_p N_7_c_86_n 4.49606e-19 $X=0.216 $Y=0.0675 $X2=0.07 $Y2=0.135
cc_58 N_6_c_67_n N_7_c_86_n 0.00250914f $X=0.324 $Y=0.0675 $X2=0.07 $Y2=0.135
cc_59 N_6_c_71_n N_7_c_86_n 0.00704516f $X=0.306 $Y=0.072 $X2=0.07 $Y2=0.135
cc_60 N_6_c_72_p N_Y_c_110_n 0.00138157f $X=0.216 $Y=0.0675 $X2=0 $Y2=0
cc_61 N_6_c_69_n N_Y_c_111_n 2.6332e-19 $X=0.243 $Y=0.072 $X2=0 $Y2=0
cc_62 N_6_c_68_n N_Y_c_114_n 2.6332e-19 $X=0.324 $Y=0.072 $X2=0.07 $Y2=0.135
cc_63 N_6_c_68_n N_Y_c_126_n 3.04405e-19 $X=0.324 $Y=0.072 $X2=0 $Y2=0
cc_64 N_7_c_97_n N_Y_c_117_n 0.00328788f $X=0.378 $Y=0.036 $X2=0.243 $Y2=0.135
cc_65 N_7_c_90_n N_Y_c_117_n 0.00250914f $X=0.486 $Y=0.036 $X2=0.243 $Y2=0.135
cc_66 N_7_c_91_n N_Y_c_117_n 0.00350515f $X=0.486 $Y=0.036 $X2=0.243 $Y2=0.135
cc_67 N_7_c_90_n N_Y_c_138_n 3.09693e-19 $X=0.486 $Y=0.036 $X2=0.297 $Y2=0.0675
cc_68 N_7_c_91_n N_Y_c_138_n 0.00337028f $X=0.486 $Y=0.036 $X2=0.297 $Y2=0.0675
cc_69 N_7_c_97_n N_Y_c_126_n 4.51951e-19 $X=0.378 $Y=0.036 $X2=0 $Y2=0
cc_70 N_7_c_90_n N_Y_c_126_n 0.00704516f $X=0.486 $Y=0.036 $X2=0 $Y2=0
cc_71 N_7_c_91_n N_Y_c_128_n 0.00233206f $X=0.486 $Y=0.036 $X2=0 $Y2=0

* END of "./NAND3x1_ASAP7_75t_R.pex.sp.NAND3X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND3x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:40:35 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND3x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND3x2_ASAP7_75t_R.pex.sp.pex"
* File: NAND3x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:40:35 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND3X2_ASAP7_75T_R%A 2 8 14 17 19 22 27 30 36 39 43 48 53 57 58 VSS
c69 58 VSS 0.0251808f $X=0.894 $Y=0.192
c70 57 VSS 0.00174297f $X=0.894 $Y=0.189
c71 53 VSS 0.00185559f $X=0.183 $Y=0.189
c72 48 VSS 0.00258491f $X=0.894 $Y=0.135
c73 43 VSS 0.00231474f $X=0.183 $Y=0.135
c74 39 VSS 0.00589537f $X=0.999 $Y=0.135
c75 36 VSS 0.0684487f $X=0.999 $Y=0.0675
c76 30 VSS 0.0649556f $X=0.945 $Y=0.0675
c77 22 VSS 0.0621952f $X=0.891 $Y=0.0675
c78 17 VSS 0.00595222f $X=0.189 $Y=0.135
c79 14 VSS 0.0623361f $X=0.189 $Y=0.0675
c80 8 VSS 0.0649686f $X=0.135 $Y=0.0675
c81 2 VSS 0.0684308f $X=0.081 $Y=0.0675
r82 57 58 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.894 $Y=0.189 $X2=0.894
+ $Y2=0.189
r83 52 58 48.2778 $w=1.8e-08 $l=7.11e-07 $layer=M2 $thickness=3.6e-08 $X=0.183
+ $Y=0.189 $X2=0.894 $Y2=0.189
r84 52 53 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.183 $Y=0.189 $X2=0.183
+ $Y2=0.189
r85 48 57 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.894
+ $Y=0.135 $X2=0.894 $Y2=0.189
r86 43 53 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.183
+ $Y=0.135 $X2=0.183 $Y2=0.189
r87 36 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.0675 $X2=0.999 $Y2=0.135
r88 33 39 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.945 $Y=0.135
+ $X2=0.999 $Y2=0.135
r89 30 33 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.945
+ $Y=0.0675 $X2=0.945 $Y2=0.135
r90 25 33 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.891 $Y=0.135
+ $X2=0.945 $Y2=0.135
r91 25 48 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.894 $Y=0.135 $X2=0.894
+ $Y2=0.135
r92 25 27 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.135 $X2=0.891 $Y2=0.2025
r93 22 25 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.0675 $X2=0.891 $Y2=0.135
r94 17 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.183 $Y=0.135 $X2=0.183
+ $Y2=0.135
r95 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r96 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r97 11 17 48 $w=2e-08 $l=4.8e-08 $layer=LIG $thickness=5e-08 $X=0.135 $Y=0.135
+ $X2=0.183 $Y2=0.135
r98 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r99 5 11 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081 $Y=0.135
+ $X2=0.135 $Y2=0.135
r100 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NAND3X2_ASAP7_75T_R%B 2 8 14 17 19 22 27 30 36 39 41 46 49 50 51 52
+ 53 55 VSS
c75 61 VSS 6.87363e-19 $X=0.734 $Y=0.1765
c76 55 VSS 0.00132227f $X=0.734 $Y=0.135
c77 53 VSS 5.96199e-19 $X=0.734 $Y=0.189
c78 52 VSS 3.49249e-19 $X=0.565 $Y=0.198
c79 51 VSS 0.00481358f $X=0.547 $Y=0.198
c80 50 VSS 9.15736e-19 $X=0.356 $Y=0.198
c81 49 VSS 0.00513351f $X=0.725 $Y=0.198
c82 48 VSS 6.87178e-19 $X=0.347 $Y=0.1765
c83 46 VSS 0.00124117f $X=0.348 $Y=0.137
c84 41 VSS 5.90119e-19 $X=0.347 $Y=0.189
c85 39 VSS 0.00836222f $X=0.837 $Y=0.135
c86 36 VSS 0.0622709f $X=0.837 $Y=0.0675
c87 30 VSS 0.0640963f $X=0.783 $Y=0.0675
c88 22 VSS 0.0630165f $X=0.729 $Y=0.0675
c89 17 VSS 0.00834409f $X=0.351 $Y=0.135
c90 14 VSS 0.0629776f $X=0.351 $Y=0.0675
c91 8 VSS 0.0640813f $X=0.297 $Y=0.0675
c92 2 VSS 0.0622537f $X=0.243 $Y=0.0675
r93 60 61 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.734
+ $Y=0.164 $X2=0.734 $Y2=0.1765
r94 55 60 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.734
+ $Y=0.135 $X2=0.734 $Y2=0.164
r95 53 61 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.734
+ $Y=0.189 $X2=0.734 $Y2=0.1765
r96 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.547
+ $Y=0.198 $X2=0.565 $Y2=0.198
r97 50 51 12.9691 $w=1.8e-08 $l=1.91e-07 $layer=M1 $thickness=3.6e-08 $X=0.356
+ $Y=0.198 $X2=0.547 $Y2=0.198
r98 49 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.725 $Y=0.198 $X2=0.734 $Y2=0.189
r99 49 52 10.8642 $w=1.8e-08 $l=1.6e-07 $layer=M1 $thickness=3.6e-08 $X=0.725
+ $Y=0.198 $X2=0.565 $Y2=0.198
r100 47 48 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.347
+ $Y=0.164 $X2=0.347 $Y2=0.1765
r101 46 47 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.347
+ $Y=0.135 $X2=0.347 $Y2=0.164
r102 41 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.347 $Y=0.189 $X2=0.356 $Y2=0.198
r103 41 48 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.347
+ $Y=0.189 $X2=0.347 $Y2=0.1765
r104 36 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.0675 $X2=0.837 $Y2=0.135
r105 33 39 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.783 $Y=0.135
+ $X2=0.837 $Y2=0.135
r106 30 33 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.135
r107 25 33 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729 $Y=0.135
+ $X2=0.783 $Y2=0.135
r108 25 55 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.734 $Y=0.135 $X2=0.734
+ $Y2=0.135
r109 25 27 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.135 $X2=0.729 $Y2=0.2025
r110 22 25 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.135
r111 17 46 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.347 $Y=0.135 $X2=0.347
+ $Y2=0.135
r112 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r113 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r114 11 17 50 $w=2e-08 $l=5e-08 $layer=LIG $thickness=5e-08 $X=0.297 $Y=0.135
+ $X2=0.347 $Y2=0.135
r115 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r116 5 11 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243 $Y=0.135
+ $X2=0.297 $Y2=0.135
r117 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_NAND3X2_ASAP7_75T_R%C 2 7 10 16 22 28 34 37 39 45 VSS
c41 45 VSS 0.00152202f $X=0.555 $Y=0.137
c42 37 VSS 0.0203793f $X=0.675 $Y=0.135
c43 34 VSS 0.062961f $X=0.675 $Y=0.0675
c44 28 VSS 0.0644377f $X=0.621 $Y=0.0675
c45 22 VSS 0.0653595f $X=0.567 $Y=0.0675
c46 16 VSS 0.06505f $X=0.513 $Y=0.0675
c47 10 VSS 0.0644495f $X=0.459 $Y=0.0675
c48 2 VSS 0.0629441f $X=0.405 $Y=0.0675
r49 43 45 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.556 $Y=0.135 $X2=0.556
+ $Y2=0.135
r50 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.2025
r51 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0675 $X2=0.675 $Y2=0.135
r52 31 37 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621 $Y=0.135
+ $X2=0.675 $Y2=0.135
r53 28 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
r54 25 31 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.567 $Y=0.135
+ $X2=0.621 $Y2=0.135
r55 25 43 11 $w=2e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.567 $Y=0.135
+ $X2=0.556 $Y2=0.135
r56 22 25 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r57 19 43 43 $w=2e-08 $l=4.3e-08 $layer=LIG $thickness=5e-08 $X=0.513 $Y=0.135
+ $X2=0.556 $Y2=0.135
r58 16 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
r59 13 19 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459 $Y=0.135
+ $X2=0.513 $Y2=0.135
r60 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r61 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405 $Y=0.135
+ $X2=0.459 $Y2=0.135
r62 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r63 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_NAND3X2_ASAP7_75T_R%6 1 2 6 7 11 12 18 22 23 24 25 28 29 30 31 VSS
c27 31 VSS 0.00267306f $X=0.29 $Y=0.036
c28 30 VSS 0.00383338f $X=0.256 $Y=0.036
c29 29 VSS 0.00475672f $X=0.324 $Y=0.036
c30 28 VSS 0.00453277f $X=0.324 $Y=0.036
c31 26 VSS 3.19325e-19 $X=0.2135 $Y=0.036
c32 25 VSS 0.00193913f $X=0.211 $Y=0.036
c33 24 VSS 0.00130548f $X=0.192 $Y=0.036
c34 23 VSS 0.00695592f $X=0.176 $Y=0.036
c35 22 VSS 0.00347287f $X=0.216 $Y=0.036
c36 18 VSS 0.00269882f $X=0.108 $Y=0.036
c37 11 VSS 7.17878e-19 $X=0.341 $Y=0.0675
c38 6 VSS 5.38922e-19 $X=0.233 $Y=0.0675
c39 1 VSS 6.4978e-19 $X=0.125 $Y=0.0675
r40 30 31 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.036 $X2=0.29 $Y2=0.036
r41 28 31 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.29 $Y2=0.036
r42 28 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r43 25 26 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.211
+ $Y=0.036 $X2=0.2135 $Y2=0.036
r44 24 25 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.192
+ $Y=0.036 $X2=0.211 $Y2=0.036
r45 23 24 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.036 $X2=0.192 $Y2=0.036
r46 21 30 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.256 $Y2=0.036
r47 21 26 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.2135 $Y2=0.036
r48 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r49 17 23 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.176 $Y2=0.036
r50 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r51 15 29 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r52 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r53 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r54 10 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r55 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r56 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r57 5 18 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r58 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r59 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends

.subckt PM_NAND3X2_ASAP7_75T_R%7 1 2 5 6 7 10 11 12 15 16 17 20 21 22 25 26 27
+ 30 38 39 43 48 49 53 54 56 59 61 VSS
c53 61 VSS 2.78809e-19 $X=0.7765 $Y=0.072
c54 59 VSS 5.17444e-19 $X=0.742 $Y=0.072
c55 58 VSS 0.00203085f $X=0.725 $Y=0.072
c56 56 VSS 2.97451e-19 $X=0.81 $Y=0.072
c57 54 VSS 7.11849e-19 $X=0.682 $Y=0.072
c58 53 VSS 0.0106025f $X=0.662 $Y=0.072
c59 49 VSS 0.00240114f $X=0.565 $Y=0.072
c60 48 VSS 0.00978135f $X=0.547 $Y=0.072
c61 44 VSS 0.0051489f $X=0.452 $Y=0.072
c62 43 VSS 0.00262736f $X=0.418 $Y=0.072
c63 39 VSS 5.46526e-19 $X=0.356 $Y=0.072
c64 38 VSS 5.72503e-19 $X=0.338 $Y=0.072
c65 30 VSS 0.0027527f $X=0.81 $Y=0.0675
c66 26 VSS 5.75435e-19 $X=0.827 $Y=0.0675
c67 25 VSS 0.0043741f $X=0.702 $Y=0.0675
c68 21 VSS 6.69874e-19 $X=0.719 $Y=0.0675
c69 20 VSS 0.0125184f $X=0.594 $Y=0.0675
c70 16 VSS 6.05897e-19 $X=0.611 $Y=0.0675
c71 15 VSS 0.0124222f $X=0.486 $Y=0.0675
c72 11 VSS 6.05897e-19 $X=0.503 $Y=0.0675
c73 10 VSS 0.00438003f $X=0.378 $Y=0.0675
c74 6 VSS 6.69874e-19 $X=0.395 $Y=0.0675
c75 5 VSS 0.00274973f $X=0.27 $Y=0.0675
c76 1 VSS 5.76015e-19 $X=0.287 $Y=0.0675
r77 60 61 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.743
+ $Y=0.072 $X2=0.7765 $Y2=0.072
r78 59 60 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.742
+ $Y=0.072 $X2=0.743 $Y2=0.072
r79 58 59 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.725
+ $Y=0.072 $X2=0.742 $Y2=0.072
r80 56 61 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.072 $X2=0.7765 $Y2=0.072
r81 53 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.662
+ $Y=0.072 $X2=0.682 $Y2=0.072
r82 51 58 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.072 $X2=0.725 $Y2=0.072
r83 51 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.072 $X2=0.682 $Y2=0.072
r84 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.547
+ $Y=0.072 $X2=0.565 $Y2=0.072
r85 46 53 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.072 $X2=0.662 $Y2=0.072
r86 46 49 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.072 $X2=0.565 $Y2=0.072
r87 43 44 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.072 $X2=0.452 $Y2=0.072
r88 41 48 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.072 $X2=0.547 $Y2=0.072
r89 41 44 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.072 $X2=0.452 $Y2=0.072
r90 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.072 $X2=0.356 $Y2=0.072
r91 36 43 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.418 $Y2=0.072
r92 36 39 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.356 $Y2=0.072
r93 32 38 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.072 $X2=0.338 $Y2=0.072
r94 30 56 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.072 $X2=0.81
+ $Y2=0.072
r95 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.0675 $X2=0.81 $Y2=0.0675
r96 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.0675 $X2=0.81 $Y2=0.0675
r97 25 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.072 $X2=0.702
+ $Y2=0.072
r98 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.0675 $X2=0.702 $Y2=0.0675
r99 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.0675 $X2=0.702 $Y2=0.0675
r100 20 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.072
+ $X2=0.594 $Y2=0.072
r101 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0675 $X2=0.594 $Y2=0.0675
r102 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0675 $X2=0.594 $Y2=0.0675
r103 15 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.072
+ $X2=0.486 $Y2=0.072
r104 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.486 $Y2=0.0675
r105 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.0675 $X2=0.486 $Y2=0.0675
r106 10 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.072
+ $X2=0.378 $Y2=0.072
r107 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.378 $Y2=0.0675
r108 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.0675 $X2=0.378 $Y2=0.0675
r109 5 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.072 $X2=0.27
+ $Y2=0.072
r110 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r111 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends

.subckt PM_NAND3X2_ASAP7_75T_R%8 1 2 6 7 11 12 18 22 23 24 26 27 30 VSS
c27 31 VSS 1.63466e-19 $X=0.904 $Y=0.036
c28 30 VSS 0.00140825f $X=0.903 $Y=0.036
c29 29 VSS 0.00181697f $X=0.885 $Y=0.036
c30 28 VSS 0.00201427f $X=0.866 $Y=0.036
c31 27 VSS 0.00269882f $X=0.972 $Y=0.036
c32 26 VSS 0.00696456f $X=0.972 $Y=0.036
c33 24 VSS 0.00181142f $X=0.844 $Y=0.036
c34 23 VSS 0.00715189f $X=0.824 $Y=0.036
c35 22 VSS 0.00341054f $X=0.864 $Y=0.036
c36 18 VSS 0.00471687f $X=0.756 $Y=0.036
c37 11 VSS 6.48198e-19 $X=0.989 $Y=0.0675
c38 6 VSS 5.38922e-19 $X=0.881 $Y=0.0675
c39 1 VSS 7.13194e-19 $X=0.773 $Y=0.0675
r40 30 31 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.903
+ $Y=0.036 $X2=0.904 $Y2=0.036
r41 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.885
+ $Y=0.036 $X2=0.903 $Y2=0.036
r42 28 29 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.866
+ $Y=0.036 $X2=0.885 $Y2=0.036
r43 26 31 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.036 $X2=0.904 $Y2=0.036
r44 26 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.036 $X2=0.972
+ $Y2=0.036
r45 23 24 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.824
+ $Y=0.036 $X2=0.844 $Y2=0.036
r46 21 28 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.866 $Y2=0.036
r47 21 24 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.036 $X2=0.844 $Y2=0.036
r48 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.036 $X2=0.864
+ $Y2=0.036
r49 17 23 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.824 $Y2=0.036
r50 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r51 15 27 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.972
+ $Y=0.0675 $X2=0.972 $Y2=0.036
r52 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.0675 $X2=0.972 $Y2=0.0675
r53 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.989 $Y=0.0675 $X2=0.972 $Y2=0.0675
r54 10 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.864
+ $Y=0.0675 $X2=0.864 $Y2=0.036
r55 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.0675 $X2=0.864 $Y2=0.0675
r56 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.0675 $X2=0.864 $Y2=0.0675
r57 5 18 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.756
+ $Y=0.0675 $X2=0.756 $Y2=0.036
r58 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
r59 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
.ends

.subckt PM_NAND3X2_ASAP7_75T_R%Y 1 4 6 7 10 11 12 15 16 19 21 24 26 27 30 31 32
+ 35 36 39 44 50 52 53 56 64 65 66 67 74 75 76 77 79 88 89 93 VSS
c76 97 VSS 4.87068e-19 $X=1.053 $Y=0.216
c77 95 VSS 6.6224e-20 $X=1.053 $Y=0.108
c78 94 VSS 0.00101778f $X=1.053 $Y=0.106
c79 93 VSS 0.00525814f $X=1.052 $Y=0.143
c80 91 VSS 4.60009e-19 $X=1.053 $Y=0.225
c81 89 VSS 7.12898e-19 $X=1.006 $Y=0.072
c82 88 VSS 6.13025e-19 $X=0.986 $Y=0.072
c83 80 VSS 0.00405642f $X=1.044 $Y=0.072
c84 79 VSS 6.76809e-19 $X=0.911 $Y=0.234
c85 77 VSS 0.00409443f $X=0.903 $Y=0.234
c86 76 VSS 0.00578947f $X=0.866 $Y=0.234
c87 75 VSS 0.0103422f $X=0.824 $Y=0.234
c88 74 VSS 0.0385756f $X=0.743 $Y=0.234
c89 67 VSS 0.0103888f $X=0.338 $Y=0.234
c90 66 VSS 0.00631091f $X=0.256 $Y=0.234
c91 65 VSS 0.00389671f $X=0.211 $Y=0.234
c92 64 VSS 0.0126481f $X=0.174 $Y=0.234
c93 57 VSS 0.00354522f $X=0.036 $Y=0.234
c94 56 VSS 0.0156892f $X=1.044 $Y=0.234
c95 53 VSS 3.04498e-19 $X=0.128 $Y=0.072
c96 52 VSS 0.00279066f $X=0.094 $Y=0.072
c97 50 VSS 4.5381e-19 $X=0.162 $Y=0.072
c98 45 VSS 0.0019505f $X=0.036 $Y=0.072
c99 44 VSS 0.00534065f $X=0.027 $Y=0.207
c100 43 VSS 0.00101778f $X=0.027 $Y=0.106
c101 42 VSS 9.47077e-19 $X=0.027 $Y=0.225
c102 39 VSS 0.00749008f $X=0.916 $Y=0.2025
c103 35 VSS 0.0105087f $X=0.702 $Y=0.2025
c104 31 VSS 5.97768e-19 $X=0.719 $Y=0.2025
c105 30 VSS 0.0106828f $X=0.378 $Y=0.2025
c106 26 VSS 5.97768e-19 $X=0.395 $Y=0.2025
c107 24 VSS 0.00716926f $X=0.164 $Y=0.2025
c108 21 VSS 5.4394e-19 $X=0.179 $Y=0.2025
c109 19 VSS 0.00107488f $X=1.024 $Y=0.0675
c110 15 VSS 0.0027527f $X=0.918 $Y=0.0675
c111 11 VSS 5.9588e-19 $X=0.935 $Y=0.0675
c112 10 VSS 0.00278521f $X=0.162 $Y=0.0675
c113 6 VSS 6.95677e-19 $X=0.179 $Y=0.0675
c114 4 VSS 7.39942e-19 $X=0.056 $Y=0.0675
c115 1 VSS 3.34937e-19 $X=0.071 $Y=0.0675
r116 96 97 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.207 $X2=1.053 $Y2=0.216
r117 94 95 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.106 $X2=1.053 $Y2=0.108
r118 93 96 4.34568 $w=1.8e-08 $l=6.4e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.143 $X2=1.053 $Y2=0.207
r119 93 95 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.143 $X2=1.053 $Y2=0.108
r120 91 97 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.225 $X2=1.053 $Y2=0.216
r121 90 94 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.081 $X2=1.053 $Y2=0.106
r122 88 89 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.986
+ $Y=0.072 $X2=1.006 $Y2=0.072
r123 86 89 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.072 $X2=1.006 $Y2=0.072
r124 82 88 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.072 $X2=0.986 $Y2=0.072
r125 80 90 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.072 $X2=1.053 $Y2=0.081
r126 80 86 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.072 $X2=1.026 $Y2=0.072
r127 78 79 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.904
+ $Y=0.234 $X2=0.911 $Y2=0.234
r128 77 78 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.903
+ $Y=0.234 $X2=0.904 $Y2=0.234
r129 76 77 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.866
+ $Y=0.234 $X2=0.903 $Y2=0.234
r130 75 76 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.824
+ $Y=0.234 $X2=0.866 $Y2=0.234
r131 74 75 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.743
+ $Y=0.234 $X2=0.824 $Y2=0.234
r132 72 79 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.234 $X2=0.911 $Y2=0.234
r133 69 74 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.234 $X2=0.743 $Y2=0.234
r134 66 67 5.5679 $w=1.8e-08 $l=8.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.234 $X2=0.338 $Y2=0.234
r135 65 66 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.211
+ $Y=0.234 $X2=0.256 $Y2=0.234
r136 64 65 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.174
+ $Y=0.234 $X2=0.211 $Y2=0.234
r137 62 69 22 $w=1.8e-08 $l=3.24e-07 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.702 $Y2=0.234
r138 62 67 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.338 $Y2=0.234
r139 59 64 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.174 $Y2=0.234
r140 57 59 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.162 $Y2=0.234
r141 56 91 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.234 $X2=1.053 $Y2=0.225
r142 56 72 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.234 $X2=0.918 $Y2=0.234
r143 52 53 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.072 $X2=0.128 $Y2=0.072
r144 50 53 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.072 $X2=0.128 $Y2=0.072
r145 47 52 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.072 $X2=0.094 $Y2=0.072
r146 45 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.072 $X2=0.054 $Y2=0.072
r147 43 44 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.106 $X2=0.027 $Y2=0.207
r148 42 57 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.225 $X2=0.036 $Y2=0.234
r149 42 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.207
r150 41 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.081 $X2=0.036 $Y2=0.072
r151 41 43 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.081 $X2=0.027 $Y2=0.106
r152 39 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.234
+ $X2=0.918 $Y2=0.234
r153 36 39 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.2025 $X2=0.916 $Y2=0.2025
r154 35 69 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.234
+ $X2=0.702 $Y2=0.234
r155 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2025 $X2=0.702 $Y2=0.2025
r156 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2025 $X2=0.702 $Y2=0.2025
r157 30 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r158 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r159 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r160 24 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r161 21 24 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.164 $Y2=0.2025
r162 19 86 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.072
+ $X2=1.026 $Y2=0.072
r163 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.0675 $X2=1.024 $Y2=0.0675
r164 15 82 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.072
+ $X2=0.918 $Y2=0.072
r165 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.0675 $X2=0.918 $Y2=0.0675
r166 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.935 $Y=0.0675 $X2=0.918 $Y2=0.0675
r167 10 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.072
+ $X2=0.162 $Y2=0.072
r168 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r169 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r170 4 47 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.072 $X2=0.054
+ $Y2=0.072
r171 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends


* END of "./NAND3x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND3x2_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 N_Y_M0_d N_A_M0_g N_6_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_Y_M1_d N_A_M1_g N_6_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_Y_M2_d N_A_M2_g N_6_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_6_M3_d N_B_M3_g N_7_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_6_M4_d N_B_M4_g N_7_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 N_6_M5_d N_B_M5_g N_7_M5_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 VSS N_C_M6_g N_7_M6_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 VSS N_C_M7_g N_7_M7_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 VSS N_C_M8_g N_7_M8_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 VSS N_C_M9_g N_7_M9_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 VSS N_C_M10_g N_7_M10_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M11 VSS N_C_M11_g N_7_M11_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M12 N_8_M12_d N_B_M12_g N_7_M12_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M13 N_8_M13_d N_B_M13_g N_7_M13_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.027
M14 N_8_M14_d N_B_M14_g N_7_M14_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.027
M15 N_Y_M15_d N_A_M15_g N_8_M15_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.027
M16 N_Y_M16_d N_A_M16_g N_8_M16_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.027
M17 N_Y_M17_d N_A_M17_g N_8_M17_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M18 VDD N_A_M18_g N_Y_M18_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M19 N_Y_M19_d N_B_M19_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M20 VDD N_C_M20_g N_Y_M20_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M21 VDD N_C_M21_g N_Y_M21_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
M22 N_Y_M22_d N_B_M22_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M23 VDD N_A_M23_g N_Y_M23_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.162
*
* 
* .include "NAND3x2_ASAP7_75t_R.pex.sp.NAND3X2_ASAP7_75T_R.pxi"
* BEGIN of "./NAND3x2_ASAP7_75t_R.pex.sp.NAND3X2_ASAP7_75T_R.pxi"
* File: NAND3x2_ASAP7_75t_R.pex.sp.NAND3X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:40:35 2017
* 
x_PM_NAND3X2_ASAP7_75T_R%A N_A_M0_g N_A_M1_g N_A_M2_g N_A_c_4_p N_A_M18_g
+ N_A_M15_g N_A_M23_g N_A_M16_g N_A_M17_g N_A_c_9_p N_A_c_12_p N_A_c_18_p
+ N_A_c_59_p N_A_c_63_p A VSS PM_NAND3X2_ASAP7_75T_R%A
x_PM_NAND3X2_ASAP7_75T_R%B N_B_M3_g N_B_M4_g N_B_M5_g N_B_c_73_n N_B_M19_g
+ N_B_M12_g N_B_M22_g N_B_M13_g N_B_M14_g N_B_c_78_n N_B_c_80_n B N_B_c_82_n
+ N_B_c_83_n N_B_c_84_n N_B_c_85_n N_B_c_86_n N_B_c_87_n VSS
+ PM_NAND3X2_ASAP7_75T_R%B
x_PM_NAND3X2_ASAP7_75T_R%C N_C_M6_g N_C_M20_g N_C_M7_g N_C_M8_g N_C_M9_g
+ N_C_M10_g N_C_M11_g N_C_c_145_n N_C_M21_g C VSS PM_NAND3X2_ASAP7_75T_R%C
x_PM_NAND3X2_ASAP7_75T_R%6 N_6_M1_s N_6_M0_s N_6_M3_d N_6_M2_s N_6_M5_d N_6_M4_d
+ N_6_c_187_n N_6_c_197_p N_6_c_188_n N_6_c_189_n N_6_c_191_n N_6_c_193_n
+ N_6_c_194_n N_6_c_195_n N_6_c_199_p VSS PM_NAND3X2_ASAP7_75T_R%6
x_PM_NAND3X2_ASAP7_75T_R%7 N_7_M4_s N_7_M3_s N_7_c_217_n N_7_M6_s N_7_M5_s
+ N_7_c_246_n N_7_M8_s N_7_M7_s N_7_c_231_n N_7_M10_s N_7_M9_s N_7_c_233_n
+ N_7_M12_s N_7_M11_s N_7_c_251_p N_7_M14_s N_7_M13_s N_7_c_219_n N_7_c_213_n
+ N_7_c_222_n N_7_c_214_n N_7_c_236_n N_7_c_238_n N_7_c_225_n N_7_c_242_n
+ N_7_c_226_n N_7_c_227_n N_7_c_215_n VSS PM_NAND3X2_ASAP7_75T_R%7
x_PM_NAND3X2_ASAP7_75T_R%8 N_8_M13_d N_8_M12_d N_8_M15_s N_8_M14_d N_8_M17_s
+ N_8_M16_s N_8_c_273_n N_8_c_280_n N_8_c_274_n N_8_c_267_n N_8_c_268_n
+ N_8_c_269_n N_8_c_270_n VSS PM_NAND3X2_ASAP7_75T_R%8
x_PM_NAND3X2_ASAP7_75T_R%Y N_Y_M0_d N_Y_c_346_n N_Y_M2_d N_Y_M1_d N_Y_c_294_n
+ N_Y_M16_d N_Y_M15_d N_Y_c_296_n N_Y_M17_d N_Y_c_364_n N_Y_M18_s N_Y_c_297_n
+ N_Y_M20_s N_Y_M19_d N_Y_c_300_n N_Y_M22_d N_Y_M21_s N_Y_c_301_n N_Y_M23_s
+ N_Y_c_302_n N_Y_c_305_n N_Y_c_307_n N_Y_c_308_n N_Y_c_352_n N_Y_c_310_n
+ N_Y_c_312_n N_Y_c_315_n N_Y_c_317_n N_Y_c_333_n N_Y_c_334_n N_Y_c_318_n
+ N_Y_c_339_n N_Y_c_319_n N_Y_c_321_n N_Y_c_322_n N_Y_c_324_n Y VSS
+ PM_NAND3X2_ASAP7_75T_R%Y
cc_1 N_A_M1_g N_B_M3_g 2.71887e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_2 N_A_M2_g N_B_M3_g 0.00333077f $X=0.189 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_3 N_A_M2_g N_B_M4_g 2.71887e-19 $X=0.189 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_4 N_A_c_4_p N_B_c_73_n 0.00148959f $X=0.189 $Y=0.135 $X2=0.351 $Y2=0.135
cc_5 A N_B_c_73_n 0.00167219f $X=0.894 $Y=0.192 $X2=0.351 $Y2=0.135
cc_6 N_A_M15_g N_B_M13_g 2.71887e-19 $X=0.891 $Y=0.0675 $X2=0.783 $Y2=0.0675
cc_7 N_A_M15_g N_B_M14_g 0.00333077f $X=0.891 $Y=0.0675 $X2=0.837 $Y2=0.0675
cc_8 N_A_M16_g N_B_M14_g 2.71887e-19 $X=0.945 $Y=0.0675 $X2=0.837 $Y2=0.0675
cc_9 N_A_c_9_p N_B_c_78_n 0.00147123f $X=0.999 $Y=0.135 $X2=0.837 $Y2=0.135
cc_10 A N_B_c_78_n 0.00167219f $X=0.894 $Y=0.192 $X2=0.837 $Y2=0.135
cc_11 A N_B_c_80_n 6.70023e-19 $X=0.894 $Y=0.192 $X2=0.347 $Y2=0.189
cc_12 N_A_c_12_p B 7.02527e-19 $X=0.183 $Y=0.135 $X2=0.348 $Y2=0.137
cc_13 A N_B_c_82_n 0.00498306f $X=0.894 $Y=0.192 $X2=0.725 $Y2=0.198
cc_14 A N_B_c_83_n 6.61822e-19 $X=0.894 $Y=0.192 $X2=0.356 $Y2=0.198
cc_15 A N_B_c_84_n 0.00522817f $X=0.894 $Y=0.192 $X2=0.547 $Y2=0.198
cc_16 A N_B_c_85_n 4.52398e-19 $X=0.894 $Y=0.192 $X2=0.565 $Y2=0.198
cc_17 A N_B_c_86_n 6.68469e-19 $X=0.894 $Y=0.192 $X2=0.734 $Y2=0.189
cc_18 N_A_c_18_p N_B_c_87_n 7.16807e-19 $X=0.894 $Y=0.135 $X2=0.734 $Y2=0.135
cc_19 A N_C_c_145_n 0.00401629f $X=0.894 $Y=0.192 $X2=0 $Y2=0
cc_20 A C 3.78779e-19 $X=0.894 $Y=0.192 $X2=0 $Y2=0
cc_21 N_A_c_4_p N_6_M1_s 3.67193e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_22 N_A_c_4_p N_6_c_187_n 0.00203185f $X=0.189 $Y=0.135 $X2=0.351 $Y2=0.2025
cc_23 N_A_M1_g N_6_c_188_n 2.65027e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_24 N_A_M2_g N_6_c_189_n 2.58643e-19 $X=0.189 $Y=0.0675 $X2=0.729 $Y2=0.135
cc_25 N_A_c_12_p N_6_c_189_n 4.7067e-19 $X=0.183 $Y=0.135 $X2=0.729 $Y2=0.135
cc_26 A N_6_c_191_n 5.9683e-19 $X=0.894 $Y=0.192 $X2=0.729 $Y2=0.135
cc_27 A N_7_c_213_n 9.00135e-19 $X=0.894 $Y=0.192 $X2=0.837 $Y2=0.135
cc_28 A N_7_c_214_n 0.00374227f $X=0.894 $Y=0.192 $X2=0.347 $Y2=0.135
cc_29 A N_7_c_215_n 8.86139e-19 $X=0.894 $Y=0.192 $X2=0.734 $Y2=0.1765
cc_30 N_A_c_9_p N_8_M17_s 3.67193e-19 $X=0.999 $Y=0.135 $X2=0.297 $Y2=0.135
cc_31 A N_8_c_267_n 5.67277e-19 $X=0.894 $Y=0.192 $X2=0.729 $Y2=0.135
cc_32 N_A_M16_g N_8_c_268_n 2.65027e-19 $X=0.945 $Y=0.0675 $X2=0.729 $Y2=0.2025
cc_33 N_A_c_9_p N_8_c_269_n 0.00203185f $X=0.999 $Y=0.135 $X2=0.729 $Y2=0.2025
cc_34 N_A_M15_g N_8_c_270_n 3.11408e-19 $X=0.891 $Y=0.0675 $X2=0.783 $Y2=0.0675
cc_35 N_A_c_18_p N_8_c_270_n 4.90094e-19 $X=0.894 $Y=0.135 $X2=0.783 $Y2=0.0675
cc_36 N_A_c_4_p N_Y_M2_d 3.39222e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_37 N_A_c_4_p N_Y_c_294_n 7.57503e-19 $X=0.189 $Y=0.135 $X2=0.297 $Y2=0.135
cc_38 N_A_c_9_p N_Y_M16_d 3.56132e-19 $X=0.999 $Y=0.135 $X2=0.297 $Y2=0.135
cc_39 N_A_c_9_p N_Y_c_296_n 7.57503e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_40 N_A_c_4_p N_Y_c_297_n 7.57503e-19 $X=0.189 $Y=0.135 $X2=0.729 $Y2=0.135
cc_41 N_A_c_12_p N_Y_c_297_n 7.78109e-19 $X=0.183 $Y=0.135 $X2=0.729 $Y2=0.135
cc_42 A N_Y_c_297_n 2.39784e-19 $X=0.894 $Y=0.192 $X2=0.729 $Y2=0.135
cc_43 A N_Y_c_300_n 3.68996e-19 $X=0.894 $Y=0.192 $X2=0.783 $Y2=0.0675
cc_44 A N_Y_c_301_n 3.68996e-19 $X=0.894 $Y=0.192 $X2=0.837 $Y2=0.0675
cc_45 N_A_c_9_p N_Y_c_302_n 7.57503e-19 $X=0.999 $Y=0.135 $X2=0.837 $Y2=0.135
cc_46 N_A_c_18_p N_Y_c_302_n 0.00136727f $X=0.894 $Y=0.135 $X2=0.837 $Y2=0.135
cc_47 A N_Y_c_302_n 2.84578e-19 $X=0.894 $Y=0.192 $X2=0.837 $Y2=0.135
cc_48 N_A_c_4_p N_Y_c_305_n 3.56528e-19 $X=0.189 $Y=0.135 $X2=0.347 $Y2=0.135
cc_49 N_A_c_12_p N_Y_c_305_n 0.00101083f $X=0.183 $Y=0.135 $X2=0.347 $Y2=0.135
cc_50 N_A_M1_g N_Y_c_307_n 3.34178e-19 $X=0.135 $Y=0.0675 $X2=0.356 $Y2=0.198
cc_51 N_A_M0_g N_Y_c_308_n 4.944e-19 $X=0.081 $Y=0.0675 $X2=0.565 $Y2=0.198
cc_52 N_A_c_4_p N_Y_c_308_n 0.0015591f $X=0.189 $Y=0.135 $X2=0.565 $Y2=0.198
cc_53 N_A_M16_g N_Y_c_310_n 4.62055e-19 $X=0.945 $Y=0.0675 $X2=0.734 $Y2=0.135
cc_54 N_A_M17_g N_Y_c_310_n 5.55762e-19 $X=0.999 $Y=0.0675 $X2=0.734 $Y2=0.135
cc_55 N_A_M0_g N_Y_c_312_n 5.55762e-19 $X=0.081 $Y=0.0675 $X2=0.297 $Y2=0.135
cc_56 N_A_M1_g N_Y_c_312_n 4.62055e-19 $X=0.135 $Y=0.0675 $X2=0.297 $Y2=0.135
cc_57 N_A_c_4_p N_Y_c_312_n 8.58361e-19 $X=0.189 $Y=0.135 $X2=0.297 $Y2=0.135
cc_58 N_A_M2_g N_Y_c_315_n 2.63908e-19 $X=0.189 $Y=0.0675 $X2=0.347 $Y2=0.135
cc_59 N_A_c_59_p N_Y_c_315_n 0.00386156f $X=0.183 $Y=0.189 $X2=0.347 $Y2=0.135
cc_60 A N_Y_c_317_n 0.00228933f $X=0.894 $Y=0.192 $X2=0 $Y2=0
cc_61 A N_Y_c_318_n 0.00223503f $X=0.894 $Y=0.192 $X2=0 $Y2=0
cc_62 N_A_M15_g N_Y_c_319_n 2.5731e-19 $X=0.891 $Y=0.0675 $X2=0 $Y2=0
cc_63 N_A_c_63_p N_Y_c_319_n 0.00387528f $X=0.894 $Y=0.189 $X2=0 $Y2=0
cc_64 N_A_c_9_p N_Y_c_321_n 8.88792e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_65 N_A_M16_g N_Y_c_322_n 3.99019e-19 $X=0.945 $Y=0.0675 $X2=0 $Y2=0
cc_66 N_A_c_9_p N_Y_c_322_n 0.00158095f $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_67 N_A_M17_g N_Y_c_324_n 4.2024e-19 $X=0.999 $Y=0.0675 $X2=0 $Y2=0
cc_68 N_A_c_9_p Y 3.57243e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_69 N_A_c_18_p Y 9.45991e-19 $X=0.894 $Y=0.135 $X2=0 $Y2=0
cc_70 N_B_M4_g N_C_M6_g 2.71887e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_71 N_B_M5_g N_C_M6_g 0.00357042f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_72 N_B_c_84_n N_C_M6_g 4.95866e-19 $X=0.547 $Y=0.198 $X2=0.081 $Y2=0.0675
cc_73 N_B_M5_g N_C_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_74 N_B_c_84_n N_C_M7_g 4.95866e-19 $X=0.547 $Y=0.198 $X2=0.135 $Y2=0.135
cc_75 N_B_c_84_n N_C_M8_g 6.8328e-19 $X=0.547 $Y=0.198 $X2=0.189 $Y2=0.135
cc_76 N_B_c_82_n N_C_M9_g 4.01427e-19 $X=0.725 $Y=0.198 $X2=0.891 $Y2=0.0675
cc_77 N_B_M12_g N_C_M10_g 2.71887e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_78 N_B_c_82_n N_C_M10_g 4.95866e-19 $X=0.725 $Y=0.198 $X2=0 $Y2=0
cc_79 N_B_M12_g N_C_M11_g 0.00357042f $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_80 N_B_M13_g N_C_M11_g 2.71887e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_81 N_B_c_82_n N_C_M11_g 4.95866e-19 $X=0.725 $Y=0.198 $X2=0 $Y2=0
cc_82 N_B_c_73_n N_C_c_145_n 0.00150454f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_83 N_B_c_78_n N_C_c_145_n 0.00151103f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_84 B N_C_c_145_n 4.22126e-19 $X=0.348 $Y=0.137 $X2=0 $Y2=0
cc_85 N_B_c_82_n N_C_c_145_n 0.00162478f $X=0.725 $Y=0.198 $X2=0 $Y2=0
cc_86 N_B_c_84_n N_C_c_145_n 0.00196905f $X=0.547 $Y=0.198 $X2=0 $Y2=0
cc_87 B C 5.00407e-19 $X=0.348 $Y=0.137 $X2=0 $Y2=0
cc_88 N_B_c_85_n C 0.00109049f $X=0.565 $Y=0.198 $X2=0 $Y2=0
cc_89 N_B_c_87_n C 5.14428e-19 $X=0.734 $Y=0.135 $X2=0 $Y2=0
cc_90 N_B_c_73_n N_6_M5_d 3.5041e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_91 N_B_M4_g N_6_c_193_n 2.2196e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_92 N_B_c_73_n N_6_c_194_n 7.57503e-19 $X=0.351 $Y=0.135 $X2=0.945 $Y2=0.0675
cc_93 N_B_M3_g N_6_c_195_n 4.61191e-19 $X=0.243 $Y=0.0675 $X2=0.945 $Y2=0.0675
cc_94 N_B_c_73_n N_6_c_195_n 2.20764e-19 $X=0.351 $Y=0.135 $X2=0.945 $Y2=0.0675
cc_95 N_B_c_73_n N_7_M4_s 3.67575e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_96 N_B_c_73_n N_7_c_217_n 0.00203185f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_97 N_B_c_78_n N_7_M14_s 3.67575e-19 $X=0.837 $Y=0.135 $X2=0.891 $Y2=0.2025
cc_98 N_B_c_78_n N_7_c_219_n 0.00203185f $X=0.837 $Y=0.135 $X2=0.945 $Y2=0.0675
cc_99 N_B_M4_g N_7_c_213_n 4.01136e-19 $X=0.297 $Y=0.0675 $X2=0.999 $Y2=0.135
cc_100 N_B_c_73_n N_7_c_213_n 0.00106723f $X=0.351 $Y=0.135 $X2=0.999 $Y2=0.135
cc_101 N_B_M5_g N_7_c_222_n 3.02555e-19 $X=0.351 $Y=0.0675 $X2=0.999 $Y2=0.135
cc_102 B N_7_c_222_n 0.00123688f $X=0.348 $Y=0.137 $X2=0.999 $Y2=0.135
cc_103 N_B_c_84_n N_7_c_214_n 9.87157e-19 $X=0.547 $Y=0.198 $X2=0.183 $Y2=0.135
cc_104 N_B_c_82_n N_7_c_225_n 9.87157e-19 $X=0.725 $Y=0.198 $X2=0.183 $Y2=0.189
cc_105 N_B_M13_g N_7_c_226_n 3.10881e-19 $X=0.783 $Y=0.0675 $X2=0.894 $Y2=0.189
cc_106 N_B_M12_g N_7_c_227_n 2.82384e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_107 N_B_c_87_n N_7_c_227_n 0.0012042f $X=0.734 $Y=0.135 $X2=0 $Y2=0
cc_108 N_B_c_78_n N_7_c_215_n 0.00105285f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_109 N_B_c_78_n N_8_M13_d 3.44816e-19 $X=0.837 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_110 N_B_c_78_n N_8_c_273_n 7.57503e-19 $X=0.837 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_111 N_B_M13_g N_8_c_274_n 2.65027e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_112 N_B_M14_g N_8_c_267_n 3.92012e-19 $X=0.837 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_113 N_B_c_78_n N_8_c_267_n 2.20618e-19 $X=0.837 $Y=0.135 $X2=0.891 $Y2=0.135
cc_114 B N_Y_c_300_n 5.80749e-19 $X=0.348 $Y=0.137 $X2=0.945 $Y2=0.0675
cc_115 N_B_c_84_n N_Y_c_300_n 0.00186448f $X=0.547 $Y=0.198 $X2=0.945 $Y2=0.0675
cc_116 N_B_c_82_n N_Y_c_301_n 0.00218056f $X=0.725 $Y=0.198 $X2=0.999 $Y2=0.0675
cc_117 N_B_c_87_n N_Y_c_301_n 5.72789e-19 $X=0.734 $Y=0.135 $X2=0.999 $Y2=0.0675
cc_118 N_B_M3_g N_Y_c_317_n 4.58673e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_119 N_B_c_73_n N_Y_c_317_n 6.40192e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_120 N_B_M4_g N_Y_c_333_n 4.62489e-19 $X=0.297 $Y=0.0675 $X2=0.945 $Y2=0.135
cc_121 N_B_M5_g N_Y_c_334_n 2.5731e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_122 N_B_M12_g N_Y_c_334_n 2.63908e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_123 N_B_c_83_n N_Y_c_334_n 0.0328889f $X=0.356 $Y=0.198 $X2=0 $Y2=0
cc_124 N_B_M13_g N_Y_c_318_n 4.62489e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_125 N_B_c_78_n N_Y_c_318_n 6.30157e-19 $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_126 N_B_M14_g N_Y_c_339_n 4.58673e-19 $X=0.837 $Y=0.0675 $X2=0 $Y2=0
cc_127 N_C_c_145_n N_7_M8_s 3.67193e-19 $X=0.675 $Y=0.135 $X2=0.135 $Y2=0.135
cc_128 N_C_c_145_n N_7_c_231_n 0.00203185f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_129 N_C_c_145_n N_7_M10_s 3.67193e-19 $X=0.675 $Y=0.135 $X2=0.189 $Y2=0.135
cc_130 N_C_c_145_n N_7_c_233_n 0.00203185f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_131 N_C_M6_g N_7_c_214_n 4.98189e-19 $X=0.405 $Y=0.0675 $X2=0.183 $Y2=0.135
cc_132 N_C_c_145_n N_7_c_214_n 0.00203644f $X=0.675 $Y=0.135 $X2=0.183 $Y2=0.135
cc_133 N_C_M7_g N_7_c_236_n 3.37351e-19 $X=0.459 $Y=0.0675 $X2=0.894 $Y2=0.135
cc_134 N_C_M8_g N_7_c_236_n 4.02808e-19 $X=0.513 $Y=0.0675 $X2=0.894 $Y2=0.135
cc_135 C N_7_c_238_n 0.00115485f $X=0.555 $Y=0.137 $X2=0.894 $Y2=0.135
cc_136 N_C_M9_g N_7_c_225_n 2.3665e-19 $X=0.567 $Y=0.0675 $X2=0.183 $Y2=0.189
cc_137 N_C_M10_g N_7_c_225_n 4.02808e-19 $X=0.621 $Y=0.0675 $X2=0.183 $Y2=0.189
cc_138 N_C_c_145_n N_7_c_225_n 0.00140374f $X=0.675 $Y=0.135 $X2=0.183 $Y2=0.189
cc_139 N_C_M11_g N_7_c_242_n 4.23461e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_140 N_C_M6_g N_Y_c_334_n 2.63908e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_141 N_C_M7_g N_Y_c_334_n 2.63908e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_142 N_C_M8_g N_Y_c_334_n 3.57615e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_143 N_C_M9_g N_Y_c_334_n 3.57615e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_144 N_C_M10_g N_Y_c_334_n 2.63908e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_145 N_C_M11_g N_Y_c_334_n 2.63908e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_146 N_6_c_197_p N_7_c_217_n 0.003312f $X=0.216 $Y=0.036 $X2=0.081 $Y2=0.135
cc_147 N_6_c_194_n N_7_c_217_n 0.00352905f $X=0.324 $Y=0.036 $X2=0.081 $Y2=0.135
cc_148 N_6_c_199_p N_7_c_217_n 0.00250914f $X=0.29 $Y=0.036 $X2=0.081 $Y2=0.135
cc_149 N_6_c_193_n N_7_c_246_n 4.49606e-19 $X=0.324 $Y=0.036 $X2=0.135 $Y2=0.135
cc_150 N_6_c_194_n N_7_c_246_n 0.00317152f $X=0.324 $Y=0.036 $X2=0.135 $Y2=0.135
cc_151 N_6_c_197_p N_7_c_213_n 4.51268e-19 $X=0.216 $Y=0.036 $X2=0.999 $Y2=0.135
cc_152 N_6_c_194_n N_7_c_213_n 0.00233206f $X=0.324 $Y=0.036 $X2=0.999 $Y2=0.135
cc_153 N_6_c_199_p N_7_c_213_n 0.00704495f $X=0.29 $Y=0.036 $X2=0.999 $Y2=0.135
cc_154 N_6_c_187_n N_Y_c_346_n 0.00337028f $X=0.108 $Y=0.036 $X2=0.081 $Y2=0.135
cc_155 N_6_c_188_n N_Y_c_346_n 3.09693e-19 $X=0.176 $Y=0.036 $X2=0.081 $Y2=0.135
cc_156 N_6_c_187_n N_Y_c_294_n 0.00352892f $X=0.108 $Y=0.036 $X2=0.135 $Y2=0.135
cc_157 N_6_c_197_p N_Y_c_294_n 0.00332044f $X=0.216 $Y=0.036 $X2=0.135 $Y2=0.135
cc_158 N_6_c_188_n N_Y_c_294_n 0.00250914f $X=0.176 $Y=0.036 $X2=0.135 $Y2=0.135
cc_159 N_6_c_197_p N_Y_c_307_n 4.48103e-19 $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_160 N_6_c_187_n N_Y_c_352_n 0.00233206f $X=0.108 $Y=0.036 $X2=0.183 $Y2=0.189
cc_161 N_6_c_188_n N_Y_c_352_n 0.00702934f $X=0.176 $Y=0.036 $X2=0.183 $Y2=0.189
cc_162 N_7_c_251_p N_8_c_273_n 0.00317169f $X=0.702 $Y=0.0675 $X2=0.189
+ $Y2=0.2025
cc_163 N_7_c_219_n N_8_c_273_n 0.00352901f $X=0.81 $Y=0.0675 $X2=0.189
+ $Y2=0.2025
cc_164 N_7_c_215_n N_8_c_273_n 0.00233206f $X=0.7765 $Y=0.072 $X2=0.189
+ $Y2=0.2025
cc_165 N_7_c_219_n N_8_c_280_n 0.00328787f $X=0.81 $Y=0.0675 $X2=0.891
+ $Y2=0.0675
cc_166 N_7_c_226_n N_8_c_280_n 4.51268e-19 $X=0.81 $Y=0.072 $X2=0.891 $Y2=0.0675
cc_167 N_7_c_251_p N_8_c_274_n 4.49606e-19 $X=0.702 $Y=0.0675 $X2=0 $Y2=0
cc_168 N_7_c_219_n N_8_c_274_n 0.00250914f $X=0.81 $Y=0.0675 $X2=0 $Y2=0
cc_169 N_7_c_215_n N_8_c_274_n 0.00697856f $X=0.7765 $Y=0.072 $X2=0 $Y2=0
cc_170 N_7_c_246_n N_Y_c_300_n 0.00158656f $X=0.378 $Y=0.0675 $X2=0.945
+ $Y2=0.0675
cc_171 N_7_c_251_p N_Y_c_301_n 0.0015999f $X=0.702 $Y=0.0675 $X2=0.999
+ $Y2=0.0675
cc_172 N_7_c_213_n N_Y_c_307_n 3.18557e-19 $X=0.338 $Y=0.072 $X2=0 $Y2=0
cc_173 N_7_c_213_n N_Y_c_333_n 4.01913e-19 $X=0.338 $Y=0.072 $X2=0.945 $Y2=0.135
cc_174 N_7_c_214_n N_Y_c_334_n 4.01913e-19 $X=0.418 $Y=0.072 $X2=0 $Y2=0
cc_175 N_7_c_215_n N_Y_c_318_n 4.01913e-19 $X=0.7765 $Y=0.072 $X2=0 $Y2=0
cc_176 N_7_c_226_n N_Y_c_322_n 3.18557e-19 $X=0.81 $Y=0.072 $X2=0 $Y2=0
cc_177 N_8_c_280_n N_Y_c_296_n 0.00328789f $X=0.864 $Y=0.036 $X2=0 $Y2=0
cc_178 N_8_c_268_n N_Y_c_296_n 0.00249187f $X=0.972 $Y=0.036 $X2=0 $Y2=0
cc_179 N_8_c_269_n N_Y_c_296_n 0.00350515f $X=0.972 $Y=0.036 $X2=0 $Y2=0
cc_180 N_8_c_268_n N_Y_c_364_n 3.09693e-19 $X=0.972 $Y=0.036 $X2=0.189
+ $Y2=0.2025
cc_181 N_8_c_269_n N_Y_c_364_n 0.00337028f $X=0.972 $Y=0.036 $X2=0.189
+ $Y2=0.2025
cc_182 N_8_c_280_n N_Y_c_322_n 4.48103e-19 $X=0.864 $Y=0.036 $X2=0 $Y2=0
cc_183 N_8_c_268_n N_Y_c_322_n 0.00704501f $X=0.972 $Y=0.036 $X2=0 $Y2=0
cc_184 N_8_c_269_n N_Y_c_322_n 0.00233206f $X=0.972 $Y=0.036 $X2=0 $Y2=0

* END of "./NAND3x2_ASAP7_75t_R.pex.sp.NAND3X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND3xp33_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:40:57 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND3xp33_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND3xp33_ASAP7_75t_R.pex.sp.pex"
* File: NAND3xp33_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:40:57 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND3XP33_ASAP7_75T_R%A 2 5 7 13 VSS
c9 13 VSS 0.00149021f $X=0.083 $Y=0.137
c10 5 VSS 0.0016745f $X=0.081 $Y=0.135
c11 2 VSS 0.0649376f $X=0.081 $Y=0.0675
r12 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r13 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NAND3XP33_ASAP7_75T_R%B 2 5 7 15 VSS
c13 15 VSS 0.00570149f $X=0.136 $Y=0.137
c14 5 VSS 0.00116826f $X=0.135 $Y=0.135
c15 2 VSS 0.0601197f $X=0.135 $Y=0.0675
r16 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_NAND3XP33_ASAP7_75T_R%C 2 7 12 13 VSS
c5 13 VSS 0.0145064f $X=0.202 $Y=0.137
c6 12 VSS 0.00522154f $X=0.2 $Y=0.135
c7 2 VSS 0.0639038f $X=0.189 $Y=0.0675
r8 12 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.2 $Y=0.135 $X2=0.2
+ $Y2=0.135
r9 5 12 11 $w=2e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.189 $Y=0.135
+ $X2=0.2 $Y2=0.135
r10 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r11 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_NAND3XP33_ASAP7_75T_R%Y 1 6 9 11 12 15 19 20 21 33 35 42 43 VSS
c12 45 VSS 9.40634e-19 $X=0.045 $Y=0.036
c13 44 VSS 0.0032947f $X=0.036 $Y=0.036
c14 43 VSS 0.00224295f $X=0.054 $Y=0.036
c15 42 VSS 0.00287833f $X=0.054 $Y=0.036
c16 36 VSS 0.00103857f $X=0.153 $Y=0.234
c17 35 VSS 0.00142296f $X=0.144 $Y=0.234
c18 34 VSS 0.00632432f $X=0.126 $Y=0.234
c19 33 VSS 0.00142296f $X=0.09 $Y=0.234
c20 32 VSS 4.19006e-19 $X=0.072 $Y=0.234
c21 31 VSS 0.00321919f $X=0.068 $Y=0.234
c22 29 VSS 0.00358469f $X=0.162 $Y=0.234
c23 24 VSS 0.00335462f $X=0.036 $Y=0.234
c24 23 VSS 4.139e-19 $X=0.027 $Y=0.2125
c25 21 VSS 0.00151641f $X=0.027 $Y=0.1065
c26 20 VSS 8.44496e-19 $X=0.027 $Y=0.07
c27 19 VSS 0.00422697f $X=0.028 $Y=0.143
c28 17 VSS 3.97344e-19 $X=0.027 $Y=0.225
c29 15 VSS 0.0075021f $X=0.162 $Y=0.216
c30 11 VSS 5.65078e-19 $X=0.179 $Y=0.216
c31 9 VSS 0.00549622f $X=0.056 $Y=0.216
c32 6 VSS 2.53241e-19 $X=0.071 $Y=0.216
c33 1 VSS 3.02808e-19 $X=0.071 $Y=0.0675
r34 44 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.045 $Y2=0.036
r35 42 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.045 $Y2=0.036
r36 42 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r37 39 44 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.036 $Y2=0.036
r38 35 36 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.153 $Y2=0.234
r39 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r40 33 34 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.126 $Y2=0.234
r41 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r42 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.068
+ $Y=0.234 $X2=0.072 $Y2=0.234
r43 29 36 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.153 $Y2=0.234
r44 26 31 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.068 $Y2=0.234
r45 24 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.054 $Y2=0.234
r46 22 23 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.2 $X2=0.027 $Y2=0.2125
r47 20 21 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.1065
r48 19 22 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.143 $X2=0.027 $Y2=0.2
r49 19 21 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.143 $X2=0.027 $Y2=0.1065
r50 17 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.225 $X2=0.036 $Y2=0.234
r51 17 23 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.2125
r52 16 39 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.036
r53 16 20 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r54 15 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r55 12 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.162 $Y2=0.216
r56 11 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.216 $X2=0.162 $Y2=0.216
r57 9 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r58 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.216 $X2=0.056 $Y2=0.216
r59 4 43 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r60 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends

.subckt PM_NAND3XP33_ASAP7_75T_R%7 1 2 VSS
c0 1 VSS 0.00221026f $X=0.125 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends

.subckt PM_NAND3XP33_ASAP7_75T_R%8 1 2 VSS
c1 1 VSS 0.00199907f $X=0.179 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.145 $Y2=0.0675
.ends


* END of "./NAND3xp33_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND3xp33_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 N_7_M0_d N_A_M0_g N_Y_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_8_M1_d N_B_M1_g N_7_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_C_M2_g N_8_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 VDD N_A_M3_g N_Y_M3_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M4 N_Y_M4_d N_B_M4_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
M5 VDD N_C_M5_g N_Y_M5_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.189
*
* 
* .include "NAND3xp33_ASAP7_75t_R.pex.sp.NAND3XP33_ASAP7_75T_R.pxi"
* BEGIN of "./NAND3xp33_ASAP7_75t_R.pex.sp.NAND3XP33_ASAP7_75T_R.pxi"
* File: NAND3xp33_ASAP7_75t_R.pex.sp.NAND3XP33_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:40:57 2017
* 
x_PM_NAND3XP33_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M3_g A VSS
+ PM_NAND3XP33_ASAP7_75T_R%A
x_PM_NAND3XP33_ASAP7_75T_R%B N_B_M1_g N_B_c_11_n N_B_M4_g B VSS
+ PM_NAND3XP33_ASAP7_75T_R%B
x_PM_NAND3XP33_ASAP7_75T_R%C N_C_M2_g N_C_M5_g N_C_c_25_n C VSS
+ PM_NAND3XP33_ASAP7_75T_R%C
x_PM_NAND3XP33_ASAP7_75T_R%Y N_Y_M0_s N_Y_M3_s N_Y_c_28_n N_Y_M5_s N_Y_M4_d
+ N_Y_c_33_n Y N_Y_c_34_n N_Y_c_29_n N_Y_c_30_n N_Y_c_35_n N_Y_c_37_n N_Y_c_32_n
+ VSS PM_NAND3XP33_ASAP7_75T_R%Y
x_PM_NAND3XP33_ASAP7_75T_R%7 N_7_M1_s N_7_M0_d VSS PM_NAND3XP33_ASAP7_75T_R%7
x_PM_NAND3XP33_ASAP7_75T_R%8 N_8_M2_s N_8_M1_d VSS PM_NAND3XP33_ASAP7_75T_R%8
cc_1 N_A_M0_g N_B_M1_g 0.00327995f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_11_n 8.52536e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A B 0.00618453f $X=0.083 $Y=0.137 $X2=0.136 $Y2=0.137
cc_4 N_A_M0_g N_C_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 A N_Y_c_28_n 3.31541e-19 $X=0.083 $Y=0.137 $X2=0 $Y2=0
cc_6 A N_Y_c_29_n 0.00548081f $X=0.083 $Y=0.137 $X2=0 $Y2=0
cc_7 N_A_M0_g N_Y_c_30_n 2.57255e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_8 A N_Y_c_30_n 0.00123619f $X=0.083 $Y=0.137 $X2=0 $Y2=0
cc_9 A N_Y_c_32_n 0.0013295f $X=0.083 $Y=0.137 $X2=0 $Y2=0
cc_10 N_B_M1_g N_C_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_11 N_B_c_11_n N_C_c_25_n 9.17588e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_12 B C 0.00690454f $X=0.136 $Y=0.137 $X2=0.083 $Y2=0.137
cc_13 B N_Y_c_33_n 3.55402e-19 $X=0.136 $Y=0.137 $X2=0 $Y2=0
cc_14 B N_Y_c_34_n 2.64182e-19 $X=0.136 $Y=0.137 $X2=0 $Y2=0
cc_15 N_B_M1_g N_Y_c_35_n 2.57255e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_16 B N_Y_c_35_n 0.00123985f $X=0.136 $Y=0.137 $X2=0 $Y2=0
cc_17 B N_Y_c_37_n 7.1001e-19 $X=0.136 $Y=0.137 $X2=0 $Y2=0
cc_18 B N_Y_c_32_n 6.83303e-19 $X=0.136 $Y=0.137 $X2=0 $Y2=0
cc_19 B N_8_M2_s 3.84149e-19 $X=0.136 $Y=0.137 $X2=0.081 $Y2=0.0675
cc_20 C N_Y_c_33_n 2.68871e-19 $X=0.202 $Y=0.137 $X2=0 $Y2=0

* END of "./NAND3xp33_ASAP7_75t_R.pex.sp.NAND3XP33_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND4xp25_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:41:20 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND4xp25_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND4xp25_ASAP7_75t_R.pex.sp.pex"
* File: NAND4xp25_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:41:20 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND4XP25_ASAP7_75T_R%D 2 5 7 19 VSS
c8 19 VSS 0.022219f $X=0.081 $Y=0.138
c9 5 VSS 0.00296916f $X=0.081 $Y=0.135
c10 2 VSS 0.0646435f $X=0.081 $Y=0.0675
r11 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r12 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r13 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NAND4XP25_ASAP7_75T_R%C 2 5 7 15 VSS
c10 15 VSS 0.00301634f $X=0.135 $Y=0.138
c11 5 VSS 0.00183837f $X=0.135 $Y=0.135
c12 2 VSS 0.0597098f $X=0.135 $Y=0.0675
r13 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_NAND4XP25_ASAP7_75T_R%B 2 5 7 15 VSS
c13 15 VSS 0.00210298f $X=0.189 $Y=0.138
c14 5 VSS 0.00106871f $X=0.189 $Y=0.135
c15 2 VSS 0.0600389f $X=0.189 $Y=0.0675
r16 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_NAND4XP25_ASAP7_75T_R%A 2 5 7 13 VSS
c9 13 VSS 0.00165342f $X=0.243 $Y=0.138
c10 5 VSS 0.00225849f $X=0.243 $Y=0.135
c11 2 VSS 0.0653596f $X=0.243 $Y=0.0675
r12 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r13 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_NAND4XP25_ASAP7_75T_R%Y 1 6 9 11 12 15 16 19 29 30 32 37 39 45 46 47
+ 52 55 VSS
c18 55 VSS 0.00396347f $X=0.288 $Y=0.036
c19 54 VSS 0.00278493f $X=0.297 $Y=0.036
c20 52 VSS 0.0022441f $X=0.27 $Y=0.036
c21 49 VSS 2.31784e-19 $X=0.297 $Y=0.207
c22 47 VSS 0.00157989f $X=0.297 $Y=0.108
c23 46 VSS 0.00129359f $X=0.297 $Y=0.07
c24 45 VSS 0.00410215f $X=0.297 $Y=0.146
c25 43 VSS 5.7946e-19 $X=0.297 $Y=0.225
c26 41 VSS 6.8347e-19 $X=0.263 $Y=0.234
c27 40 VSS 3.38363e-19 $X=0.256 $Y=0.234
c28 39 VSS 0.00146362f $X=0.252 $Y=0.234
c29 38 VSS 0.00631478f $X=0.234 $Y=0.234
c30 37 VSS 0.00146362f $X=0.198 $Y=0.234
c31 36 VSS 0.00377397f $X=0.18 $Y=0.234
c32 32 VSS 0.00146362f $X=0.144 $Y=0.234
c33 31 VSS 0.00575705f $X=0.126 $Y=0.234
c34 30 VSS 0.00322775f $X=0.095 $Y=0.234
c35 29 VSS 0.0024767f $X=0.057 $Y=0.234
c36 21 VSS 0.00591782f $X=0.288 $Y=0.234
c37 19 VSS 0.00574816f $X=0.268 $Y=0.216
c38 15 VSS 0.0079209f $X=0.162 $Y=0.216
c39 11 VSS 5.3314e-19 $X=0.179 $Y=0.216
c40 9 VSS 0.0058471f $X=0.056 $Y=0.216
c41 6 VSS 4.86827e-19 $X=0.071 $Y=0.216
c42 4 VSS 3.74006e-19 $X=0.268 $Y=0.0675
r43 55 56 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.2925 $Y2=0.036
r44 54 56 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.036 $X2=0.2925 $Y2=0.036
r45 51 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.288 $Y2=0.036
r46 51 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r47 48 49 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.2 $X2=0.297 $Y2=0.207
r48 46 47 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.07 $X2=0.297 $Y2=0.108
r49 45 48 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.146 $X2=0.297 $Y2=0.2
r50 45 47 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.146 $X2=0.297 $Y2=0.108
r51 43 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.207
r52 42 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.036
r53 42 46 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.07
r54 40 41 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.234 $X2=0.263 $Y2=0.234
r55 39 40 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.256 $Y2=0.234
r56 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r57 37 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.234 $Y2=0.234
r58 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r59 34 41 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.263 $Y2=0.234
r60 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r61 30 31 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.234 $X2=0.126 $Y2=0.234
r62 29 30 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.057
+ $Y=0.234 $X2=0.095 $Y2=0.234
r63 27 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r64 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.144 $Y2=0.234
r65 23 29 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.057 $Y2=0.234
r66 21 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.234 $X2=0.297 $Y2=0.225
r67 21 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.27 $Y2=0.234
r68 19 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r69 16 19 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.216 $X2=0.268 $Y2=0.216
r70 15 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r71 12 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.162 $Y2=0.216
r72 11 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.216 $X2=0.162 $Y2=0.216
r73 9 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r74 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.216 $X2=0.056 $Y2=0.216
r75 4 52 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r76 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.268 $Y2=0.0675
.ends

.subckt PM_NAND4XP25_ASAP7_75T_R%8 1 2 VSS
c0 1 VSS 0.00233476f $X=0.125 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends

.subckt PM_NAND4XP25_ASAP7_75T_R%9 1 2 VSS
c0 1 VSS 0.00228146f $X=0.179 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.145 $Y2=0.0675
.ends

.subckt PM_NAND4XP25_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00228146f $X=0.233 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.199 $Y2=0.0675
.ends


* END of "./NAND4xp25_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND4xp25_ASAP7_75t_R  VSS VDD D C B A Y
* 
* Y	Y
* A	A
* B	B
* C	C
* D	D
M0 N_8_M0_d N_D_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_9_M1_d N_C_M1_g N_8_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_10_M2_d N_B_M2_g N_9_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_Y_M3_d N_A_M3_g N_10_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 VDD N_D_M4_g N_Y_M4_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M5 N_Y_M5_d N_C_M5_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
M6 VDD N_B_M6_g N_Y_M6_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.189
M7 N_Y_M7_d N_A_M7_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.189
*
* 
* .include "NAND4xp25_ASAP7_75t_R.pex.sp.NAND4XP25_ASAP7_75T_R.pxi"
* BEGIN of "./NAND4xp25_ASAP7_75t_R.pex.sp.NAND4XP25_ASAP7_75T_R.pxi"
* File: NAND4xp25_ASAP7_75t_R.pex.sp.NAND4XP25_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:41:20 2017
* 
x_PM_NAND4XP25_ASAP7_75T_R%D N_D_M0_g N_D_c_2_p N_D_M4_g D VSS
+ PM_NAND4XP25_ASAP7_75T_R%D
x_PM_NAND4XP25_ASAP7_75T_R%C N_C_M1_g N_C_c_10_n N_C_M5_g C VSS
+ PM_NAND4XP25_ASAP7_75T_R%C
x_PM_NAND4XP25_ASAP7_75T_R%B N_B_M2_g N_B_c_21_n N_B_M6_g B VSS
+ PM_NAND4XP25_ASAP7_75T_R%B
x_PM_NAND4XP25_ASAP7_75T_R%A N_A_M3_g N_A_c_34_n N_A_M7_g A VSS
+ PM_NAND4XP25_ASAP7_75T_R%A
x_PM_NAND4XP25_ASAP7_75T_R%Y N_Y_M3_d N_Y_M4_s N_Y_c_41_n N_Y_M6_s N_Y_M5_d
+ N_Y_c_45_n N_Y_M7_d N_Y_c_54_n N_Y_c_42_n N_Y_c_43_n N_Y_c_46_n N_Y_c_49_n
+ N_Y_c_55_n Y N_Y_c_51_n N_Y_c_57_n N_Y_c_52_n N_Y_c_53_n VSS
+ PM_NAND4XP25_ASAP7_75T_R%Y
x_PM_NAND4XP25_ASAP7_75T_R%8 N_8_M1_s N_8_M0_d VSS PM_NAND4XP25_ASAP7_75T_R%8
x_PM_NAND4XP25_ASAP7_75T_R%9 N_9_M2_s N_9_M1_d VSS PM_NAND4XP25_ASAP7_75T_R%9
x_PM_NAND4XP25_ASAP7_75T_R%10 N_10_M3_s N_10_M2_d VSS
+ PM_NAND4XP25_ASAP7_75T_R%10
cc_1 N_D_M0_g N_C_M1_g 0.0032073f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_D_c_2_p N_C_c_10_n 0.00101358f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 D C 0.00294306f $X=0.081 $Y=0.138 $X2=0.135 $Y2=0.138
cc_4 N_D_M0_g N_B_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 D N_Y_c_41_n 0.00214868f $X=0.081 $Y=0.138 $X2=0 $Y2=0
cc_6 D N_Y_c_42_n 0.00194715f $X=0.081 $Y=0.138 $X2=0 $Y2=0
cc_7 N_D_M0_g N_Y_c_43_n 4.31632e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_8 D N_Y_c_43_n 3.65373e-19 $X=0.081 $Y=0.138 $X2=0 $Y2=0
cc_9 N_C_M1_g N_B_M2_g 0.0035196f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_10 N_C_c_10_n N_B_c_21_n 7.51247e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_11 C B 0.00814915f $X=0.135 $Y=0.138 $X2=0.081 $Y2=0.135
cc_12 N_C_M1_g N_A_M3_g 2.71887e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_13 C N_Y_c_45_n 3.24828e-19 $X=0.135 $Y=0.138 $X2=0.081 $Y2=0.135
cc_14 N_C_M1_g N_Y_c_46_n 2.64924e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 C N_Y_c_46_n 0.00125705f $X=0.135 $Y=0.138 $X2=0 $Y2=0
cc_16 N_B_M2_g N_A_M3_g 0.00333077f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 N_B_c_21_n N_A_c_34_n 7.51046e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_18 B A 0.00620922f $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_19 B N_Y_c_45_n 3.31541e-19 $X=0.189 $Y=0.138 $X2=0.081 $Y2=0.135
cc_20 N_B_M2_g N_Y_c_49_n 2.64606e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_21 B N_Y_c_49_n 0.0012569f $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_22 B N_Y_c_51_n 2.69891e-19 $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_23 B N_Y_c_52_n 4.68998e-19 $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_24 B N_Y_c_53_n 4.44922e-19 $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_25 A N_Y_c_54_n 3.31541e-19 $X=0.243 $Y=0.138 $X2=0 $Y2=0
cc_26 N_A_M3_g N_Y_c_55_n 2.64924e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_27 A N_Y_c_55_n 0.00125383f $X=0.243 $Y=0.138 $X2=0 $Y2=0
cc_28 A N_Y_c_57_n 0.0054927f $X=0.243 $Y=0.138 $X2=0 $Y2=0
cc_29 A N_Y_c_52_n 0.0013295f $X=0.243 $Y=0.138 $X2=0 $Y2=0

* END of "./NAND4xp25_ASAP7_75t_R.pex.sp.NAND4XP25_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND4xp75_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:41:42 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND4xp75_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND4xp75_ASAP7_75t_R.pex.sp.pex"
* File: NAND4xp75_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:41:42 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND4XP75_ASAP7_75T_R%D 2 7 10 15 18 21 23 41 VSS
c16 41 VSS 0.0314045f $X=0.081 $Y=0.138
c17 21 VSS 0.0109493f $X=0.189 $Y=0.135
c18 18 VSS 0.0622597f $X=0.189 $Y=0.0675
c19 10 VSS 0.0638991f $X=0.135 $Y=0.0675
c20 2 VSS 0.0646334f $X=0.081 $Y=0.0675
r21 21 23 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r22 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r23 13 21 60 $w=1.8e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135 $Y=0.135
+ $X2=0.189 $Y2=0.135
r24 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r25 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r26 5 13 60 $w=1.8e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081 $Y=0.135
+ $X2=0.135 $Y2=0.135
r27 5 41 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r28 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r29 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NAND4XP75_ASAP7_75T_R%C 2 7 10 15 18 21 23 33 VSS
c35 33 VSS 0.00488597f $X=0.3 $Y=0.138
c36 21 VSS 0.00619913f $X=0.351 $Y=0.135
c37 18 VSS 0.0624063f $X=0.351 $Y=0.0675
c38 10 VSS 0.0636165f $X=0.297 $Y=0.0675
c39 2 VSS 0.0620301f $X=0.243 $Y=0.0675
r40 21 23 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.216
r41 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r42 13 21 60 $w=1.8e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297 $Y=0.135
+ $X2=0.351 $Y2=0.135
r43 13 33 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r44 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.216
r45 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r46 5 13 60 $w=1.8e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243 $Y=0.135
+ $X2=0.297 $Y2=0.135
r47 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r48 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_NAND4XP75_ASAP7_75T_R%B 2 7 10 15 18 21 23 29 VSS
c34 29 VSS 0.00265618f $X=0.521 $Y=0.138
c35 21 VSS 0.00647024f $X=0.513 $Y=0.135
c36 18 VSS 0.0621861f $X=0.513 $Y=0.0675
c37 10 VSS 0.0640813f $X=0.459 $Y=0.0675
c38 2 VSS 0.0623945f $X=0.405 $Y=0.0675
r39 21 29 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r40 21 23 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.216
r41 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
r42 13 21 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459 $Y=0.135
+ $X2=0.513 $Y2=0.135
r43 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.216
r44 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r45 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405 $Y=0.135
+ $X2=0.459 $Y2=0.135
r46 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.216
r47 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_NAND4XP75_ASAP7_75T_R%A 2 7 10 15 18 21 23 31 VSS
c27 31 VSS 0.00148865f $X=0.621 $Y=0.138
c28 21 VSS 0.00699989f $X=0.675 $Y=0.135
c29 18 VSS 0.066303f $X=0.675 $Y=0.0675
c30 10 VSS 0.0636276f $X=0.621 $Y=0.0675
c31 2 VSS 0.0627233f $X=0.567 $Y=0.0675
r32 21 23 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.216
r33 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0675 $X2=0.675 $Y2=0.135
r34 13 21 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621 $Y=0.135
+ $X2=0.675 $Y2=0.135
r35 13 31 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r36 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.216
r37 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
r38 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.567 $Y=0.135
+ $X2=0.621 $Y2=0.135
r39 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.216
r40 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
.ends

.subckt PM_NAND4XP75_ASAP7_75T_R%7 1 2 6 7 11 12 17 18 24 25 26 28 29 31 VSS
c28 31 VSS 0.0024855f $X=0.256 $Y=0.036
c29 30 VSS 9.70579e-19 $X=0.225 $Y=0.036
c30 29 VSS 0.00283956f $X=0.324 $Y=0.036
c31 28 VSS 0.00708487f $X=0.324 $Y=0.036
c32 26 VSS 3.3597e-19 $X=0.2115 $Y=0.036
c33 25 VSS 0.0118841f $X=0.207 $Y=0.036
c34 24 VSS 0.00618448f $X=0.216 $Y=0.036
c35 18 VSS 0.00903596f $X=0.108 $Y=0.036
c36 17 VSS 0.00160315f $X=0.108 $Y=0.036
c37 11 VSS 6.1922e-19 $X=0.341 $Y=0.0675
c38 6 VSS 6.20841e-19 $X=0.233 $Y=0.0675
c39 1 VSS 5.24403e-19 $X=0.125 $Y=0.0675
r40 30 31 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.036 $X2=0.256 $Y2=0.036
r41 28 31 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.256 $Y2=0.036
r42 28 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r43 25 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.036 $X2=0.2115 $Y2=0.036
r44 23 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.225 $Y2=0.036
r45 23 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.2115 $Y2=0.036
r46 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r47 17 25 6.72222 $w=1.8e-08 $l=9.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.207 $Y2=0.036
r48 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r49 15 29 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r50 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r51 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r52 10 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r53 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r54 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r55 5 18 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r56 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r57 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends

.subckt PM_NAND4XP75_ASAP7_75T_R%8 1 2 5 6 7 10 11 12 15 23 24 26 28 29 VSS
c31 29 VSS 3.56711e-19 $X=0.4485 $Y=0.072
c32 28 VSS 0.00305582f $X=0.412 $Y=0.072
c33 26 VSS 4.07927e-19 $X=0.485 $Y=0.072
c34 24 VSS 3.19402e-19 $X=0.34 $Y=0.072
c35 23 VSS 8.46035e-21 $X=0.306 $Y=0.072
c36 15 VSS 0.00387497f $X=0.486 $Y=0.0675
c37 11 VSS 5.71502e-19 $X=0.503 $Y=0.0675
c38 10 VSS 0.00180298f $X=0.378 $Y=0.0675
c39 6 VSS 7.40637e-19 $X=0.395 $Y=0.0675
c40 5 VSS 0.00353193f $X=0.27 $Y=0.0675
c41 1 VSS 6.21322e-19 $X=0.287 $Y=0.0675
r42 28 29 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.412
+ $Y=0.072 $X2=0.4485 $Y2=0.072
r43 26 29 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.485
+ $Y=0.072 $X2=0.4485 $Y2=0.072
r44 23 24 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.072 $X2=0.34 $Y2=0.072
r45 21 28 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.412 $Y2=0.072
r46 21 24 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.34 $Y2=0.072
r47 17 23 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.072 $X2=0.306 $Y2=0.072
r48 15 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.485 $Y=0.072 $X2=0.485
+ $Y2=0.072
r49 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.486 $Y2=0.0675
r50 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.0675 $X2=0.486 $Y2=0.0675
r51 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.072 $X2=0.378
+ $Y2=0.072
r52 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.378 $Y2=0.0675
r53 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.0675 $X2=0.378 $Y2=0.0675
r54 5 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.072 $X2=0.27
+ $Y2=0.072
r55 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
r56 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends

.subckt PM_NAND4XP75_ASAP7_75T_R%9 1 2 6 7 11 12 18 22 23 25 26 28 29 31 VSS
c33 31 VSS 0.00288066f $X=0.58 $Y=0.036
c34 30 VSS 9.70579e-19 $X=0.549 $Y=0.036
c35 29 VSS 0.00276854f $X=0.648 $Y=0.036
c36 28 VSS 0.00738141f $X=0.648 $Y=0.036
c37 26 VSS 3.3597e-19 $X=0.5355 $Y=0.036
c38 25 VSS 0.00212432f $X=0.531 $Y=0.036
c39 24 VSS 6.07508e-19 $X=0.504 $Y=0.036
c40 23 VSS 0.00739746f $X=0.499 $Y=0.036
c41 22 VSS 0.00216821f $X=0.54 $Y=0.036
c42 18 VSS 0.00283848f $X=0.432 $Y=0.036
c43 11 VSS 6.30433e-19 $X=0.665 $Y=0.0675
c44 6 VSS 6.20841e-19 $X=0.557 $Y=0.0675
c45 1 VSS 6.25349e-19 $X=0.449 $Y=0.0675
r46 30 31 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.549
+ $Y=0.036 $X2=0.58 $Y2=0.036
r47 28 31 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.58 $Y2=0.036
r48 28 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036 $X2=0.648
+ $Y2=0.036
r49 25 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.531
+ $Y=0.036 $X2=0.5355 $Y2=0.036
r50 24 25 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.531 $Y2=0.036
r51 23 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.499
+ $Y=0.036 $X2=0.504 $Y2=0.036
r52 21 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.549 $Y2=0.036
r53 21 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.5355 $Y2=0.036
r54 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r55 17 23 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.499 $Y2=0.036
r56 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r57 15 29 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.648
+ $Y=0.0675 $X2=0.648 $Y2=0.036
r58 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.648 $Y2=0.0675
r59 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0675 $X2=0.648 $Y2=0.0675
r60 10 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r61 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r62 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r63 5 18 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r64 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.432 $Y2=0.0675
r65 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.449
+ $Y=0.0675 $X2=0.432 $Y2=0.0675
.ends

.subckt PM_NAND4XP75_ASAP7_75T_R%Y 1 2 5 6 9 11 12 15 16 17 20 21 22 25 26 27 30
+ 31 32 35 36 37 40 41 43 51 52 56 57 64 66 67 72 74 83 84 85 86 90 92 VSS
c58 94 VSS 7.14098e-19 $X=0.729 $Y=0.2125
c59 92 VSS 0.00110969f $X=0.729 $Y=0.126
c60 91 VSS 0.00116545f $X=0.729 $Y=0.106
c61 90 VSS 0.00379407f $X=0.732 $Y=0.146
c62 88 VSS 6.07272e-19 $X=0.729 $Y=0.225
c63 86 VSS 6.39993e-19 $X=0.6845 $Y=0.072
c64 85 VSS 3.43772e-19 $X=0.666 $Y=0.072
c65 84 VSS 8.46035e-21 $X=0.63 $Y=0.072
c66 83 VSS 3.77963e-19 $X=0.612 $Y=0.072
c67 75 VSS 0.00367873f $X=0.72 $Y=0.072
c68 74 VSS 0.00146362f $X=0.63 $Y=0.234
c69 73 VSS 0.00501797f $X=0.612 $Y=0.234
c70 72 VSS 0.00285554f $X=0.58 $Y=0.234
c71 71 VSS 0.00172044f $X=0.549 $Y=0.234
c72 67 VSS 8.32314e-19 $X=0.531 $Y=0.234
c73 66 VSS 0.00142296f $X=0.522 $Y=0.234
c74 65 VSS 5.34627e-19 $X=0.504 $Y=0.234
c75 64 VSS 0.0214141f $X=0.499 $Y=0.234
c76 57 VSS 0.00146362f $X=0.306 $Y=0.234
c77 56 VSS 0.00900134f $X=0.288 $Y=0.234
c78 52 VSS 4.42399e-19 $X=0.2115 $Y=0.234
c79 51 VSS 0.0117964f $X=0.207 $Y=0.234
c80 43 VSS 0.00128823f $X=0.108 $Y=0.234
c81 41 VSS 0.0134649f $X=0.72 $Y=0.234
c82 40 VSS 0.00824104f $X=0.648 $Y=0.216
c83 36 VSS 5.3314e-19 $X=0.665 $Y=0.216
c84 35 VSS 0.00775062f $X=0.54 $Y=0.216
c85 31 VSS 5.3314e-19 $X=0.557 $Y=0.216
c86 30 VSS 0.00774743f $X=0.432 $Y=0.216
c87 26 VSS 5.3314e-19 $X=0.449 $Y=0.216
c88 25 VSS 0.00820645f $X=0.324 $Y=0.216
c89 21 VSS 5.3314e-19 $X=0.341 $Y=0.216
c90 20 VSS 0.0073284f $X=0.216 $Y=0.216
c91 16 VSS 5.3314e-19 $X=0.233 $Y=0.216
c92 15 VSS 0.00750643f $X=0.108 $Y=0.216
c93 11 VSS 5.5175e-19 $X=0.125 $Y=0.216
c94 9 VSS 0.00220041f $X=0.7 $Y=0.0675
c95 5 VSS 0.00395433f $X=0.594 $Y=0.0675
c96 1 VSS 5.7545e-19 $X=0.611 $Y=0.0675
r97 93 94 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.2 $X2=0.729 $Y2=0.2125
r98 91 92 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.106 $X2=0.729 $Y2=0.126
r99 90 93 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.146 $X2=0.729 $Y2=0.2
r100 90 92 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.146 $X2=0.729 $Y2=0.126
r101 88 94 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.225 $X2=0.729 $Y2=0.2125
r102 87 91 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.081 $X2=0.729 $Y2=0.106
r103 85 86 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.072 $X2=0.6845 $Y2=0.072
r104 84 85 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.072 $X2=0.666 $Y2=0.072
r105 83 84 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.072 $X2=0.63 $Y2=0.072
r106 81 86 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.703
+ $Y=0.072 $X2=0.6845 $Y2=0.072
r107 77 83 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.072 $X2=0.612 $Y2=0.072
r108 75 87 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.072 $X2=0.729 $Y2=0.081
r109 75 81 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.072 $X2=0.703 $Y2=0.072
r110 73 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.63 $Y2=0.234
r111 72 73 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.58
+ $Y=0.234 $X2=0.612 $Y2=0.234
r112 71 72 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.549
+ $Y=0.234 $X2=0.58 $Y2=0.234
r113 69 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.63 $Y2=0.234
r114 66 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.234 $X2=0.531 $Y2=0.234
r115 65 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.522 $Y2=0.234
r116 64 65 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.499
+ $Y=0.234 $X2=0.504 $Y2=0.234
r117 62 71 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.549 $Y2=0.234
r118 62 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.531 $Y2=0.234
r119 59 64 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.499 $Y2=0.234
r120 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.306 $Y2=0.234
r121 54 59 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r122 54 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.306 $Y2=0.234
r123 51 52 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.234 $X2=0.2115 $Y2=0.234
r124 49 56 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.288 $Y2=0.234
r125 49 52 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.2115 $Y2=0.234
r126 43 51 6.72222 $w=1.8e-08 $l=9.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.207 $Y2=0.234
r127 41 88 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.234 $X2=0.729 $Y2=0.225
r128 41 69 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.234 $X2=0.648 $Y2=0.234
r129 40 69 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234
+ $X2=0.648 $Y2=0.234
r130 37 40 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.216 $X2=0.648 $Y2=0.216
r131 36 40 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.216 $X2=0.648 $Y2=0.216
r132 35 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r133 32 35 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.216 $X2=0.54 $Y2=0.216
r134 31 35 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.216 $X2=0.54 $Y2=0.216
r135 30 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r136 27 30 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.216 $X2=0.432 $Y2=0.216
r137 26 30 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.216 $X2=0.432 $Y2=0.216
r138 25 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r139 22 25 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.216 $X2=0.324 $Y2=0.216
r140 21 25 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.216 $X2=0.324 $Y2=0.216
r141 20 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r142 17 20 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.216 $X2=0.216 $Y2=0.216
r143 16 20 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.216 $X2=0.216 $Y2=0.216
r144 15 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r145 12 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.216 $X2=0.108 $Y2=0.216
r146 11 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.216 $X2=0.108 $Y2=0.216
r147 9 81 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.703 $Y=0.072 $X2=0.703
+ $Y2=0.072
r148 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.0675 $X2=0.7 $Y2=0.0675
r149 5 77 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.072 $X2=0.594
+ $Y2=0.072
r150 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0675 $X2=0.594 $Y2=0.0675
r151 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.0675 $X2=0.594 $Y2=0.0675
.ends


* END of "./NAND4xp75_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND4xp75_ASAP7_75t_R  VSS VDD D C B A Y
* 
* Y	Y
* A	A
* B	B
* C	C
* D	D
M0 N_7_M0_d N_D_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_7_M1_d N_D_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_7_M2_d N_D_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_8_M3_d N_C_M3_g N_7_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_8_M4_d N_C_M4_g N_7_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 N_8_M5_d N_C_M5_g N_7_M5_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 N_9_M6_d N_B_M6_g N_8_M6_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_9_M7_d N_B_M7_g N_8_M7_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_9_M8_d N_B_M8_g N_8_M8_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 N_Y_M9_d N_A_M9_g N_9_M9_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M10 N_Y_M10_d N_A_M10_g N_9_M10_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M11 N_Y_M11_d N_A_M11_g N_9_M11_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M12 N_Y_M12_d N_D_M12_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M13 N_Y_M13_d N_D_M13_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M14 N_Y_M14_d N_D_M14_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M15 VDD N_C_M15_g N_Y_M15_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M16 VDD N_C_M16_g N_Y_M16_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.189
M17 VDD N_C_M17_g N_Y_M17_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341
+ $Y=0.189
M18 N_Y_M18_d N_B_M18_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.395
+ $Y=0.189
M19 N_Y_M19_d N_B_M19_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.449
+ $Y=0.189
M20 N_Y_M20_d N_B_M20_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.503
+ $Y=0.189
M21 VDD N_A_M21_g N_Y_M21_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.557
+ $Y=0.189
M22 VDD N_A_M22_g N_Y_M22_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.611
+ $Y=0.189
M23 VDD N_A_M23_g N_Y_M23_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.665
+ $Y=0.189
*
* 
* .include "NAND4xp75_ASAP7_75t_R.pex.sp.NAND4XP75_ASAP7_75T_R.pxi"
* BEGIN of "./NAND4xp75_ASAP7_75t_R.pex.sp.NAND4XP75_ASAP7_75T_R.pxi"
* File: NAND4xp75_ASAP7_75t_R.pex.sp.NAND4XP75_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:41:42 2017
* 
x_PM_NAND4XP75_ASAP7_75T_R%D N_D_M0_g N_D_M12_g N_D_M1_g N_D_M13_g N_D_M2_g
+ N_D_c_4_p N_D_M14_g D VSS PM_NAND4XP75_ASAP7_75T_R%D
x_PM_NAND4XP75_ASAP7_75T_R%C N_C_M3_g N_C_M15_g N_C_M4_g N_C_M16_g N_C_M5_g
+ N_C_c_20_n N_C_M17_g C VSS PM_NAND4XP75_ASAP7_75T_R%C
x_PM_NAND4XP75_ASAP7_75T_R%B N_B_M6_g N_B_M18_g N_B_M7_g N_B_M19_g N_B_M8_g
+ N_B_c_55_n N_B_M20_g B VSS PM_NAND4XP75_ASAP7_75T_R%B
x_PM_NAND4XP75_ASAP7_75T_R%A N_A_M9_g N_A_M21_g N_A_M10_g N_A_M22_g N_A_M11_g
+ N_A_c_89_n N_A_M23_g A VSS PM_NAND4XP75_ASAP7_75T_R%A
x_PM_NAND4XP75_ASAP7_75T_R%7 N_7_M1_d N_7_M0_d N_7_M3_s N_7_M2_d N_7_M5_s
+ N_7_M4_s N_7_c_114_n N_7_c_116_n N_7_c_120_n N_7_c_117_n N_7_c_121_n
+ N_7_c_122_n N_7_c_123_n N_7_c_125_n VSS PM_NAND4XP75_ASAP7_75T_R%7
x_PM_NAND4XP75_ASAP7_75T_R%8 N_8_M4_d N_8_M3_d N_8_c_142_n N_8_M6_s N_8_M5_d
+ N_8_c_158_n N_8_M8_s N_8_M7_s N_8_c_149_n N_8_c_144_n N_8_c_146_n N_8_c_151_n
+ N_8_c_147_n N_8_c_165_p VSS PM_NAND4XP75_ASAP7_75T_R%8
x_PM_NAND4XP75_ASAP7_75T_R%9 N_9_M7_d N_9_M6_d N_9_M9_s N_9_M8_d N_9_M11_s
+ N_9_M10_s N_9_c_173_n N_9_c_174_n N_9_c_175_n N_9_c_177_n N_9_c_179_n
+ N_9_c_181_n N_9_c_182_n N_9_c_183_n VSS PM_NAND4XP75_ASAP7_75T_R%9
x_PM_NAND4XP75_ASAP7_75T_R%Y N_Y_M10_d N_Y_M9_d N_Y_c_230_n N_Y_M11_d
+ N_Y_c_255_n N_Y_M13_d N_Y_M12_d N_Y_c_205_n N_Y_M15_s N_Y_M14_d N_Y_c_247_n
+ N_Y_M17_s N_Y_M16_s N_Y_c_210_n N_Y_M19_d N_Y_M18_d N_Y_c_220_n N_Y_M21_s
+ N_Y_M20_d N_Y_c_221_n N_Y_M23_s N_Y_M22_s N_Y_c_231_n N_Y_c_233_n N_Y_c_206_n
+ N_Y_c_208_n N_Y_c_212_n N_Y_c_213_n N_Y_c_216_n N_Y_c_218_n N_Y_c_225_n
+ N_Y_c_227_n N_Y_c_235_n N_Y_c_237_n N_Y_c_228_n N_Y_c_240_n N_Y_c_242_n
+ N_Y_c_243_n Y N_Y_c_245_n VSS PM_NAND4XP75_ASAP7_75T_R%Y
cc_1 N_D_M1_g N_C_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_2 N_D_M2_g N_C_M3_g 0.00344695f $X=0.189 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_3 N_D_M2_g N_C_M4_g 2.66145e-19 $X=0.189 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_4 N_D_c_4_p N_C_c_20_n 0.00139993f $X=0.189 $Y=0.135 $X2=0.351 $Y2=0.135
cc_5 D C 2.41551e-19 $X=0.081 $Y=0.138 $X2=0.3 $Y2=0.138
cc_6 N_D_c_4_p N_7_M1_d 3.47207e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_7 N_D_c_4_p N_7_c_114_n 0.00129866f $X=0.189 $Y=0.135 $X2=0.351 $Y2=0.0675
cc_8 D N_7_c_114_n 7.8813e-19 $X=0.081 $Y=0.138 $X2=0.351 $Y2=0.0675
cc_9 N_D_c_4_p N_7_c_116_n 8.23937e-19 $X=0.189 $Y=0.135 $X2=0.351 $Y2=0.0675
cc_10 N_D_M1_g N_7_c_117_n 4.637e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_11 N_D_M2_g N_7_c_117_n 4.637e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_12 N_D_c_4_p N_Y_c_205_n 3.69297e-19 $X=0.189 $Y=0.135 $X2=0.297 $Y2=0.216
cc_13 N_D_c_4_p N_Y_c_206_n 0.00126095f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_14 D N_Y_c_206_n 7.47007e-19 $X=0.081 $Y=0.138 $X2=0 $Y2=0
cc_15 N_D_M1_g N_Y_c_208_n 4.637e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_16 N_D_M2_g N_Y_c_208_n 4.637e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_17 N_C_M4_g N_B_M6_g 2.71887e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_18 N_C_M5_g N_B_M6_g 0.00333077f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_19 N_C_M5_g N_B_M7_g 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_20 N_C_c_20_n N_B_c_55_n 0.00136412f $X=0.351 $Y=0.135 $X2=0.189 $Y2=0.135
cc_21 C B 6.03898e-19 $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_22 N_C_c_20_n N_7_M5_s 3.53818e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_23 C N_7_c_120_n 0.00300227f $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_24 C N_7_c_121_n 0.00101769f $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_25 N_C_M4_g N_7_c_122_n 2.38737e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_C_c_20_n N_7_c_123_n 8.23937e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_27 C N_7_c_123_n 2.5649e-19 $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_28 N_C_M3_g N_7_c_125_n 3.88389e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_29 C N_7_c_125_n 9.37582e-19 $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_30 N_C_c_20_n N_8_M4_d 3.46366e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_31 N_C_c_20_n N_8_c_142_n 8.23937e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_32 C N_8_c_142_n 0.00158145f $X=0.3 $Y=0.138 $X2=0.081 $Y2=0.135
cc_33 N_C_M4_g N_8_c_144_n 2.60457e-19 $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.216
cc_34 C N_8_c_144_n 0.00445699f $X=0.3 $Y=0.138 $X2=0.189 $Y2=0.216
cc_35 N_C_c_20_n N_8_c_146_n 8.71744e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_36 N_C_M5_g N_8_c_147_n 4.99916e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_C_c_20_n N_Y_c_210_n 3.69297e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_38 C N_Y_c_210_n 3.86867e-19 $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_39 C N_Y_c_212_n 5.24578e-19 $X=0.3 $Y=0.138 $X2=0.135 $Y2=0.135
cc_40 N_C_M3_g N_Y_c_213_n 4.5519e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_41 N_C_c_20_n N_Y_c_213_n 6.79963e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_42 C N_Y_c_213_n 5.24578e-19 $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_43 N_C_M4_g N_Y_c_216_n 2.64924e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_44 C N_Y_c_216_n 0.00124933f $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_45 N_C_M5_g N_Y_c_218_n 4.67322e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_46 N_C_c_20_n N_Y_c_218_n 5.37353e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_47 N_B_M7_g N_A_M9_g 2.71887e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_48 N_B_M8_g N_A_M9_g 0.00357042f $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_49 N_B_M8_g N_A_M10_g 2.71887e-19 $X=0.513 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_50 N_B_c_55_n N_A_c_89_n 0.00121234f $X=0.513 $Y=0.135 $X2=0.189 $Y2=0.135
cc_51 B A 0.00191741f $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_52 N_B_c_55_n N_8_M8_s 3.67702e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_53 N_B_c_55_n N_8_c_149_n 8.69026e-19 $X=0.513 $Y=0.135 $X2=0.135 $Y2=0.216
cc_54 B N_8_c_149_n 2.62694e-19 $X=0.521 $Y=0.138 $X2=0.135 $Y2=0.216
cc_55 N_B_M7_g N_8_c_151_n 4.0114e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_56 B N_8_c_151_n 4.95077e-19 $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_57 N_B_M6_g N_8_c_147_n 4.15837e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_B_c_55_n N_8_c_147_n 0.00156237f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_59 N_B_c_55_n N_9_M7_d 3.67193e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_60 N_B_c_55_n N_9_c_173_n 8.69026e-19 $X=0.513 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_61 B N_9_c_174_n 0.00274509f $X=0.521 $Y=0.138 $X2=0.189 $Y2=0.216
cc_62 N_B_M6_g N_9_c_175_n 2.16933e-19 $X=0.405 $Y=0.0675 $X2=0.189 $Y2=0.216
cc_63 N_B_M7_g N_9_c_175_n 2.65027e-19 $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.216
cc_64 N_B_M8_g N_9_c_177_n 3.43821e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_65 B N_9_c_177_n 8.36482e-19 $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_66 B N_9_c_179_n 0.00101769f $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_67 N_B_c_55_n N_Y_c_220_n 3.75758e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_68 B N_Y_c_221_n 3.83412e-19 $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_69 N_B_M6_g N_Y_c_218_n 4.65034e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_70 N_B_M7_g N_Y_c_218_n 4.65034e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_71 N_B_c_55_n N_Y_c_218_n 0.00126591f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_72 N_B_M8_g N_Y_c_225_n 2.57255e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_73 B N_Y_c_225_n 0.00123176f $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_74 B N_Y_c_227_n 4.04735e-19 $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_75 B N_Y_c_228_n 6.57587e-19 $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_76 N_A_c_89_n N_9_M11_s 3.67193e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_77 N_A_M10_g N_9_c_181_n 2.38524e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_78 N_A_c_89_n N_9_c_182_n 8.69026e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_79 N_A_M9_g N_9_c_183_n 4.61191e-19 $X=0.567 $Y=0.0675 $X2=0.297 $Y2=0.135
cc_80 N_A_c_89_n N_9_c_183_n 2.50471e-19 $X=0.675 $Y=0.135 $X2=0.297 $Y2=0.135
cc_81 N_A_c_89_n N_Y_M10_d 3.67575e-19 $X=0.675 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_82 N_A_c_89_n N_Y_c_230_n 8.69026e-19 $X=0.675 $Y=0.135 $X2=0.243 $Y2=0.135
cc_83 N_A_c_89_n N_Y_c_231_n 3.75758e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_84 A N_Y_c_231_n 3.83412e-19 $X=0.621 $Y=0.138 $X2=0 $Y2=0
cc_85 N_A_M11_g N_Y_c_233_n 4.38953e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_86 N_A_c_89_n N_Y_c_233_n 5.32086e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_87 N_A_M9_g N_Y_c_235_n 4.61191e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_88 N_A_c_89_n N_Y_c_235_n 7.74107e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_89 N_A_M10_g N_Y_c_237_n 2.64606e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_90 A N_Y_c_237_n 0.0012482f $X=0.621 $Y=0.138 $X2=0 $Y2=0
cc_91 N_A_c_89_n N_Y_c_228_n 4.94606e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_92 N_A_M10_g N_Y_c_240_n 2.77224e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_93 A N_Y_c_240_n 0.00123371f $X=0.621 $Y=0.138 $X2=0 $Y2=0
cc_94 N_A_c_89_n N_Y_c_242_n 8.61062e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_95 N_A_M11_g N_Y_c_243_n 4.5732e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_96 A Y 8.29133e-19 $X=0.621 $Y=0.138 $X2=0 $Y2=0
cc_97 A N_Y_c_245_n 8.29133e-19 $X=0.621 $Y=0.138 $X2=0 $Y2=0
cc_98 N_7_c_120_n N_8_c_142_n 0.00379429f $X=0.216 $Y=0.036 $X2=0.081 $Y2=0.135
cc_99 N_7_c_122_n N_8_c_142_n 0.00250918f $X=0.324 $Y=0.036 $X2=0.081 $Y2=0.135
cc_100 N_7_c_123_n N_8_c_142_n 0.00361461f $X=0.324 $Y=0.036 $X2=0.081 $Y2=0.135
cc_101 N_7_c_122_n N_8_c_158_n 4.51105e-19 $X=0.324 $Y=0.036 $X2=0.135
+ $Y2=0.0675
cc_102 N_7_c_123_n N_8_c_158_n 0.0032677f $X=0.324 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_103 N_7_c_120_n N_8_c_144_n 2.68768e-19 $X=0.216 $Y=0.036 $X2=0.189 $Y2=0.216
cc_104 N_7_c_122_n N_8_c_144_n 0.00723013f $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.216
cc_105 N_7_c_123_n N_8_c_146_n 0.00233206f $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_106 N_7_c_122_n N_9_c_175_n 3.33393e-19 $X=0.324 $Y=0.036 $X2=0.189 $Y2=0.216
cc_107 N_7_c_116_n N_Y_c_205_n 9.19308e-19 $X=0.108 $Y=0.036 $X2=0.135 $Y2=0.216
cc_108 N_7_c_120_n N_Y_c_247_n 7.34324e-19 $X=0.216 $Y=0.036 $X2=0.189 $Y2=0.135
cc_109 N_7_c_123_n N_Y_c_210_n 9.98826e-19 $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_110 N_7_c_114_n N_Y_c_206_n 2.27785e-19 $X=0.108 $Y=0.036 $X2=0 $Y2=0
cc_111 N_7_c_117_n N_Y_c_206_n 2.27785e-19 $X=0.207 $Y=0.036 $X2=0 $Y2=0
cc_112 N_8_c_158_n N_9_c_173_n 0.00317784f $X=0.378 $Y=0.0675 $X2=0.351
+ $Y2=0.0675
cc_113 N_8_c_149_n N_9_c_173_n 0.00358852f $X=0.486 $Y=0.0675 $X2=0.351
+ $Y2=0.0675
cc_114 N_8_c_165_p N_9_c_173_n 0.00233206f $X=0.4485 $Y=0.072 $X2=0.351
+ $Y2=0.0675
cc_115 N_8_c_149_n N_9_c_174_n 0.00363127f $X=0.486 $Y=0.0675 $X2=0.351
+ $Y2=0.216
cc_116 N_8_c_151_n N_9_c_174_n 3.19711e-19 $X=0.485 $Y=0.072 $X2=0.351 $Y2=0.216
cc_117 N_8_c_158_n N_9_c_175_n 4.73069e-19 $X=0.378 $Y=0.0675 $X2=0.351
+ $Y2=0.216
cc_118 N_8_c_149_n N_9_c_175_n 0.00250051f $X=0.486 $Y=0.0675 $X2=0.351
+ $Y2=0.216
cc_119 N_8_c_165_p N_9_c_175_n 0.00744433f $X=0.4485 $Y=0.072 $X2=0.351
+ $Y2=0.216
cc_120 N_8_c_146_n N_Y_c_218_n 0.00103693f $X=0.34 $Y=0.072 $X2=0 $Y2=0
cc_121 N_9_c_174_n N_Y_c_230_n 0.00362498f $X=0.54 $Y=0.036 $X2=0.405 $Y2=0.135
cc_122 N_9_c_181_n N_Y_c_230_n 0.00250914f $X=0.648 $Y=0.036 $X2=0.405 $Y2=0.135
cc_123 N_9_c_182_n N_Y_c_230_n 0.00348914f $X=0.648 $Y=0.036 $X2=0.405 $Y2=0.135
cc_124 N_9_c_181_n N_Y_c_255_n 2.9219e-19 $X=0.648 $Y=0.036 $X2=0.459 $Y2=0.0675
cc_125 N_9_c_182_n N_Y_c_255_n 0.00339247f $X=0.648 $Y=0.036 $X2=0.459
+ $Y2=0.0675
cc_126 N_9_c_173_n N_Y_c_220_n 9.98826e-19 $X=0.432 $Y=0.036 $X2=0 $Y2=0
cc_127 N_9_c_174_n N_Y_c_221_n 7.31912e-19 $X=0.54 $Y=0.036 $X2=0.513 $Y2=0.135
cc_128 N_9_c_182_n N_Y_c_231_n 9.98826e-19 $X=0.648 $Y=0.036 $X2=0 $Y2=0
cc_129 N_9_c_174_n N_Y_c_228_n 3.22784e-19 $X=0.54 $Y=0.036 $X2=0 $Y2=0
cc_130 N_9_c_181_n N_Y_c_228_n 0.00739153f $X=0.648 $Y=0.036 $X2=0 $Y2=0
cc_131 N_9_c_182_n N_Y_c_242_n 0.00233206f $X=0.648 $Y=0.036 $X2=0 $Y2=0

* END of "./NAND4xp75_ASAP7_75t_R.pex.sp.NAND4XP75_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NAND5xp2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:42:05 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NAND5xp2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NAND5xp2_ASAP7_75t_R.pex.sp.pex"
* File: NAND5xp2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:42:05 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NAND5XP2_ASAP7_75T_R%A 2 5 7 13 VSS
c10 13 VSS 0.00172694f $X=0.081 $Y=0.135
c11 5 VSS 0.00325747f $X=0.081 $Y=0.134
c12 2 VSS 0.0653596f $X=0.081 $Y=0.0675
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.134 $X2=0.081
+ $Y2=0.134
r14 5 7 307.213 $w=2e-08 $l=8.2e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.134 $X2=0.081 $Y2=0.216
r15 2 5 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.134
.ends

.subckt PM_NAND5XP2_ASAP7_75T_R%B 2 5 7 15 VSS
c12 15 VSS 0.0024522f $X=0.135 $Y=0.135
c13 5 VSS 0.0017107f $X=0.135 $Y=0.1345
c14 2 VSS 0.0604599f $X=0.135 $Y=0.0675
r15 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.134 $X2=0.135
+ $Y2=0.134
r16 5 7 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1345 $X2=0.135 $Y2=0.216
r17 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1345
.ends

.subckt PM_NAND5XP2_ASAP7_75T_R%C 2 5 7 13 VSS
c11 13 VSS 0.00220204f $X=0.189 $Y=0.135
c12 5 VSS 0.00160244f $X=0.189 $Y=0.1345
c13 2 VSS 0.0597904f $X=0.189 $Y=0.0675
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.134 $X2=0.189
+ $Y2=0.134
r15 5 7 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1345 $X2=0.189 $Y2=0.216
r16 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.1345
.ends

.subckt PM_NAND5XP2_ASAP7_75T_R%D 2 5 7 13 VSS
c10 13 VSS 0.00239098f $X=0.243 $Y=0.135
c11 5 VSS 0.0016285f $X=0.243 $Y=0.1345
c12 2 VSS 0.0597219f $X=0.243 $Y=0.0675
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.134 $X2=0.243
+ $Y2=0.134
r14 5 7 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1345 $X2=0.243 $Y2=0.216
r15 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.1345
.ends

.subckt PM_NAND5XP2_ASAP7_75T_R%E 2 5 7 13 VSS
c7 13 VSS 0.00581766f $X=0.297 $Y=0.135
c8 5 VSS 0.00255331f $X=0.297 $Y=0.1345
c9 2 VSS 0.0624574f $X=0.297 $Y=0.0675
r10 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.134 $X2=0.297
+ $Y2=0.134
r11 5 7 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.1345 $X2=0.297 $Y2=0.216
r12 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.1345
.ends

.subckt PM_NAND5XP2_ASAP7_75T_R%Y 1 6 9 11 12 15 16 17 20 24 26 31 32 43 45 48
+ 51 53 VSS
c20 53 VSS 0.00146362f $X=0.252 $Y=0.234
c21 52 VSS 0.00631462f $X=0.234 $Y=0.234
c22 51 VSS 0.00146362f $X=0.198 $Y=0.234
c23 50 VSS 0.00284382f $X=0.18 $Y=0.234
c24 48 VSS 0.00904588f $X=0.27 $Y=0.234
c25 46 VSS 9.64186e-19 $X=0.153 $Y=0.234
c26 45 VSS 0.00142296f $X=0.144 $Y=0.234
c27 44 VSS 0.00636214f $X=0.126 $Y=0.234
c28 43 VSS 0.00142296f $X=0.09 $Y=0.234
c29 42 VSS 1.68773e-19 $X=0.072 $Y=0.234
c30 41 VSS 0.00470185f $X=0.07 $Y=0.234
c31 34 VSS 0.00324955f $X=0.027 $Y=0.234
c32 32 VSS 0.00244555f $X=0.054 $Y=0.036
c33 31 VSS 0.00545273f $X=0.054 $Y=0.036
c34 29 VSS 0.00317163f $X=0.027 $Y=0.036
c35 28 VSS 4.98571e-19 $X=0.018 $Y=0.2125
c36 26 VSS 0.00127013f $X=0.018 $Y=0.0995
c37 25 VSS 0.00117262f $X=0.018 $Y=0.07
c38 24 VSS 0.00478829f $X=0.025 $Y=0.129
c39 22 VSS 5.68738e-19 $X=0.018 $Y=0.225
c40 20 VSS 0.00791579f $X=0.27 $Y=0.216
c41 16 VSS 5.3314e-19 $X=0.287 $Y=0.216
c42 15 VSS 0.00792006f $X=0.162 $Y=0.216
c43 11 VSS 5.3314e-19 $X=0.179 $Y=0.216
c44 9 VSS 0.00523518f $X=0.056 $Y=0.216
c45 6 VSS 2.53241e-19 $X=0.071 $Y=0.216
c46 1 VSS 4.49354e-19 $X=0.071 $Y=0.0675
r47 52 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r48 51 52 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.234 $Y2=0.234
r49 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r50 48 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.252 $Y2=0.234
r51 45 46 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.153 $Y2=0.234
r52 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r53 43 44 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.126 $Y2=0.234
r54 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r55 41 42 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.07
+ $Y=0.234 $X2=0.072 $Y2=0.234
r56 39 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r57 39 46 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.153 $Y2=0.234
r58 36 41 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.07 $Y2=0.234
r59 34 36 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.054 $Y2=0.234
r60 31 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r61 29 31 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.054 $Y2=0.036
r62 27 28 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.2 $X2=0.018 $Y2=0.2125
r63 25 26 2.00309 $w=1.8e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.0995
r64 24 27 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.129 $X2=0.018 $Y2=0.2
r65 24 26 2.00309 $w=1.8e-08 $l=2.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.129 $X2=0.018 $Y2=0.0995
r66 22 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r67 22 28 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2125
r68 21 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r69 21 25 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r70 20 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r71 17 20 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.216 $X2=0.27 $Y2=0.216
r72 16 20 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.216 $X2=0.27 $Y2=0.216
r73 15 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r74 12 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.162 $Y2=0.216
r75 11 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.216 $X2=0.162 $Y2=0.216
r76 9 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r77 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.216 $X2=0.056 $Y2=0.216
r78 4 32 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r79 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends

.subckt PM_NAND5XP2_ASAP7_75T_R%9 1 2 VSS
c0 1 VSS 0.00228332f $X=0.125 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends

.subckt PM_NAND5XP2_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00228332f $X=0.179 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.145 $Y2=0.0675
.ends

.subckt PM_NAND5XP2_ASAP7_75T_R%11 1 2 VSS
c0 1 VSS 0.00228332f $X=0.233 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.199 $Y2=0.0675
.ends

.subckt PM_NAND5XP2_ASAP7_75T_R%12 1 2 VSS
c0 1 VSS 0.00228332f $X=0.287 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.253 $Y2=0.0675
.ends


* END of "./NAND5xp2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NAND5xp2_ASAP7_75t_R  VSS VDD A B C D E Y
* 
* Y	Y
* E	E
* D	D
* C	C
* B	B
* A	A
M0 N_9_M0_d N_A_M0_g N_Y_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_10_M1_d N_B_M1_g N_9_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_11_M2_d N_C_M2_g N_10_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_12_M3_d N_D_M3_g N_11_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 VSS N_E_M4_g N_12_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 VDD N_A_M5_g N_Y_M5_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M6 N_Y_M6_d N_B_M6_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
M7 VDD N_C_M7_g N_Y_M7_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.189
M8 N_Y_M8_d N_D_M8_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.189
M9 VDD N_E_M9_g N_Y_M9_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287 $Y=0.189
*
* 
* .include "NAND5xp2_ASAP7_75t_R.pex.sp.NAND5XP2_ASAP7_75T_R.pxi"
* BEGIN of "./NAND5xp2_ASAP7_75t_R.pex.sp.NAND5XP2_ASAP7_75T_R.pxi"
* File: NAND5xp2_ASAP7_75t_R.pex.sp.NAND5XP2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:42:05 2017
* 
x_PM_NAND5XP2_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M5_g A VSS
+ PM_NAND5XP2_ASAP7_75T_R%A
x_PM_NAND5XP2_ASAP7_75T_R%B N_B_M1_g N_B_c_12_n N_B_M6_g B VSS
+ PM_NAND5XP2_ASAP7_75T_R%B
x_PM_NAND5XP2_ASAP7_75T_R%C N_C_M2_g N_C_c_25_n N_C_M7_g C VSS
+ PM_NAND5XP2_ASAP7_75T_R%C
x_PM_NAND5XP2_ASAP7_75T_R%D N_D_M3_g N_D_c_36_n N_D_M8_g D VSS
+ PM_NAND5XP2_ASAP7_75T_R%D
x_PM_NAND5XP2_ASAP7_75T_R%E N_E_M4_g N_E_c_46_n N_E_M9_g E VSS
+ PM_NAND5XP2_ASAP7_75T_R%E
x_PM_NAND5XP2_ASAP7_75T_R%Y N_Y_M0_s N_Y_M5_s N_Y_c_51_n N_Y_M7_s N_Y_M6_d
+ N_Y_c_57_n N_Y_M9_s N_Y_M8_d N_Y_c_65_n Y N_Y_c_52_n N_Y_c_58_n N_Y_c_53_n
+ N_Y_c_55_n N_Y_c_60_n N_Y_c_69_n N_Y_c_63_n N_Y_c_66_n VSS
+ PM_NAND5XP2_ASAP7_75T_R%Y
x_PM_NAND5XP2_ASAP7_75T_R%9 N_9_M1_s N_9_M0_d VSS PM_NAND5XP2_ASAP7_75T_R%9
x_PM_NAND5XP2_ASAP7_75T_R%10 N_10_M2_s N_10_M1_d VSS PM_NAND5XP2_ASAP7_75T_R%10
x_PM_NAND5XP2_ASAP7_75T_R%11 N_11_M3_s N_11_M2_d VSS PM_NAND5XP2_ASAP7_75T_R%11
x_PM_NAND5XP2_ASAP7_75T_R%12 N_12_M4_s N_12_M3_d VSS PM_NAND5XP2_ASAP7_75T_R%12
cc_1 N_A_M0_g N_B_M1_g 0.00333077f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_12_n 7.98811e-19 $X=0.081 $Y=0.134 $X2=0.135 $Y2=0.1345
cc_3 A B 0.00621434f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A_M0_g N_C_M2_g 2.71887e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 A N_Y_c_51_n 3.52002e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_6 A N_Y_c_52_n 0.00436078f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_7 N_A_c_2_p N_Y_c_53_n 3.06446e-19 $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_8 A N_Y_c_53_n 0.00134508f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_A_M0_g N_Y_c_55_n 2.57864e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_10 A N_Y_c_55_n 0.00123648f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 N_B_M1_g N_C_M2_g 0.00357042f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_12 N_B_c_12_n N_C_c_25_n 7.92653e-19 $X=0.135 $Y=0.1345 $X2=0.081 $Y2=0.134
cc_13 B C 0.00817592f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 N_B_M1_g N_D_M3_g 2.71887e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_15 B N_Y_c_57_n 3.31541e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_16 B N_Y_c_58_n 4.64233e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_17 B N_Y_c_53_n 5.56013e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_18 N_B_M1_g N_Y_c_60_n 2.57565e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 B N_Y_c_60_n 0.00123952f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_20 N_C_M2_g N_D_M3_g 0.00327995f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_21 N_C_c_25_n N_D_c_36_n 7.90494e-19 $X=0.189 $Y=0.1345 $X2=0.081 $Y2=0.134
cc_22 C D 0.00819209f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 N_C_M2_g N_E_M4_g 2.66145e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_24 C N_Y_c_57_n 3.31541e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_25 N_C_M2_g N_Y_c_63_n 2.64924e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 C N_Y_c_63_n 0.00125705f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_27 N_D_M3_g N_E_M4_g 0.00344695f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_28 N_D_c_36_n N_E_c_46_n 8.31912e-19 $X=0.243 $Y=0.1345 $X2=0.135 $Y2=0.1345
cc_29 D E 0.00809651f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_30 D N_Y_c_65_n 3.31541e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 N_D_M3_g N_Y_c_66_n 2.64924e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_32 D N_Y_c_66_n 0.00125705f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_33 E N_Y_c_65_n 3.31541e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_34 N_E_M4_g N_Y_c_69_n 2.63571e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_35 E N_Y_c_69_n 0.00125705f $X=0.297 $Y=0.135 $X2=0 $Y2=0

* END of "./NAND5xp2_ASAP7_75t_R.pex.sp.NAND5XP2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR2x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:42:27 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR2x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR2x1_ASAP7_75t_R.pex.sp.pex"
* File: NOR2x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:42:27 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR2X1_ASAP7_75T_R%A 2 5 8 11 13 23 VSS
c17 23 VSS 0.0172609f $X=0.07 $Y=0.134
c18 11 VSS 0.00965183f $X=0.135 $Y=0.1355
c19 8 VSS 0.0631147f $X=0.135 $Y=0.0675
c20 2 VSS 0.0689981f $X=0.081 $Y=0.1355
r21 23 27 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.07 $Y=0.135 $X2=0.07
+ $Y2=0.135
r22 11 13 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.2025
r23 8 11 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1355
r24 2 11 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1355 $X2=0.135 $Y2=0.1355
r25 2 27 9.56522 $w=2.3e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1355 $X2=0.07 $Y2=0.1355
r26 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1355 $X2=0.081 $Y2=0.2025
.ends

.subckt PM_NOR2X1_ASAP7_75T_R%B 2 7 10 13 21 VSS
c28 21 VSS 0.0066475f $X=0.215 $Y=0.134
c29 10 VSS 0.072767f $X=0.243 $Y=0.135
c30 2 VSS 0.0623886f $X=0.189 $Y=0.0675
r31 21 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.216 $Y=0.135 $X2=0.216
+ $Y2=0.135
r32 10 25 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.216 $Y2=0.135
r33 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r34 5 25 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.216 $Y2=0.135
r35 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r36 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_NOR2X1_ASAP7_75T_R%5 1 4 6 7 10 11 14 17 25 28 30 32 33 VSS
c19 33 VSS 0.00267294f $X=0.236 $Y=0.234
c20 32 VSS 0.00469192f $X=0.202 $Y=0.234
c21 30 VSS 0.00500972f $X=0.27 $Y=0.234
c22 28 VSS 0.00429696f $X=0.144 $Y=0.234
c23 27 VSS 0.00231585f $X=0.107 $Y=0.234
c24 26 VSS 9.61037e-19 $X=0.094 $Y=0.234
c25 25 VSS 0.00270713f $X=0.084 $Y=0.234
c26 17 VSS 0.00190113f $X=0.054 $Y=0.234
c27 14 VSS 0.00266486f $X=0.268 $Y=0.2025
c28 10 VSS 0.00699137f $X=0.162 $Y=0.2025
c29 6 VSS 7.1893e-19 $X=0.179 $Y=0.2025
c30 4 VSS 0.00621518f $X=0.056 $Y=0.2025
c31 1 VSS 4.64427e-19 $X=0.071 $Y=0.2025
r32 32 33 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.234 $X2=0.236 $Y2=0.234
r33 30 33 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.236 $Y2=0.234
r34 27 28 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.234 $X2=0.144 $Y2=0.234
r35 26 27 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.234 $X2=0.107 $Y2=0.234
r36 25 26 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.084
+ $Y=0.234 $X2=0.094 $Y2=0.234
r37 23 32 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.202 $Y2=0.234
r38 23 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.144 $Y2=0.234
r39 17 25 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.084 $Y2=0.234
r40 14 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r41 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.268 $Y2=0.2025
r42 10 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r43 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r44 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r45 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r46 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
.ends

.subckt PM_NOR2X1_ASAP7_75T_R%Y 1 6 11 12 15 18 19 26 27 28 29 35 36 38 40 42 44
+ VSS
c28 44 VSS 7.82225e-19 $X=0.297 $Y=0.144
c29 42 VSS 0.00145953f $X=0.297 $Y=0.094
c30 41 VSS 0.00104959f $X=0.297 $Y=0.063
c31 40 VSS 0.00168609f $X=0.298 $Y=0.125
c32 38 VSS 0.00224035f $X=0.297 $Y=0.189
c33 36 VSS 3.80778e-19 $X=0.284 $Y=0.198
c34 35 VSS 7.56861e-20 $X=0.23 $Y=0.198
c35 30 VSS 0.00215853f $X=0.288 $Y=0.198
c36 29 VSS 0.00275922f $X=0.259 $Y=0.036
c37 28 VSS 0.00393886f $X=0.23 $Y=0.036
c38 27 VSS 0.0057393f $X=0.18 $Y=0.036
c39 26 VSS 0.00286718f $X=0.144 $Y=0.036
c40 25 VSS 0.00609008f $X=0.216 $Y=0.036
c41 19 VSS 0.00816231f $X=0.108 $Y=0.036
c42 18 VSS 0.00195467f $X=0.108 $Y=0.036
c43 16 VSS 0.00628356f $X=0.288 $Y=0.036
c44 15 VSS 0.00288208f $X=0.216 $Y=0.2025
c45 11 VSS 5.71396e-19 $X=0.233 $Y=0.2025
c46 9 VSS 4.5957e-19 $X=0.214 $Y=0.0675
c47 1 VSS 5.07509e-19 $X=0.125 $Y=0.0675
r48 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.144
r49 41 42 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.063 $X2=0.297 $Y2=0.094
r50 40 43 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.125 $X2=0.297 $Y2=0.126
r51 40 42 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.125 $X2=0.297 $Y2=0.094
r52 38 44 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.144
r53 37 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.063
r54 35 36 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.198 $X2=0.284 $Y2=0.198
r55 32 35 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.23 $Y2=0.198
r56 30 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.198 $X2=0.297 $Y2=0.189
r57 30 36 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.284 $Y2=0.198
r58 28 29 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.036 $X2=0.259 $Y2=0.036
r59 26 27 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.18 $Y2=0.036
r60 24 28 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.23 $Y2=0.036
r61 24 27 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.18 $Y2=0.036
r62 24 25 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r63 18 26 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.144 $Y2=0.036
r64 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r65 16 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r66 16 29 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.259 $Y2=0.036
r67 15 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r68 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r69 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r70 9 25 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r71 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.214 $Y2=0.0675
r72 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r73 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.11 $Y2=0.0675
.ends


* END of "./NOR2x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR2x1_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 VSS N_A_M0_g N_Y_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M1 N_Y_M1_d N_B_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M2 VDD N_A_M2_g N_5_M2_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M3 VDD N_A_M3_g N_5_M3_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M4 N_Y_M4_d N_B_M4_g N_5_M4_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M5 N_Y_M5_d N_B_M5_g N_5_M5_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
*
* 
* .include "NOR2x1_ASAP7_75t_R.pex.sp.NOR2X1_ASAP7_75T_R.pxi"
* BEGIN of "./NOR2x1_ASAP7_75t_R.pex.sp.NOR2X1_ASAP7_75T_R.pxi"
* File: NOR2x1_ASAP7_75t_R.pex.sp.NOR2X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:42:27 2017
* 
x_PM_NOR2X1_ASAP7_75T_R%A N_A_c_1_p N_A_M2_g N_A_M0_g N_A_c_4_p N_A_M3_g A VSS
+ PM_NOR2X1_ASAP7_75T_R%A
x_PM_NOR2X1_ASAP7_75T_R%B N_B_M1_g N_B_M4_g N_B_c_20_n N_B_M5_g B VSS
+ PM_NOR2X1_ASAP7_75T_R%B
x_PM_NOR2X1_ASAP7_75T_R%5 N_5_M2_s N_5_c_46_n N_5_M4_s N_5_M3_s N_5_c_52_n
+ N_5_M5_s N_5_c_58_p N_5_c_47_n N_5_c_48_n N_5_c_51_n N_5_c_54_n N_5_c_55_n
+ N_5_c_59_p VSS PM_NOR2X1_ASAP7_75T_R%5
x_PM_NOR2X1_ASAP7_75T_R%Y N_Y_M0_s N_Y_M1_d N_Y_M5_d N_Y_M4_d N_Y_c_85_n
+ N_Y_c_65_n N_Y_c_66_n N_Y_c_68_n N_Y_c_72_n N_Y_c_74_n N_Y_c_76_n N_Y_c_77_n
+ N_Y_c_79_n N_Y_c_80_n Y N_Y_c_83_n N_Y_c_84_n VSS PM_NOR2X1_ASAP7_75T_R%Y
cc_1 N_A_c_1_p N_B_M1_g 2.31381e-19 $X=0.081 $Y=0.1355 $X2=0.189 $Y2=0.0675
cc_2 N_A_M0_g N_B_M1_g 0.0032073f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A_M0_g N_B_c_20_n 2.66145e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_4 N_A_c_4_p N_B_c_20_n 0.00207153f $X=0.135 $Y=0.1355 $X2=0.243 $Y2=0.135
cc_5 N_A_M0_g B 6.63451e-19 $X=0.135 $Y=0.0675 $X2=0.215 $Y2=0.134
cc_6 N_A_c_4_p B 0.0033047f $X=0.135 $Y=0.1355 $X2=0.215 $Y2=0.134
cc_7 A B 0.002325f $X=0.07 $Y=0.134 $X2=0.215 $Y2=0.134
cc_8 A N_5_c_46_n 0.00201602f $X=0.07 $Y=0.134 $X2=0.189 $Y2=0.135
cc_9 A N_5_c_47_n 0.00116786f $X=0.07 $Y=0.134 $X2=0 $Y2=0
cc_10 N_A_c_1_p N_5_c_48_n 2.7229e-19 $X=0.081 $Y=0.1355 $X2=0.216 $Y2=0.135
cc_11 N_A_c_4_p N_5_c_48_n 4.85349e-19 $X=0.135 $Y=0.1355 $X2=0.216 $Y2=0.135
cc_12 A N_5_c_48_n 2.11212e-19 $X=0.07 $Y=0.134 $X2=0.216 $Y2=0.135
cc_13 N_A_M0_g N_5_c_51_n 2.38073e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_14 A N_Y_c_65_n 8.40589e-19 $X=0.07 $Y=0.134 $X2=0 $Y2=0
cc_15 N_A_c_4_p N_Y_c_66_n 8.01479e-19 $X=0.135 $Y=0.1355 $X2=0 $Y2=0
cc_16 A N_Y_c_66_n 0.0011434f $X=0.07 $Y=0.134 $X2=0 $Y2=0
cc_17 N_A_M0_g N_Y_c_68_n 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_18 B N_5_c_52_n 0.00125734f $X=0.215 $Y=0.134 $X2=0.135 $Y2=0.1355
cc_19 B N_5_c_51_n 0.00377172f $X=0.215 $Y=0.134 $X2=0 $Y2=0
cc_20 N_B_c_20_n N_5_c_54_n 2.21754e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_21 N_B_M1_g N_5_c_55_n 4.28653e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_22 B N_5_c_55_n 0.0010249f $X=0.215 $Y=0.134 $X2=0 $Y2=0
cc_23 N_B_c_20_n N_Y_M5_d 3.80404e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.1355
cc_24 B N_Y_c_66_n 0.00224872f $X=0.215 $Y=0.134 $X2=0 $Y2=0
cc_25 B N_Y_c_68_n 0.00377239f $X=0.215 $Y=0.134 $X2=0.07 $Y2=0.135
cc_26 N_B_c_20_n N_Y_c_72_n 4.02626e-19 $X=0.243 $Y=0.135 $X2=0.07 $Y2=0.135
cc_27 B N_Y_c_72_n 6.70107e-19 $X=0.215 $Y=0.134 $X2=0.07 $Y2=0.135
cc_28 N_B_M1_g N_Y_c_74_n 4.01862e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_29 B N_Y_c_74_n 6.70107e-19 $X=0.215 $Y=0.134 $X2=0 $Y2=0
cc_30 N_B_c_20_n N_Y_c_76_n 4.59758e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_31 N_B_c_20_n N_Y_c_77_n 5.08727e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_32 B N_Y_c_77_n 0.00101392f $X=0.215 $Y=0.134 $X2=0 $Y2=0
cc_33 N_B_c_20_n N_Y_c_79_n 3.95625e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.1355
cc_34 B N_Y_c_80_n 2.20656e-19 $X=0.215 $Y=0.134 $X2=0 $Y2=0
cc_35 N_B_c_20_n Y 4.69449e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_36 B Y 2.00696e-19 $X=0.215 $Y=0.134 $X2=0 $Y2=0
cc_37 B N_Y_c_83_n 2.00696e-19 $X=0.215 $Y=0.134 $X2=0 $Y2=0
cc_38 B N_Y_c_84_n 4.07779e-19 $X=0.215 $Y=0.134 $X2=0 $Y2=0
cc_39 N_5_c_52_n N_Y_c_85_n 0.00367277f $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_40 N_5_c_58_p N_Y_c_85_n 0.00368895f $X=0.268 $Y=0.2025 $X2=0 $Y2=0
cc_41 N_5_c_59_p N_Y_c_85_n 0.0025091f $X=0.236 $Y=0.234 $X2=0 $Y2=0
cc_42 N_5_c_52_n N_Y_c_77_n 3.96143e-19 $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_43 N_5_c_59_p N_Y_c_77_n 0.00353849f $X=0.236 $Y=0.234 $X2=0 $Y2=0
cc_44 N_5_c_58_p N_Y_c_79_n 0.00285496f $X=0.268 $Y=0.2025 $X2=0.081 $Y2=0.1355
cc_45 N_5_c_54_n N_Y_c_79_n 0.00353849f $X=0.27 $Y=0.234 $X2=0.081 $Y2=0.1355
cc_46 N_5_c_58_p N_Y_c_80_n 3.52384e-19 $X=0.268 $Y=0.2025 $X2=0 $Y2=0

* END of "./NOR2x1_ASAP7_75t_R.pex.sp.NOR2X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR2x1p5_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:42:49 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR2x1p5_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR2x1p5_ASAP7_75t_R.pex.sp.pex"
* File: NOR2x1p5_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:42:49 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR2X1P5_ASAP7_75T_R%A 5 8 13 16 19 21 37 VSS
c22 37 VSS 0.0246493f $X=0.07 $Y=0.136
c23 19 VSS 0.0122813f $X=0.189 $Y=0.1355
c24 16 VSS 0.0622543f $X=0.189 $Y=0.054
c25 8 VSS 0.0638575f $X=0.135 $Y=0.0675
c26 2 VSS 0.067082f $X=0.081 $Y=0.1355
r27 34 37 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.07 $Y=0.135 $X2=0.07
+ $Y2=0.135
r28 19 21 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1355 $X2=0.189 $Y2=0.2025
r29 16 19 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.1355
r30 11 19 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.1355 $X2=0.189 $Y2=0.1355
r31 11 13 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.2025
r32 8 11 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1355
r33 2 11 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1355 $X2=0.135 $Y2=0.1355
r34 2 34 9.56522 $w=2.3e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1355 $X2=0.07 $Y2=0.1355
r35 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1355 $X2=0.081 $Y2=0.2025
.ends

.subckt PM_NOR2X1P5_ASAP7_75T_R%B 2 7 10 15 18 21 29 31 32 39 VSS
c33 39 VSS 0.00657098f $X=0.135 $Y=0.136
c34 32 VSS 1.63059e-19 $X=0.202 $Y=0.135
c35 31 VSS 1.06681e-21 $X=0.163 $Y=0.135
c36 29 VSS 6.5551e-19 $X=0.243 $Y=0.135
c37 18 VSS 0.0770878f $X=0.351 $Y=0.135
c38 10 VSS 0.0645037f $X=0.297 $Y=0.0675
c39 2 VSS 0.0621762f $X=0.243 $Y=0.054
r40 31 32 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.163
+ $Y=0.135 $X2=0.202 $Y2=0.135
r41 29 32 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.202 $Y2=0.135
r42 27 39 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.135 $Y2=0.135
r43 27 31 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.135 $X2=0.163 $Y2=0.135
r44 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r45 13 18 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r46 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r47 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r48 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r49 5 29 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r50 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r51 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_NOR2X1P5_ASAP7_75T_R%5 1 2 5 6 7 10 11 12 15 17 23 25 26 33 35 36 37
+ 38 VSS
c29 38 VSS 5.12412e-19 $X=0.2925 $Y=0.198
c30 37 VSS 2.79488e-19 $X=0.261 $Y=0.198
c31 36 VSS 9.73694e-19 $X=0.257 $Y=0.198
c32 35 VSS 4.97766e-19 $X=0.225 $Y=0.198
c33 33 VSS 2.92324e-19 $X=0.324 $Y=0.198
c34 26 VSS 0.0074475f $X=0.202 $Y=0.234
c35 25 VSS 0.00286574f $X=0.144 $Y=0.234
c36 23 VSS 0.0022696f $X=0.216 $Y=0.234
c37 17 VSS 0.0021938f $X=0.108 $Y=0.234
c38 15 VSS 0.0026225f $X=0.324 $Y=0.2025
c39 11 VSS 5.75221e-19 $X=0.341 $Y=0.2025
c40 10 VSS 0.00603836f $X=0.216 $Y=0.2025
c41 6 VSS 7.04766e-19 $X=0.233 $Y=0.2025
c42 5 VSS 0.0105454f $X=0.108 $Y=0.2025
c43 1 VSS 6.18024e-19 $X=0.125 $Y=0.2025
r44 37 38 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.198 $X2=0.2925 $Y2=0.198
r45 36 37 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.257
+ $Y=0.198 $X2=0.261 $Y2=0.198
r46 35 36 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.198 $X2=0.257 $Y2=0.198
r47 33 38 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.2925 $Y2=0.198
r48 29 35 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.225 $Y2=0.198
r49 25 26 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.202 $Y2=0.234
r50 23 26 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.202 $Y2=0.234
r51 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r52 17 25 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.144 $Y2=0.234
r53 15 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198 $X2=0.324
+ $Y2=0.198
r54 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r55 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r56 10 24 31.0714 $w=2.4e-08 $l=3.6e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.198 $X2=0.216 $Y2=0.234
r57 10 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r58 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r59 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r60 5 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r61 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.2025 $X2=0.108 $Y2=0.2025
r62 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.108 $Y2=0.2025
.ends

.subckt PM_NOR2X1P5_ASAP7_75T_R%Y 1 6 7 10 11 16 17 20 21 24 28 29 37 40 41 43
+ 44 53 54 58 61 64 VSS
c32 64 VSS 6.86417e-19 $X=0.405 $Y=0.207
c33 62 VSS 9.22213e-19 $X=0.405 $Y=0.144
c34 61 VSS 0.00243102f $X=0.405 $Y=0.126
c35 60 VSS 7.83596e-19 $X=0.405 $Y=0.081
c36 59 VSS 0.00104959f $X=0.405 $Y=0.063
c37 58 VSS 0.00237618f $X=0.405 $Y=0.145
c38 56 VSS 8.85605e-19 $X=0.405 $Y=0.225
c39 54 VSS 0.00175149f $X=0.358 $Y=0.234
c40 53 VSS 0.00657771f $X=0.338 $Y=0.234
c41 45 VSS 0.00707768f $X=0.396 $Y=0.234
c42 44 VSS 0.00266146f $X=0.367 $Y=0.036
c43 43 VSS 0.00425376f $X=0.338 $Y=0.036
c44 42 VSS 0.00567501f $X=0.2905 $Y=0.036
c45 41 VSS 0.0089446f $X=0.257 $Y=0.036
c46 40 VSS 0.00626831f $X=0.324 $Y=0.036
c47 37 VSS 0.00429709f $X=0.163 $Y=0.036
c48 36 VSS 0.00163196f $X=0.126 $Y=0.036
c49 29 VSS 0.00671331f $X=0.108 $Y=0.036
c50 28 VSS 0.00187319f $X=0.108 $Y=0.036
c51 26 VSS 0.00634021f $X=0.396 $Y=0.036
c52 24 VSS 0.00307995f $X=0.376 $Y=0.2025
c53 20 VSS 0.00488081f $X=0.27 $Y=0.2025
c54 16 VSS 6.56704e-19 $X=0.287 $Y=0.2025
c55 14 VSS 4.59792e-19 $X=0.322 $Y=0.0675
c56 10 VSS 0.00783498f $X=0.216 $Y=0.054
c57 6 VSS 5.3314e-19 $X=0.233 $Y=0.054
c58 1 VSS 4.6121e-19 $X=0.125 $Y=0.0675
r59 63 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.207
r60 61 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.126 $X2=0.405 $Y2=0.144
r61 60 61 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.081 $X2=0.405 $Y2=0.126
r62 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.063 $X2=0.405 $Y2=0.081
r63 58 63 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.145 $X2=0.405 $Y2=0.189
r64 58 62 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.145 $X2=0.405 $Y2=0.144
r65 56 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.207
r66 55 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.063
r67 53 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.234 $X2=0.358 $Y2=0.234
r68 51 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.358 $Y2=0.234
r69 47 53 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.338 $Y2=0.234
r70 45 56 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r71 45 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.378 $Y2=0.234
r72 43 44 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.036 $X2=0.367 $Y2=0.036
r73 41 42 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.257
+ $Y=0.036 $X2=0.2905 $Y2=0.036
r74 39 43 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.338 $Y2=0.036
r75 39 42 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.2905 $Y2=0.036
r76 39 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r77 36 37 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.163 $Y2=0.036
r78 34 41 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.257 $Y2=0.036
r79 34 37 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.163 $Y2=0.036
r80 28 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r81 28 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r82 26 55 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r83 26 44 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.367 $Y2=0.036
r84 24 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r85 21 24 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.376 $Y2=0.2025
r86 20 47 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r87 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r88 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r89 14 40 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r90 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.322 $Y2=0.0675
r91 10 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r92 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.054 $X2=0.216 $Y2=0.054
r93 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.054 $X2=0.216 $Y2=0.054
r94 4 29 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r95 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.11 $Y2=0.0675
.ends


* END of "./NOR2x1p5_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR2x1p5_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 VSS N_A_M0_g N_Y_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M1 VSS N_A_M1_g N_Y_M1_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M2 VSS N_B_M2_g N_Y_M2_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M3 VSS N_B_M3_g N_Y_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M4 N_5_M4_d N_A_M4_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M5 N_5_M5_d N_A_M5_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M6 N_5_M6_d N_A_M6_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M7 N_Y_M7_d N_B_M7_g N_5_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M8 N_Y_M8_d N_B_M8_g N_5_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M9 N_Y_M9_d N_B_M9_g N_5_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "NOR2x1p5_ASAP7_75t_R.pex.sp.NOR2X1P5_ASAP7_75T_R.pxi"
* BEGIN of "./NOR2x1p5_ASAP7_75t_R.pex.sp.NOR2X1P5_ASAP7_75T_R.pxi"
* File: NOR2x1p5_ASAP7_75t_R.pex.sp.NOR2X1P5_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:42:49 2017
* 
x_PM_NOR2X1P5_ASAP7_75T_R%A N_A_M4_g N_A_M0_g N_A_M5_g N_A_M1_g N_A_c_4_p
+ N_A_M6_g A VSS PM_NOR2X1P5_ASAP7_75T_R%A
x_PM_NOR2X1P5_ASAP7_75T_R%B N_B_M2_g N_B_M7_g N_B_M3_g N_B_M8_g N_B_c_26_n
+ N_B_M9_g N_B_c_39_p N_B_c_27_n N_B_c_28_n B VSS PM_NOR2X1P5_ASAP7_75T_R%B
x_PM_NOR2X1P5_ASAP7_75T_R%5 N_5_M5_d N_5_M4_d N_5_c_57_n N_5_M7_s N_5_M6_d
+ N_5_c_72_p N_5_M9_s N_5_M8_s N_5_c_64_n N_5_c_58_n N_5_c_82_p N_5_c_59_n
+ N_5_c_60_n N_5_c_67_n N_5_c_68_n N_5_c_70_n N_5_c_75_p N_5_c_76_p VSS
+ PM_NOR2X1P5_ASAP7_75T_R%5
x_PM_NOR2X1P5_ASAP7_75T_R%Y N_Y_M0_s N_Y_M2_s N_Y_M1_s N_Y_c_104_n N_Y_M3_s
+ N_Y_M8_d N_Y_M7_d N_Y_c_92_n N_Y_M9_d N_Y_c_109_n N_Y_c_85_n N_Y_c_87_n
+ N_Y_c_89_n N_Y_c_95_n N_Y_c_90_n N_Y_c_99_n N_Y_c_100_n N_Y_c_101_n
+ N_Y_c_102_n Y N_Y_c_103_n N_Y_c_116_n VSS PM_NOR2X1P5_ASAP7_75T_R%Y
cc_1 N_A_M0_g N_B_M2_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.054
cc_2 N_A_M1_g N_B_M2_g 0.00344695f $X=0.189 $Y=0.054 $X2=0.243 $Y2=0.054
cc_3 N_A_M1_g N_B_M3_g 2.66145e-19 $X=0.189 $Y=0.054 $X2=0.297 $Y2=0.0675
cc_4 N_A_c_4_p N_B_c_26_n 0.0020914f $X=0.189 $Y=0.1355 $X2=0.351 $Y2=0.135
cc_5 N_A_c_4_p N_B_c_27_n 0.00109734f $X=0.189 $Y=0.1355 $X2=0.163 $Y2=0.135
cc_6 N_A_M1_g N_B_c_28_n 7.24562e-19 $X=0.189 $Y=0.054 $X2=0.202 $Y2=0.135
cc_7 N_A_c_4_p N_B_c_28_n 0.00297492f $X=0.189 $Y=0.1355 $X2=0.202 $Y2=0.135
cc_8 N_A_M0_g B 6.18619e-19 $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.136
cc_9 N_A_c_4_p B 0.00239456f $X=0.189 $Y=0.1355 $X2=0.135 $Y2=0.136
cc_10 A B 0.00188437f $X=0.07 $Y=0.136 $X2=0.135 $Y2=0.136
cc_11 N_A_c_4_p N_5_M5_d 3.8991e-19 $X=0.189 $Y=0.1355 $X2=0.243 $Y2=0.054
cc_12 N_A_c_4_p N_5_c_57_n 8.45347e-19 $X=0.189 $Y=0.1355 $X2=0.243 $Y2=0.135
cc_13 A N_5_c_58_n 5.26979e-19 $X=0.07 $Y=0.136 $X2=0.351 $Y2=0.135
cc_14 N_A_M0_g N_5_c_59_n 2.34767e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 N_A_M1_g N_5_c_60_n 4.27122e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_16 N_A_c_4_p N_5_c_60_n 2.13568e-19 $X=0.189 $Y=0.1355 $X2=0 $Y2=0
cc_17 N_A_c_4_p N_Y_c_85_n 3.08716e-19 $X=0.189 $Y=0.1355 $X2=0.243 $Y2=0.135
cc_18 A N_Y_c_85_n 8.43259e-19 $X=0.07 $Y=0.136 $X2=0.243 $Y2=0.135
cc_19 N_A_c_4_p N_Y_c_87_n 8.01479e-19 $X=0.189 $Y=0.1355 $X2=0.243 $Y2=0.135
cc_20 A N_Y_c_87_n 0.0013808f $X=0.07 $Y=0.136 $X2=0.243 $Y2=0.135
cc_21 N_A_M0_g N_Y_c_89_n 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_22 N_A_M1_g N_Y_c_90_n 4.28653e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_23 B N_5_c_57_n 0.00216211f $X=0.135 $Y=0.136 $X2=0.081 $Y2=0.2025
cc_24 N_B_c_26_n N_5_M9_s 3.80371e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.1355
cc_25 N_B_c_26_n N_5_c_64_n 8.0006e-19 $X=0.351 $Y=0.135 $X2=0.189 $Y2=0.054
cc_26 B N_5_c_59_n 0.00372796f $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_27 N_B_c_27_n N_5_c_60_n 8.54443e-19 $X=0.163 $Y=0.135 $X2=0 $Y2=0
cc_28 N_B_M3_g N_5_c_67_n 2.83374e-19 $X=0.297 $Y=0.0675 $X2=0.07 $Y2=0.135
cc_29 N_B_c_39_p N_5_c_68_n 0.00189395f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_30 B N_5_c_68_n 3.68725e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_31 N_B_M2_g N_5_c_70_n 4.27107e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_32 N_B_c_26_n N_5_c_70_n 0.00133835f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_33 N_B_c_26_n N_Y_M8_d 3.80413e-19 $X=0.351 $Y=0.135 $X2=0.189 $Y2=0.054
cc_34 N_B_c_26_n N_Y_c_92_n 8.0006e-19 $X=0.351 $Y=0.135 $X2=0.189 $Y2=0.2025
cc_35 B N_Y_c_87_n 0.00157124f $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_36 B N_Y_c_89_n 0.00377179f $X=0.135 $Y=0.136 $X2=0.07 $Y2=0.136
cc_37 N_B_c_26_n N_Y_c_95_n 8.0006e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_38 N_B_M2_g N_Y_c_90_n 4.28653e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_39 N_B_c_26_n N_Y_c_90_n 0.00129524f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_40 N_B_c_28_n N_Y_c_90_n 0.00157481f $X=0.202 $Y=0.135 $X2=0 $Y2=0
cc_41 N_B_M3_g N_Y_c_99_n 3.58606e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_42 N_B_c_26_n N_Y_c_100_n 4.59284e-19 $X=0.351 $Y=0.135 $X2=0.07 $Y2=0.1355
cc_43 N_B_M3_g N_Y_c_101_n 2.64781e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_B_c_26_n N_Y_c_102_n 6.43639e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_45 N_B_c_26_n N_Y_c_103_n 3.35167e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_46 N_5_c_72_p N_Y_c_104_n 0.00103326f $X=0.216 $Y=0.2025 $X2=0.135 $Y2=0.1355
cc_47 N_5_c_72_p N_Y_c_92_n 0.00328977f $X=0.216 $Y=0.2025 $X2=0.189 $Y2=0.2025
cc_48 N_5_c_64_n N_Y_c_92_n 0.00350506f $X=0.324 $Y=0.2025 $X2=0.189 $Y2=0.2025
cc_49 N_5_c_75_p N_Y_c_92_n 5.59832e-19 $X=0.261 $Y=0.198 $X2=0.189 $Y2=0.2025
cc_50 N_5_c_76_p N_Y_c_92_n 0.00175493f $X=0.2925 $Y=0.198 $X2=0.189 $Y2=0.2025
cc_51 N_5_c_64_n N_Y_c_109_n 0.00374846f $X=0.324 $Y=0.2025 $X2=0 $Y2=0
cc_52 N_5_c_67_n N_Y_c_109_n 3.97701e-19 $X=0.324 $Y=0.198 $X2=0 $Y2=0
cc_53 N_5_c_57_n N_Y_c_87_n 0.00122007f $X=0.108 $Y=0.2025 $X2=0 $Y2=0
cc_54 N_5_c_64_n N_Y_c_95_n 0.00137166f $X=0.324 $Y=0.2025 $X2=0 $Y2=0
cc_55 N_5_c_64_n N_Y_c_101_n 0.0025091f $X=0.324 $Y=0.2025 $X2=0 $Y2=0
cc_56 N_5_c_82_p N_Y_c_101_n 6.95286e-19 $X=0.216 $Y=0.234 $X2=0 $Y2=0
cc_57 N_5_c_76_p N_Y_c_101_n 0.00640856f $X=0.2925 $Y=0.198 $X2=0 $Y2=0
cc_58 N_5_c_67_n N_Y_c_116_n 3.4706e-19 $X=0.324 $Y=0.198 $X2=0 $Y2=0

* END of "./NOR2x1p5_ASAP7_75t_R.pex.sp.NOR2X1P5_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR2x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:43:12 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR2x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR2x2_ASAP7_75t_R.pex.sp.pex"
* File: NOR2x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:43:12 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR2X2_ASAP7_75T_R%B 2 5 8 11 13 16 21 24 27 32 35 36 37 38 39 41 42
+ 43 44 45 46 47 49 50 51 52 53 54 VSS
c73 54 VSS 5.56748e-19 $X=0.459 $Y=0.153
c74 53 VSS 2.64552e-19 $X=0.434 $Y=0.162
c75 52 VSS 0.00120695f $X=0.418 $Y=0.162
c76 51 VSS 0.00127853f $X=0.34 $Y=0.162
c77 50 VSS 2.97889e-19 $X=0.45 $Y=0.162
c78 49 VSS 6.6029e-19 $X=0.331 $Y=0.189
c79 47 VSS 3.12831e-19 $X=0.3005 $Y=0.198
c80 46 VSS 8.46035e-21 $X=0.279 $Y=0.198
c81 45 VSS 3.14008e-19 $X=0.261 $Y=0.198
c82 44 VSS 0.00152288f $X=0.242 $Y=0.198
c83 43 VSS 7.41509e-19 $X=0.218 $Y=0.198
c84 42 VSS 0.0022087f $X=0.322 $Y=0.198
c85 41 VSS 6.6029e-19 $X=0.209 $Y=0.189
c86 39 VSS 2.13186e-19 $X=0.122 $Y=0.162
c87 38 VSS 9.36999e-20 $X=0.109 $Y=0.162
c88 37 VSS 6.87104e-20 $X=0.09 $Y=0.162
c89 36 VSS 0.00248547f $X=0.2 $Y=0.162
c90 32 VSS 0.00126201f $X=0.081 $Y=0.135
c91 24 VSS 0.0718082f $X=0.459 $Y=0.135
c92 16 VSS 0.0623886f $X=0.405 $Y=0.0675
c93 11 VSS 0.00381086f $X=0.135 $Y=0.135
c94 8 VSS 0.0623954f $X=0.135 $Y=0.0675
c95 2 VSS 0.0680685f $X=0.081 $Y=0.135
r96 54 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.153 $X2=0.459 $Y2=0.135
r97 52 53 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.162 $X2=0.434 $Y2=0.162
r98 51 52 5.2963 $w=1.8e-08 $l=7.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.34
+ $Y=0.162 $X2=0.418 $Y2=0.162
r99 50 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.162 $X2=0.459 $Y2=0.153
r100 50 53 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.162 $X2=0.434 $Y2=0.162
r101 48 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.331 $Y=0.171 $X2=0.34 $Y2=0.162
r102 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.331
+ $Y=0.171 $X2=0.331 $Y2=0.189
r103 46 47 1.45988 $w=1.8e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.198 $X2=0.3005 $Y2=0.198
r104 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.198 $X2=0.279 $Y2=0.198
r105 44 45 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.242
+ $Y=0.198 $X2=0.261 $Y2=0.198
r106 43 44 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.218
+ $Y=0.198 $X2=0.242 $Y2=0.198
r107 42 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.322 $Y=0.198 $X2=0.331 $Y2=0.189
r108 42 47 1.45988 $w=1.8e-08 $l=2.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.322
+ $Y=0.198 $X2=0.3005 $Y2=0.198
r109 41 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.209 $Y=0.189 $X2=0.218 $Y2=0.198
r110 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.209
+ $Y=0.171 $X2=0.209 $Y2=0.189
r111 38 39 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.162 $X2=0.122 $Y2=0.162
r112 37 38 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.162 $X2=0.109 $Y2=0.162
r113 36 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.2 $Y=0.162 $X2=0.209 $Y2=0.171
r114 36 39 5.2963 $w=1.8e-08 $l=7.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.2
+ $Y=0.162 $X2=0.122 $Y2=0.162
r115 32 35 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.152
r116 30 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.153 $X2=0.09 $Y2=0.162
r117 30 35 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.153 $X2=0.081 $Y2=0.152
r118 24 56 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r119 24 27 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r120 19 24 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r121 19 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r122 16 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r123 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r124 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r125 2 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r126 2 32 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r127 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
.ends

.subckt PM_NOR2X2_ASAP7_75T_R%A 2 7 10 13 16 19 22 25 27 35 VSS
c39 35 VSS 0.00226955f $X=0.272 $Y=0.136
c40 25 VSS 0.0123218f $X=0.351 $Y=0.1355
c41 22 VSS 0.062303f $X=0.351 $Y=0.0675
c42 16 VSS 0.0643897f $X=0.297 $Y=0.1355
c43 10 VSS 0.0645813f $X=0.243 $Y=0.1355
c44 2 VSS 0.0622987f $X=0.189 $Y=0.0675
r45 32 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.27 $Y=0.135 $X2=0.27
+ $Y2=0.135
r46 25 27 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.1355 $X2=0.351 $Y2=0.2025
r47 22 25 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.1355
r48 16 25 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.1355 $X2=0.351 $Y2=0.1355
r49 16 32 23.4783 $w=2.3e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.1355 $X2=0.27 $Y2=0.1355
r50 16 19 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.1355 $X2=0.297 $Y2=0.2025
r51 10 32 23.4783 $w=2.3e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.1355 $X2=0.27 $Y2=0.1355
r52 10 13 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1355 $X2=0.243 $Y2=0.2025
r53 5 10 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.1355 $X2=0.243 $Y2=0.1355
r54 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1355 $X2=0.189 $Y2=0.2025
r55 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.1355
.ends

.subckt PM_NOR2X2_ASAP7_75T_R%5 1 4 6 7 10 11 12 15 16 17 20 21 24 33 34 38 39
+ 43 44 46 48 49 VSS
c40 49 VSS 0.00261806f $X=0.452 $Y=0.234
c41 48 VSS 0.00456882f $X=0.418 $Y=0.234
c42 46 VSS 0.00500247f $X=0.486 $Y=0.234
c43 44 VSS 0.0015425f $X=0.359 $Y=0.234
c44 43 VSS 0.0107037f $X=0.34 $Y=0.234
c45 39 VSS 0.00520575f $X=0.235 $Y=0.234
c46 38 VSS 0.0044884f $X=0.2 $Y=0.234
c47 34 VSS 0.00162279f $X=0.142 $Y=0.234
c48 33 VSS 0.00762831f $X=0.122 $Y=0.234
c49 24 VSS 0.00262643f $X=0.484 $Y=0.2025
c50 20 VSS 0.00713099f $X=0.378 $Y=0.2025
c51 16 VSS 7.6997e-19 $X=0.395 $Y=0.2025
c52 15 VSS 0.0100322f $X=0.27 $Y=0.2025
c53 11 VSS 6.26354e-19 $X=0.287 $Y=0.2025
c54 10 VSS 0.00713099f $X=0.162 $Y=0.2025
c55 6 VSS 7.6997e-19 $X=0.179 $Y=0.2025
c56 4 VSS 0.00228092f $X=0.056 $Y=0.2025
c57 1 VSS 3.4551e-19 $X=0.071 $Y=0.2025
r58 48 49 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.234 $X2=0.452 $Y2=0.234
r59 46 49 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.452 $Y2=0.234
r60 43 44 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.34
+ $Y=0.234 $X2=0.359 $Y2=0.234
r61 41 48 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.418 $Y2=0.234
r62 41 44 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.359 $Y2=0.234
r63 38 39 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.2
+ $Y=0.234 $X2=0.235 $Y2=0.234
r64 36 43 4.75309 $w=1.8e-08 $l=7e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.34 $Y2=0.234
r65 36 39 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.235 $Y2=0.234
r66 33 34 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.122
+ $Y=0.234 $X2=0.142 $Y2=0.234
r67 31 38 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.2 $Y2=0.234
r68 31 34 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.142 $Y2=0.234
r69 27 33 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.122 $Y2=0.234
r70 24 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r71 21 24 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.484 $Y2=0.2025
r72 20 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r73 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r74 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r75 15 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r76 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r77 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r78 10 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r79 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r80 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r81 4 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r82 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
.ends

.subckt PM_NOR2X2_ASAP7_75T_R%Y 1 6 11 16 21 22 25 26 27 30 34 39 41 44 45 46 49
+ 50 51 52 53 56 57 58 61 64 71 72 76 VSS
c62 80 VSS 3.80356e-19 $X=0.513 $Y=0.18
c63 78 VSS 0.00130599f $X=0.513 $Y=0.093
c64 77 VSS 9.03568e-19 $X=0.513 $Y=0.063
c65 76 VSS 0.00332325f $X=0.514 $Y=0.145
c66 74 VSS 3.59225e-19 $X=0.513 $Y=0.189
c67 72 VSS 4.78169e-19 $X=0.5 $Y=0.198
c68 71 VSS 8.46035e-21 $X=0.468 $Y=0.198
c69 66 VSS 0.00220485f $X=0.504 $Y=0.198
c70 64 VSS 4.78169e-19 $X=0.072 $Y=0.198
c71 63 VSS 2.76758e-19 $X=0.04 $Y=0.198
c72 61 VSS 8.46035e-21 $X=0.108 $Y=0.198
c73 59 VSS 0.00192809f $X=0.036 $Y=0.198
c74 58 VSS 0.00146362f $X=0.468 $Y=0.036
c75 57 VSS 0.0137555f $X=0.45 $Y=0.036
c76 56 VSS 0.0064565f $X=0.432 $Y=0.036
c77 53 VSS 0.00395819f $X=0.322 $Y=0.036
c78 52 VSS 0.00324847f $X=0.279 $Y=0.036
c79 51 VSS 0.00226617f $X=0.242 $Y=0.036
c80 50 VSS 0.00608839f $X=0.218 $Y=0.036
c81 49 VSS 0.0071986f $X=0.324 $Y=0.036
c82 46 VSS 0.00606865f $X=0.1625 $Y=0.036
c83 45 VSS 0.00142953f $X=0.109 $Y=0.036
c84 44 VSS 0.0071979f $X=0.216 $Y=0.036
c85 41 VSS 0.00146362f $X=0.09 $Y=0.036
c86 40 VSS 0.00346625f $X=0.072 $Y=0.036
c87 39 VSS 0.0069473f $X=0.108 $Y=0.036
c88 36 VSS 0.00350046f $X=0.036 $Y=0.036
c89 35 VSS 0.00696671f $X=0.504 $Y=0.036
c90 34 VSS 0.00462133f $X=0.027 $Y=0.171
c91 33 VSS 9.03568e-19 $X=0.027 $Y=0.063
c92 32 VSS 7.39581e-19 $X=0.027 $Y=0.189
c93 30 VSS 0.00283195f $X=0.432 $Y=0.2025
c94 26 VSS 6.19444e-19 $X=0.449 $Y=0.2025
c95 25 VSS 0.00283195f $X=0.108 $Y=0.2025
c96 21 VSS 6.18143e-19 $X=0.125 $Y=0.2025
c97 19 VSS 4.59792e-19 $X=0.43 $Y=0.0675
c98 11 VSS 4.6121e-19 $X=0.341 $Y=0.0675
c99 9 VSS 4.6121e-19 $X=0.214 $Y=0.0675
c100 1 VSS 4.59792e-19 $X=0.125 $Y=0.0675
r101 79 80 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.171 $X2=0.513 $Y2=0.18
r102 77 78 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.063 $X2=0.513 $Y2=0.093
r103 76 79 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.145 $X2=0.513 $Y2=0.171
r104 76 78 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.145 $X2=0.513 $Y2=0.093
r105 74 80 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.513 $Y2=0.18
r106 73 77 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.063
r107 71 72 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.198 $X2=0.5 $Y2=0.198
r108 68 71 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.468 $Y2=0.198
r109 66 74 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.198 $X2=0.513 $Y2=0.189
r110 66 72 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.198 $X2=0.5 $Y2=0.198
r111 63 64 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.198 $X2=0.072 $Y2=0.198
r112 61 64 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.198 $X2=0.072 $Y2=0.198
r113 59 63 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.198 $X2=0.04 $Y2=0.198
r114 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r115 55 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r116 55 56 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r117 52 53 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.036 $X2=0.322 $Y2=0.036
r118 51 52 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.242
+ $Y=0.036 $X2=0.279 $Y2=0.036
r119 50 51 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.218
+ $Y=0.036 $X2=0.242 $Y2=0.036
r120 48 55 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r121 48 53 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.322 $Y2=0.036
r122 48 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r123 45 46 3.63272 $w=1.8e-08 $l=5.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.036 $X2=0.1625 $Y2=0.036
r124 43 50 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.218 $Y2=0.036
r125 43 46 3.63272 $w=1.8e-08 $l=5.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.1625 $Y2=0.036
r126 43 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r127 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r128 38 45 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.109 $Y2=0.036
r129 38 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.09 $Y2=0.036
r130 38 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r131 36 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.072 $Y2=0.036
r132 35 73 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.036 $X2=0.513 $Y2=0.045
r133 35 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.468 $Y2=0.036
r134 33 34 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.063 $X2=0.027 $Y2=0.171
r135 32 59 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.189 $X2=0.036 $Y2=0.198
r136 32 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.027 $Y2=0.171
r137 31 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r138 31 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.063
r139 30 68 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198
+ $X2=0.432 $Y2=0.198
r140 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r141 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r142 25 61 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.198
+ $X2=0.108 $Y2=0.198
r143 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r144 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r145 19 56 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r146 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.43 $Y2=0.0675
r147 14 49 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r148 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.326 $Y2=0.0675
r149 9 44 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r150 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.214 $Y2=0.0675
r151 4 39 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r152 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.11 $Y2=0.0675
.ends


* END of "./NOR2x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR2x2_ASAP7_75t_R  VSS VDD B A Y
* 
* Y	Y
* A	A
* B	B
M0 VSS N_B_M0_g N_Y_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M1 N_Y_M1_d N_A_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M2 N_Y_M2_d N_A_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M3 VSS N_B_M3_g N_Y_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M4 N_Y_M4_d N_B_M4_g N_5_M4_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 N_Y_M5_d N_B_M5_g N_5_M5_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 VDD N_A_M6_g N_5_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M7 VDD N_A_M7_g N_5_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M8 VDD N_A_M8_g N_5_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
M9 VDD N_A_M9_g N_5_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.162
M10 N_Y_M10_d N_B_M10_g N_5_M10_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M11 N_Y_M11_d N_B_M11_g N_5_M11_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "NOR2x2_ASAP7_75t_R.pex.sp.NOR2X2_ASAP7_75T_R.pxi"
* BEGIN of "./NOR2x2_ASAP7_75t_R.pex.sp.NOR2X2_ASAP7_75T_R.pxi"
* File: NOR2x2_ASAP7_75t_R.pex.sp.NOR2X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:43:12 2017
* 
x_PM_NOR2X2_ASAP7_75T_R%B N_B_c_1_p N_B_M4_g N_B_M0_g N_B_c_11_p N_B_M5_g
+ N_B_M3_g N_B_M10_g N_B_c_9_p N_B_M11_g N_B_c_17_p B N_B_c_3_p N_B_c_22_p
+ N_B_c_42_p N_B_c_43_p N_B_c_24_p N_B_c_70_p N_B_c_34_p N_B_c_14_p N_B_c_5_p
+ N_B_c_19_p N_B_c_7_p N_B_c_28_p N_B_c_30_p N_B_c_16_p N_B_c_10_p N_B_c_47_p
+ N_B_c_21_p VSS PM_NOR2X2_ASAP7_75T_R%B
x_PM_NOR2X2_ASAP7_75T_R%A N_A_M1_g N_A_M6_g N_A_c_77_n N_A_M7_g N_A_c_79_n
+ N_A_M8_g N_A_M2_g N_A_c_84_n N_A_M9_g A VSS PM_NOR2X2_ASAP7_75T_R%A
x_PM_NOR2X2_ASAP7_75T_R%5 N_5_M4_s N_5_c_113_n N_5_M6_s N_5_M5_s N_5_c_114_n
+ N_5_M8_s N_5_M7_s N_5_c_116_n N_5_M10_s N_5_M9_s N_5_c_119_n N_5_M11_s
+ N_5_c_121_n N_5_c_122_n N_5_c_123_n N_5_c_133_n N_5_c_125_n N_5_c_126_n
+ N_5_c_127_n N_5_c_128_n N_5_c_129_n N_5_c_142_p VSS PM_NOR2X2_ASAP7_75T_R%5
x_PM_NOR2X2_ASAP7_75T_R%Y N_Y_M0_s N_Y_M1_d N_Y_M2_d N_Y_M3_s N_Y_M5_d N_Y_M4_d
+ N_Y_c_155_n N_Y_M11_d N_Y_M10_d N_Y_c_159_n N_Y_c_162_n N_Y_c_164_n
+ N_Y_c_166_n N_Y_c_188_n N_Y_c_168_n N_Y_c_169_n N_Y_c_190_n N_Y_c_172_n
+ N_Y_c_194_n N_Y_c_195_n N_Y_c_196_n N_Y_c_173_n N_Y_c_175_n N_Y_c_178_n
+ N_Y_c_180_n N_Y_c_207_n N_Y_c_183_n N_Y_c_212_n Y VSS PM_NOR2X2_ASAP7_75T_R%Y
cc_1 N_B_c_1_p N_A_M1_g 2.66145e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_2 N_B_M0_g N_A_M1_g 0.0032073f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_B_c_3_p N_A_M1_g 4.19577e-19 $X=0.2 $Y=0.162 $X2=0.189 $Y2=0.0675
cc_4 N_B_M0_g N_A_c_77_n 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.1355
cc_5 N_B_c_5_p N_A_c_77_n 2.1804e-19 $X=0.261 $Y=0.198 $X2=0.243 $Y2=0.1355
cc_6 N_B_M3_g N_A_c_79_n 2.31381e-19 $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.1355
cc_7 N_B_c_7_p N_A_c_79_n 2.66132e-19 $X=0.3005 $Y=0.198 $X2=0.297 $Y2=0.1355
cc_8 N_B_M3_g N_A_M2_g 0.0032073f $X=0.405 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_9 N_B_c_9_p N_A_M2_g 2.66145e-19 $X=0.459 $Y=0.135 $X2=0.351 $Y2=0.0675
cc_10 N_B_c_10_p N_A_M2_g 4.19577e-19 $X=0.418 $Y=0.162 $X2=0.351 $Y2=0.0675
cc_11 N_B_c_11_p N_A_c_84_n 0.00227362f $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.1355
cc_12 N_B_c_9_p N_A_c_84_n 0.00227362f $X=0.459 $Y=0.135 $X2=0.351 $Y2=0.1355
cc_13 N_B_c_3_p N_A_c_84_n 0.00124067f $X=0.2 $Y=0.162 $X2=0.351 $Y2=0.1355
cc_14 N_B_c_14_p N_A_c_84_n 8.12001e-19 $X=0.242 $Y=0.198 $X2=0.351 $Y2=0.1355
cc_15 N_B_c_7_p N_A_c_84_n 8.41977e-19 $X=0.3005 $Y=0.198 $X2=0.351 $Y2=0.1355
cc_16 N_B_c_16_p N_A_c_84_n 0.00124067f $X=0.34 $Y=0.162 $X2=0.351 $Y2=0.1355
cc_17 N_B_c_17_p A 5.12949e-19 $X=0.081 $Y=0.135 $X2=0.272 $Y2=0.136
cc_18 N_B_c_3_p A 4.78502e-19 $X=0.2 $Y=0.162 $X2=0.272 $Y2=0.136
cc_19 N_B_c_19_p A 0.00101457f $X=0.279 $Y=0.198 $X2=0.272 $Y2=0.136
cc_20 N_B_c_16_p A 6.38258e-19 $X=0.34 $Y=0.162 $X2=0.272 $Y2=0.136
cc_21 N_B_c_21_p A 4.34071e-19 $X=0.459 $Y=0.153 $X2=0.272 $Y2=0.136
cc_22 N_B_c_22_p N_5_c_113_n 2.78572e-19 $X=0.09 $Y=0.162 $X2=0.189 $Y2=0.1355
cc_23 N_B_c_3_p N_5_c_114_n 0.00201076f $X=0.2 $Y=0.162 $X2=0.243 $Y2=0.1355
cc_24 N_B_c_24_p N_5_c_114_n 7.67394e-19 $X=0.209 $Y=0.189 $X2=0.243 $Y2=0.1355
cc_25 N_B_c_5_p N_5_c_116_n 5.61323e-19 $X=0.261 $Y=0.198 $X2=0.297 $Y2=0.1355
cc_26 N_B_c_19_p N_5_c_116_n 0.00124096f $X=0.279 $Y=0.198 $X2=0.297 $Y2=0.1355
cc_27 N_B_c_7_p N_5_c_116_n 5.58359e-19 $X=0.3005 $Y=0.198 $X2=0.297 $Y2=0.1355
cc_28 N_B_c_28_p N_5_c_119_n 7.67394e-19 $X=0.331 $Y=0.189 $X2=0 $Y2=0
cc_29 N_B_c_10_p N_5_c_119_n 0.00201076f $X=0.418 $Y=0.162 $X2=0 $Y2=0
cc_30 N_B_c_30_p N_5_c_121_n 2.78572e-19 $X=0.45 $Y=0.162 $X2=0.351 $Y2=0.1355
cc_31 N_B_c_1_p N_5_c_122_n 2.38303e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_32 N_B_M0_g N_5_c_123_n 3.24635e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_33 N_B_c_3_p N_5_c_123_n 0.00230303f $X=0.2 $Y=0.162 $X2=0 $Y2=0
cc_34 N_B_c_34_p N_5_c_125_n 0.0059448f $X=0.218 $Y=0.198 $X2=0 $Y2=0
cc_35 N_B_c_19_p N_5_c_126_n 0.0059448f $X=0.279 $Y=0.198 $X2=0.27 $Y2=0.1355
cc_36 N_B_c_10_p N_5_c_127_n 0.00230302f $X=0.418 $Y=0.162 $X2=0.297 $Y2=0.1355
cc_37 N_B_c_9_p N_5_c_128_n 2.08515e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_38 N_B_M3_g N_5_c_129_n 3.81924e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_B_c_17_p N_Y_M0_s 2.0764e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_40 N_B_c_11_p N_Y_M5_d 3.70143e-19 $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.0675
cc_41 N_B_c_11_p N_Y_c_155_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.1355
cc_42 N_B_c_42_p N_Y_c_155_n 7.62637e-19 $X=0.109 $Y=0.162 $X2=0.351 $Y2=0.1355
cc_43 N_B_c_43_p N_Y_c_155_n 8.29904e-19 $X=0.122 $Y=0.162 $X2=0.351 $Y2=0.1355
cc_44 N_B_c_9_p N_Y_M11_d 3.70143e-19 $X=0.459 $Y=0.135 $X2=0.351 $Y2=0.2025
cc_45 N_B_c_9_p N_Y_c_159_n 8.0006e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_46 N_B_c_30_p N_Y_c_159_n 6.01614e-19 $X=0.45 $Y=0.162 $X2=0 $Y2=0
cc_47 N_B_c_47_p N_Y_c_159_n 9.90927e-19 $X=0.434 $Y=0.162 $X2=0 $Y2=0
cc_48 N_B_c_11_p N_Y_c_162_n 3.39417e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_49 N_B_c_17_p N_Y_c_162_n 0.00519692f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_50 N_B_c_11_p N_Y_c_164_n 8.00061e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_51 N_B_c_17_p N_Y_c_164_n 0.00261434f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_52 N_B_c_1_p N_Y_c_166_n 2.38303e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_53 N_B_c_17_p N_Y_c_166_n 0.00371886f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_54 N_B_c_42_p N_Y_c_168_n 4.64167e-19 $X=0.109 $Y=0.162 $X2=0.351 $Y2=0.1355
cc_55 N_B_M0_g N_Y_c_169_n 4.52603e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_56 N_B_c_11_p N_Y_c_169_n 3.30932e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_57 N_B_c_43_p N_Y_c_169_n 4.64167e-19 $X=0.122 $Y=0.162 $X2=0 $Y2=0
cc_58 N_B_c_3_p N_Y_c_172_n 4.64167e-19 $X=0.2 $Y=0.162 $X2=0 $Y2=0
cc_59 N_B_c_9_p N_Y_c_173_n 8.0006e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_60 N_B_c_21_p N_Y_c_173_n 5.27536e-19 $X=0.459 $Y=0.153 $X2=0 $Y2=0
cc_61 N_B_M3_g N_Y_c_175_n 4.52603e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_62 N_B_c_9_p N_Y_c_175_n 4.74833e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_63 N_B_c_16_p N_Y_c_175_n 0.00160573f $X=0.34 $Y=0.162 $X2=0 $Y2=0
cc_64 N_B_c_9_p N_Y_c_178_n 3.30638e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_65 N_B_c_21_p N_Y_c_178_n 6.86694e-19 $X=0.459 $Y=0.153 $X2=0 $Y2=0
cc_66 N_B_c_1_p N_Y_c_180_n 2.52885e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_67 N_B_c_22_p N_Y_c_180_n 0.00408818f $X=0.09 $Y=0.162 $X2=0 $Y2=0
cc_68 N_B_c_34_p N_Y_c_180_n 2.95701e-19 $X=0.218 $Y=0.198 $X2=0 $Y2=0
cc_69 N_B_c_9_p N_Y_c_183_n 2.52885e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_70 N_B_c_70_p N_Y_c_183_n 2.95701e-19 $X=0.322 $Y=0.198 $X2=0 $Y2=0
cc_71 N_B_c_47_p N_Y_c_183_n 0.00407975f $X=0.434 $Y=0.162 $X2=0 $Y2=0
cc_72 N_B_c_9_p Y 3.39417e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_73 N_B_c_21_p Y 0.00372982f $X=0.459 $Y=0.153 $X2=0 $Y2=0
cc_74 N_A_c_84_n N_5_M8_s 3.89915e-19 $X=0.351 $Y=0.1355 $X2=0.135 $Y2=0.135
cc_75 N_A_c_84_n N_5_c_116_n 0.00227427f $X=0.351 $Y=0.1355 $X2=0.405 $Y2=0.0675
cc_76 A N_5_c_116_n 0.0438982f $X=0.272 $Y=0.136 $X2=0.405 $Y2=0.0675
cc_77 N_A_M1_g N_5_c_133_n 3.80935e-19 $X=0.189 $Y=0.0675 $X2=0.109 $Y2=0.162
cc_78 N_A_c_77_n N_5_c_126_n 2.34767e-19 $X=0.243 $Y=0.1355 $X2=0.218 $Y2=0.198
cc_79 N_A_c_79_n N_5_c_126_n 2.64526e-19 $X=0.297 $Y=0.1355 $X2=0.218 $Y2=0.198
cc_80 N_A_M2_g N_5_c_127_n 3.42841e-19 $X=0.351 $Y=0.0675 $X2=0.242 $Y2=0.198
cc_81 N_A_c_84_n N_Y_c_188_n 8.01479e-19 $X=0.351 $Y=0.1355 $X2=0.242 $Y2=0.198
cc_82 A N_Y_c_188_n 0.0010607f $X=0.272 $Y=0.136 $X2=0.242 $Y2=0.198
cc_83 N_A_c_84_n N_Y_c_190_n 8.01479e-19 $X=0.351 $Y=0.1355 $X2=0.331 $Y2=0.189
cc_84 A N_Y_c_190_n 0.00105555f $X=0.272 $Y=0.136 $X2=0.331 $Y2=0.189
cc_85 N_A_M1_g N_Y_c_172_n 4.52603e-19 $X=0.189 $Y=0.0675 $X2=0.45 $Y2=0.162
cc_86 N_A_c_84_n N_Y_c_172_n 5.47817e-19 $X=0.351 $Y=0.1355 $X2=0.45 $Y2=0.162
cc_87 N_A_c_77_n N_Y_c_194_n 2.08223e-19 $X=0.243 $Y=0.1355 $X2=0.34 $Y2=0.162
cc_88 A N_Y_c_195_n 0.0035884f $X=0.272 $Y=0.136 $X2=0.418 $Y2=0.162
cc_89 N_A_c_79_n N_Y_c_196_n 4.62717e-19 $X=0.297 $Y=0.1355 $X2=0.434 $Y2=0.162
cc_90 N_A_c_84_n N_Y_c_196_n 7.12009e-19 $X=0.351 $Y=0.1355 $X2=0.434 $Y2=0.162
cc_91 N_A_M2_g N_Y_c_175_n 4.52603e-19 $X=0.351 $Y=0.0675 $X2=0.459 $Y2=0.135
cc_92 N_5_c_113_n N_Y_c_155_n 0.00384463f $X=0.056 $Y=0.2025 $X2=0 $Y2=0
cc_93 N_5_c_114_n N_Y_c_155_n 0.00363853f $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_94 N_5_c_122_n N_Y_c_155_n 0.0025091f $X=0.122 $Y=0.234 $X2=0 $Y2=0
cc_95 N_5_c_119_n N_Y_c_159_n 0.00363853f $X=0.378 $Y=0.2025 $X2=0.081 $Y2=0.153
cc_96 N_5_c_121_n N_Y_c_159_n 0.00384463f $X=0.484 $Y=0.2025 $X2=0.081 $Y2=0.153
cc_97 N_5_c_142_p N_Y_c_159_n 0.0025091f $X=0.452 $Y=0.234 $X2=0.081 $Y2=0.153
cc_98 N_5_c_113_n N_Y_c_162_n 2.86097e-19 $X=0.056 $Y=0.2025 $X2=0.081 $Y2=0.152
cc_99 N_5_c_114_n N_Y_c_180_n 4.45525e-19 $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_100 N_5_M4_s N_Y_c_207_n 2.53396e-19 $X=0.071 $Y=0.2025 $X2=0.405 $Y2=0.135
cc_101 N_5_c_113_n N_Y_c_207_n 0.00263302f $X=0.056 $Y=0.2025 $X2=0.405
+ $Y2=0.135
cc_102 N_5_c_122_n N_Y_c_207_n 0.00709175f $X=0.122 $Y=0.234 $X2=0.405 $Y2=0.135
cc_103 N_5_c_119_n N_Y_c_183_n 4.45525e-19 $X=0.378 $Y=0.2025 $X2=0 $Y2=0
cc_104 N_5_c_142_p N_Y_c_183_n 0.00354594f $X=0.452 $Y=0.234 $X2=0 $Y2=0
cc_105 N_5_c_121_n N_Y_c_212_n 0.00288641f $X=0.484 $Y=0.2025 $X2=0 $Y2=0
cc_106 N_5_c_128_n N_Y_c_212_n 0.00354594f $X=0.486 $Y=0.234 $X2=0 $Y2=0
cc_107 N_5_c_121_n Y 2.85653e-19 $X=0.484 $Y=0.2025 $X2=0 $Y2=0

* END of "./NOR2x2_ASAP7_75t_R.pex.sp.NOR2X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR2xp33_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:43:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR2xp33_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR2xp33_ASAP7_75t_R.pex.sp.pex"
* File: NOR2xp33_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:43:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR2XP33_ASAP7_75T_R%A 2 5 7 19 VSS
c5 19 VSS 0.0263471f $X=0.06 $Y=0.135
c6 5 VSS 0.00582264f $X=0.081 $Y=0.135
c7 2 VSS 0.0643819f $X=0.081 $Y=0.0405
r8 19 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r9 5 23 18.8889 $w=1.8e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r10 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r11 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0405 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NOR2XP33_ASAP7_75T_R%B 2 5 7 12 VSS
c10 12 VSS 0.00423739f $X=0.135 $Y=0.135
c11 5 VSS 0.00156845f $X=0.135 $Y=0.135
c12 2 VSS 0.0638285f $X=0.135 $Y=0.0405
r13 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r14 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r15 2 5 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0405 $X2=0.135 $Y2=0.135
.ends

.subckt PM_NOR2XP33_ASAP7_75T_R%Y 1 2 6 9 13 18 22 30 32 VSS
c8 34 VSS 4.55454e-19 $X=0.189 $Y=0.216
c9 32 VSS 0.00158366f $X=0.189 $Y=0.099
c10 31 VSS 8.85605e-19 $X=0.189 $Y=0.063
c11 30 VSS 0.00483084f $X=0.19 $Y=0.135
c12 28 VSS 4.30151e-19 $X=0.189 $Y=0.225
c13 22 VSS 0.00166239f $X=0.162 $Y=0.234
c14 20 VSS 0.00607663f $X=0.18 $Y=0.234
c15 19 VSS 0.00303662f $X=0.162 $Y=0.036
c16 18 VSS 0.00288209f $X=0.144 $Y=0.036
c17 13 VSS 0.0023094f $X=0.108 $Y=0.036
c18 11 VSS 0.00621531f $X=0.18 $Y=0.036
c19 9 VSS 0.0041197f $X=0.16 $Y=0.216
c20 5 VSS 0.00562504f $X=0.108 $Y=0.0405
c21 1 VSS 6.15566e-19 $X=0.125 $Y=0.0405
r22 33 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.207 $X2=0.189 $Y2=0.216
r23 31 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.063 $X2=0.189 $Y2=0.099
r24 30 33 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.207
r25 30 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.099
r26 28 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.216
r27 27 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.045 $X2=0.189 $Y2=0.063
r28 20 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.234 $X2=0.189 $Y2=0.225
r29 20 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.162 $Y2=0.234
r30 18 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.162 $Y2=0.036
r31 13 18 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.144 $Y2=0.036
r32 11 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.036 $X2=0.189 $Y2=0.045
r33 11 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.162 $Y2=0.036
r34 9 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r35 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.145
+ $Y=0.216 $X2=0.16 $Y2=0.216
r36 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r37 2 5 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0405 $X2=0.108 $Y2=0.0405
r38 1 5 25.1852 $w=2.7e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0405 $X2=0.108 $Y2=0.0405
.ends

.subckt PM_NOR2XP33_ASAP7_75T_R%6 1 2 VSS
c1 1 VSS 0.00221012f $X=0.125 $Y=0.216
r2 1 2 25.1852 $w=5.4e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.216 $X2=0.091 $Y2=0.216
.ends


* END of "./NOR2xp33_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR2xp33_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_RVT L=2e-08 W=2.7e-08 NFIN=1 $X=0.071 $Y=0.027
M1 VSS N_B_M1_g N_Y_M1_s VSS NMOS_RVT L=2e-08 W=2.7e-08 NFIN=1 $X=0.125 $Y=0.027
M2 N_6_M2_d N_A_M2_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M3 N_Y_M3_d N_B_M3_g N_6_M3_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
*
* 
* .include "NOR2xp33_ASAP7_75t_R.pex.sp.NOR2XP33_ASAP7_75T_R.pxi"
* BEGIN of "./NOR2xp33_ASAP7_75t_R.pex.sp.NOR2XP33_ASAP7_75T_R.pxi"
* File: NOR2xp33_ASAP7_75t_R.pex.sp.NOR2XP33_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:43:34 2017
* 
x_PM_NOR2XP33_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M2_g A VSS
+ PM_NOR2XP33_ASAP7_75T_R%A
x_PM_NOR2XP33_ASAP7_75T_R%B N_B_M1_g N_B_c_7_n N_B_M3_g B VSS
+ PM_NOR2XP33_ASAP7_75T_R%B
x_PM_NOR2XP33_ASAP7_75T_R%Y N_Y_M1_s N_Y_M0_d N_Y_M3_d N_Y_c_18_n N_Y_c_16_n
+ N_Y_c_19_n N_Y_c_17_n Y N_Y_c_23_n VSS PM_NOR2XP33_ASAP7_75T_R%Y
x_PM_NOR2XP33_ASAP7_75T_R%6 N_6_M3_s N_6_M2_d VSS PM_NOR2XP33_ASAP7_75T_R%6
cc_1 N_A_M0_g N_B_M1_g 0.00344695f $X=0.081 $Y=0.0405 $X2=0.135 $Y2=0.0405
cc_2 N_A_c_2_p N_B_c_7_n 8.71247e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A B 0.0027917f $X=0.06 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 A N_Y_c_16_n 5.24213e-19 $X=0.06 $Y=0.135 $X2=0 $Y2=0
cc_5 A N_Y_c_17_n 2.61367e-19 $X=0.06 $Y=0.135 $X2=0 $Y2=0
cc_6 B N_Y_c_18_n 6.42527e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_7 N_B_M1_g N_Y_c_19_n 2.25474e-19 $X=0.135 $Y=0.0405 $X2=0 $Y2=0
cc_8 B N_Y_c_19_n 0.0036051f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_9 N_B_M1_g N_Y_c_17_n 3.14377e-19 $X=0.135 $Y=0.0405 $X2=0.064 $Y2=0.135
cc_10 B Y 0.00340691f $X=0.135 $Y=0.135 $X2=0.064 $Y2=0.135
cc_11 B N_Y_c_23_n 0.00340691f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_12 B N_6_M3_s 2.75518e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.0405

* END of "./NOR2xp33_ASAP7_75t_R.pex.sp.NOR2XP33_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR2xp67_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:43:57 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR2xp67_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR2xp67_ASAP7_75t_R.pex.sp.pex"
* File: NOR2xp67_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:43:57 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR2XP67_ASAP7_75T_R%A 2 7 10 13 23 VSS
c12 23 VSS 0.0198655f $X=0.081 $Y=0.13
c13 10 VSS 0.0708673f $X=0.135 $Y=0.136
c14 2 VSS 0.067081f $X=0.081 $Y=0.054
r15 10 13 299.72 $w=2e-08 $l=8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.136 $X2=0.135 $Y2=0.216
r16 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.136 $X2=0.135 $Y2=0.136
r17 5 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.136 $X2=0.081
+ $Y2=0.136
r18 5 7 299.72 $w=2e-08 $l=8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.136 $X2=0.081 $Y2=0.216
r19 2 5 307.213 $w=2e-08 $l=8.2e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.136
.ends

.subckt PM_NOR2XP67_ASAP7_75T_R%B 2 7 10 13 23 VSS
c22 23 VSS 0.00635012f $X=0.243 $Y=0.134
c23 10 VSS 0.0738524f $X=0.243 $Y=0.136
c24 2 VSS 0.0631829f $X=0.189 $Y=0.054
r25 10 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r26 10 13 299.72 $w=2e-08 $l=8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.136 $X2=0.243 $Y2=0.216
r27 5 10 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.136 $X2=0.243 $Y2=0.136
r28 5 7 299.72 $w=2e-08 $l=8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.136 $X2=0.189 $Y2=0.216
r29 2 5 307.213 $w=2e-08 $l=8.2e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.136
.ends

.subckt PM_NOR2XP67_ASAP7_75T_R%5 1 4 6 7 10 11 14 17 25 27 28 30 32 33 VSS
c20 33 VSS 0.00261791f $X=0.236 $Y=0.234
c21 32 VSS 0.00398061f $X=0.202 $Y=0.234
c22 30 VSS 0.00495854f $X=0.27 $Y=0.234
c23 28 VSS 7.47399e-19 $X=0.153 $Y=0.234
c24 27 VSS 0.00420751f $X=0.144 $Y=0.234
c25 26 VSS 0.00242309f $X=0.107 $Y=0.234
c26 25 VSS 0.00361761f $X=0.095 $Y=0.234
c27 17 VSS 0.00190391f $X=0.054 $Y=0.234
c28 14 VSS 0.00248344f $X=0.268 $Y=0.216
c29 10 VSS 0.00500461f $X=0.162 $Y=0.216
c30 6 VSS 5.3314e-19 $X=0.179 $Y=0.216
c31 4 VSS 0.00605643f $X=0.056 $Y=0.216
c32 1 VSS 2.6657e-19 $X=0.071 $Y=0.216
r33 32 33 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.234 $X2=0.236 $Y2=0.234
r34 30 33 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.236 $Y2=0.234
r35 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.153 $Y2=0.234
r36 26 27 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.234 $X2=0.144 $Y2=0.234
r37 25 26 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.234 $X2=0.107 $Y2=0.234
r38 23 32 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.202 $Y2=0.234
r39 23 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.153 $Y2=0.234
r40 17 25 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.095 $Y2=0.234
r41 14 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r42 11 14 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.216 $X2=0.268 $Y2=0.216
r43 10 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r44 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.162 $Y2=0.216
r45 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.216 $X2=0.162 $Y2=0.216
r46 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r47 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.216 $X2=0.056 $Y2=0.216
.ends

.subckt PM_NOR2XP67_ASAP7_75T_R%Y 1 6 9 11 12 15 21 22 28 29 33 36 37 VSS
c20 37 VSS 7.46755e-19 $X=0.297 $Y=0.144
c21 36 VSS 0.00266718f $X=0.297 $Y=0.126
c22 35 VSS 0.00111622f $X=0.297 $Y=0.081
c23 34 VSS 0.00104959f $X=0.297 $Y=0.063
c24 33 VSS 0.00249264f $X=0.296 $Y=0.164
c25 29 VSS 3.03827e-19 $X=0.284 $Y=0.198
c26 28 VSS 1.1404e-19 $X=0.257 $Y=0.198
c27 23 VSS 0.00215853f $X=0.288 $Y=0.198
c28 22 VSS 0.010489f $X=0.257 $Y=0.036
c29 21 VSS 0.00199353f $X=0.163 $Y=0.036
c30 16 VSS 0.00694576f $X=0.288 $Y=0.036
c31 15 VSS 0.00324684f $X=0.216 $Y=0.216
c32 11 VSS 5.65575e-19 $X=0.233 $Y=0.216
c33 9 VSS 0.0241392f $X=0.164 $Y=0.054
c34 6 VSS 2.6657e-19 $X=0.179 $Y=0.054
c35 4 VSS 3.19801e-19 $X=0.106 $Y=0.054
r36 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.144
r37 35 36 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.081 $X2=0.297 $Y2=0.126
r38 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.063 $X2=0.297 $Y2=0.081
r39 33 37 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.164 $X2=0.297 $Y2=0.144
r40 31 33 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.164
r41 30 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.063
r42 28 29 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.257
+ $Y=0.198 $X2=0.284 $Y2=0.198
r43 25 28 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.257 $Y2=0.198
r44 23 31 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.198 $X2=0.297 $Y2=0.189
r45 23 29 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.284 $Y2=0.198
r46 21 22 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.163
+ $Y=0.036 $X2=0.257 $Y2=0.036
r47 18 21 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.163 $Y2=0.036
r48 16 30 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r49 16 22 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.257 $Y2=0.036
r50 15 25 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r51 12 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.216 $X2=0.216 $Y2=0.216
r52 11 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.216 $X2=0.216 $Y2=0.216
r53 9 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r54 6 9 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.054 $X2=0.164 $Y2=0.054
r55 4 9 21.4815 $w=5.4e-08 $l=5.6e-08 $layer=LISD $thickness=2.8e-08 $X=0.106
+ $Y=0.054 $X2=0.162 $Y2=0.054
r56 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.054 $X2=0.106 $Y2=0.054
.ends


* END of "./NOR2xp67_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR2xp67_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 VSS N_B_M1_g N_Y_M1_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M2 VDD N_A_M2_g N_5_M2_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M3 VDD N_A_M3_g N_5_M3_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
M4 N_Y_M4_d N_B_M4_g N_5_M4_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M5 N_Y_M5_d N_B_M5_g N_5_M5_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
*
* 
* .include "NOR2xp67_ASAP7_75t_R.pex.sp.NOR2XP67_ASAP7_75T_R.pxi"
* BEGIN of "./NOR2xp67_ASAP7_75t_R.pex.sp.NOR2XP67_ASAP7_75T_R.pxi"
* File: NOR2xp67_ASAP7_75t_R.pex.sp.NOR2XP67_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:43:57 2017
* 
x_PM_NOR2XP67_ASAP7_75T_R%A N_A_M0_g N_A_M2_g N_A_c_2_p N_A_M3_g A VSS
+ PM_NOR2XP67_ASAP7_75T_R%A
x_PM_NOR2XP67_ASAP7_75T_R%B N_B_M1_g N_B_M4_g N_B_c_15_n N_B_M5_g B VSS
+ PM_NOR2XP67_ASAP7_75T_R%B
x_PM_NOR2XP67_ASAP7_75T_R%5 N_5_M2_s N_5_c_35_n N_5_M4_s N_5_M3_s N_5_c_41_n
+ N_5_M5_s N_5_c_49_p N_5_c_36_n N_5_c_37_n N_5_c_40_n N_5_c_43_n N_5_c_44_n
+ N_5_c_45_n N_5_c_50_p VSS PM_NOR2XP67_ASAP7_75T_R%5
x_PM_NOR2XP67_ASAP7_75T_R%Y N_Y_M0_d N_Y_M1_s N_Y_c_55_n N_Y_M5_d N_Y_M4_d
+ N_Y_c_68_n N_Y_c_57_n N_Y_c_58_n N_Y_c_61_n N_Y_c_73_n Y N_Y_c_64_n N_Y_c_65_n
+ VSS PM_NOR2XP67_ASAP7_75T_R%Y
cc_1 N_A_M0_g N_B_M1_g 2.60402e-19 $X=0.081 $Y=0.054 $X2=0.189 $Y2=0.054
cc_2 N_A_c_2_p N_B_M1_g 0.0035196f $X=0.135 $Y=0.136 $X2=0.189 $Y2=0.054
cc_3 N_A_c_2_p N_B_c_15_n 0.00183132f $X=0.135 $Y=0.136 $X2=0.243 $Y2=0.136
cc_4 N_A_c_2_p B 0.00437697f $X=0.135 $Y=0.136 $X2=0.243 $Y2=0.134
cc_5 A B 0.00298589f $X=0.081 $Y=0.13 $X2=0.243 $Y2=0.134
cc_6 A N_5_c_35_n 0.00130836f $X=0.081 $Y=0.13 $X2=0.189 $Y2=0.136
cc_7 A N_5_c_36_n 0.0013084f $X=0.081 $Y=0.13 $X2=0 $Y2=0
cc_8 N_A_M0_g N_5_c_37_n 3.94108e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_9 N_A_c_2_p N_5_c_37_n 4.52377e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_10 A N_5_c_37_n 2.8148e-19 $X=0.081 $Y=0.13 $X2=0 $Y2=0
cc_11 N_A_c_2_p N_5_c_40_n 2.34767e-19 $X=0.135 $Y=0.136 $X2=0.243 $Y2=0.135
cc_12 N_A_c_2_p N_Y_c_55_n 0.00464573f $X=0.135 $Y=0.136 $X2=0.243 $Y2=0.136
cc_13 B N_5_c_41_n 6.13941e-19 $X=0.243 $Y=0.134 $X2=0.135 $Y2=0.136
cc_14 B N_5_c_40_n 0.00375045f $X=0.243 $Y=0.134 $X2=0.081 $Y2=0.136
cc_15 B N_5_c_43_n 5.32529e-19 $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_16 N_B_c_15_n N_5_c_44_n 2.2154e-19 $X=0.243 $Y=0.136 $X2=0 $Y2=0
cc_17 N_B_M1_g N_5_c_45_n 4.27122e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_18 B N_5_c_45_n 5.32529e-19 $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_19 B N_Y_c_55_n 0.00386626f $X=0.243 $Y=0.134 $X2=0.135 $Y2=0.136
cc_20 B N_Y_c_57_n 0.00142656f $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_21 N_B_M1_g N_Y_c_58_n 4.30157e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_22 N_B_c_15_n N_Y_c_58_n 7.71399e-19 $X=0.243 $Y=0.136 $X2=0 $Y2=0
cc_23 B N_Y_c_58_n 0.00155911f $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_24 N_B_c_15_n N_Y_c_61_n 5.61351e-19 $X=0.243 $Y=0.136 $X2=0 $Y2=0
cc_25 B N_Y_c_61_n 0.00198568f $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_26 B Y 2.97361e-19 $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_27 B N_Y_c_64_n 5.36266e-19 $X=0.243 $Y=0.134 $X2=0.135 $Y2=0.136
cc_28 N_B_c_15_n N_Y_c_65_n 5.18378e-19 $X=0.243 $Y=0.136 $X2=0 $Y2=0
cc_29 B N_Y_c_65_n 0.00103289f $X=0.243 $Y=0.134 $X2=0 $Y2=0
cc_30 N_5_c_41_n N_Y_c_55_n 5.3737e-19 $X=0.162 $Y=0.216 $X2=0.135 $Y2=0.136
cc_31 N_5_c_41_n N_Y_c_68_n 0.00288888f $X=0.162 $Y=0.216 $X2=0 $Y2=0
cc_32 N_5_c_49_p N_Y_c_68_n 0.00302498f $X=0.268 $Y=0.216 $X2=0 $Y2=0
cc_33 N_5_c_50_p N_Y_c_68_n 0.00250906f $X=0.236 $Y=0.234 $X2=0 $Y2=0
cc_34 N_5_c_41_n N_Y_c_61_n 3.96143e-19 $X=0.162 $Y=0.216 $X2=0 $Y2=0
cc_35 N_5_c_50_p N_Y_c_61_n 0.00352737f $X=0.236 $Y=0.234 $X2=0 $Y2=0
cc_36 N_5_c_49_p N_Y_c_73_n 0.00413386f $X=0.268 $Y=0.216 $X2=0 $Y2=0
cc_37 N_5_c_44_n N_Y_c_73_n 0.00352737f $X=0.27 $Y=0.234 $X2=0 $Y2=0

* END of "./NOR2xp67_ASAP7_75t_R.pex.sp.NOR2XP67_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR3x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:44:19 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR3x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR3x1_ASAP7_75t_R.pex.sp.pex"
* File: NOR3x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:44:19 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR3X1_ASAP7_75T_R%C 5 8 11 14 17 19 31 VSS
c10 31 VSS 0.0226821f $X=0.069 $Y=0.133
c11 17 VSS 0.0141154f $X=0.189 $Y=0.135
c12 14 VSS 0.0633654f $X=0.189 $Y=0.0675
c13 8 VSS 0.0651217f $X=0.135 $Y=0.135
c14 2 VSS 0.0675439f $X=0.081 $Y=0.135
r15 31 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.07 $Y=0.135 $X2=0.07
+ $Y2=0.135
r16 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r18 8 17 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135 $Y=0.135
+ $X2=0.189 $Y2=0.135
r19 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r20 2 8 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081 $Y=0.135
+ $X2=0.135 $Y2=0.135
r21 2 35 11 $w=2e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.081 $Y=0.135
+ $X2=0.07 $Y2=0.135
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
.ends

.subckt PM_NOR3X1_ASAP7_75T_R%B 2 7 10 13 16 19 28 VSS
c27 28 VSS 0.00521604f $X=0.296 $Y=0.133
c28 16 VSS 0.070107f $X=0.351 $Y=0.135
c29 10 VSS 0.0637068f $X=0.297 $Y=0.135
c30 2 VSS 0.0625081f $X=0.243 $Y=0.0675
r31 16 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r32 10 16 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297 $Y=0.135
+ $X2=0.351 $Y2=0.135
r33 10 28 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r34 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r35 5 10 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243 $Y=0.135
+ $X2=0.297 $Y2=0.135
r36 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r37 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_NOR3X1_ASAP7_75T_R%A 2 7 10 13 16 19 30 VSS
c29 30 VSS 0.00203075f $X=0.459 $Y=0.133
c30 16 VSS 0.0741408f $X=0.513 $Y=0.135
c31 10 VSS 0.0645812f $X=0.459 $Y=0.135
c32 2 VSS 0.061821f $X=0.405 $Y=0.0675
r33 16 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r34 10 16 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459 $Y=0.135
+ $X2=0.513 $Y2=0.135
r35 10 30 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r36 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r37 5 10 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405 $Y=0.135
+ $X2=0.459 $Y2=0.135
r38 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r39 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_NOR3X1_ASAP7_75T_R%6 1 2 5 6 7 10 11 12 15 23 24 26 28 29 30 31 VSS
c25 31 VSS 6.15197e-20 $X=0.315 $Y=0.198
c26 30 VSS 7.1588e-20 $X=0.306 $Y=0.198
c27 29 VSS 6.54394e-19 $X=0.256 $Y=0.198
c28 28 VSS 0.0014247f $X=0.234 $Y=0.198
c29 26 VSS 1.81636e-19 $X=0.324 $Y=0.198
c30 24 VSS 0.00103795f $X=0.202 $Y=0.198
c31 23 VSS 0.0106365f $X=0.176 $Y=0.198
c32 15 VSS 0.00275365f $X=0.324 $Y=0.2025
c33 11 VSS 5.7545e-19 $X=0.341 $Y=0.2025
c34 10 VSS 0.00456849f $X=0.216 $Y=0.2025
c35 6 VSS 6.69874e-19 $X=0.233 $Y=0.2025
c36 5 VSS 0.0122657f $X=0.108 $Y=0.2025
c37 1 VSS 6.89902e-19 $X=0.125 $Y=0.2025
r38 30 31 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.198 $X2=0.315 $Y2=0.198
r39 29 30 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.198 $X2=0.306 $Y2=0.198
r40 28 29 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.256 $Y2=0.198
r41 26 31 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.198 $X2=0.315 $Y2=0.198
r42 23 24 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.198 $X2=0.202 $Y2=0.198
r43 21 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.234 $Y2=0.198
r44 21 24 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.202 $Y2=0.198
r45 17 23 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.198 $X2=0.176 $Y2=0.198
r46 15 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198 $X2=0.324
+ $Y2=0.198
r47 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r48 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r49 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r50 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r51 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r52 5 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.198 $X2=0.108
+ $Y2=0.198
r53 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.2025 $X2=0.108 $Y2=0.2025
r54 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.108 $Y2=0.2025
.ends

.subckt PM_NOR3X1_ASAP7_75T_R%7 1 2 5 6 7 10 11 12 15 23 24 26 29 VSS
c28 29 VSS 0.00178544f $X=0.418 $Y=0.234
c29 28 VSS 0.00392508f $X=0.396 $Y=0.234
c30 26 VSS 0.00691197f $X=0.486 $Y=0.234
c31 24 VSS 0.00192468f $X=0.358 $Y=0.234
c32 23 VSS 0.00710134f $X=0.338 $Y=0.234
c33 15 VSS 0.00269882f $X=0.486 $Y=0.2025
c34 11 VSS 6.4978e-19 $X=0.503 $Y=0.2025
c35 10 VSS 0.00329808f $X=0.378 $Y=0.2025
c36 6 VSS 5.38922e-19 $X=0.395 $Y=0.2025
c37 5 VSS 0.00397608f $X=0.27 $Y=0.2025
c38 1 VSS 7.12816e-19 $X=0.287 $Y=0.2025
r39 28 29 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.418 $Y2=0.234
r40 26 29 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.418 $Y2=0.234
r41 23 24 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.234 $X2=0.358 $Y2=0.234
r42 21 28 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r43 21 24 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.358 $Y2=0.234
r44 17 23 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.338 $Y2=0.234
r45 15 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r46 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.486 $Y2=0.2025
r47 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.2025 $X2=0.486 $Y2=0.2025
r48 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r49 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r50 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r51 5 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r52 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.2025 $X2=0.27 $Y2=0.2025
r53 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.27 $Y2=0.2025
.ends

.subckt PM_NOR3X1_ASAP7_75T_R%Y 1 2 6 9 11 12 15 16 19 21 24 28 29 30 31 32 33
+ 34 35 43 44 48 50 VSS
c35 52 VSS 4.55454e-19 $X=0.567 $Y=0.18
c36 50 VSS 0.00151026f $X=0.567 $Y=0.095
c37 49 VSS 0.00104959f $X=0.567 $Y=0.063
c38 48 VSS 0.00374358f $X=0.566 $Y=0.127
c39 46 VSS 4.30151e-19 $X=0.567 $Y=0.189
c40 44 VSS 2.77631e-19 $X=0.5 $Y=0.198
c41 43 VSS 8.46035e-21 $X=0.468 $Y=0.198
c42 35 VSS 0.00420063f $X=0.558 $Y=0.198
c43 34 VSS 0.00414532f $X=0.513 $Y=0.036
c44 33 VSS 0.00575891f $X=0.468 $Y=0.036
c45 32 VSS 0.00868347f $X=0.396 $Y=0.036
c46 31 VSS 0.00311736f $X=0.338 $Y=0.036
c47 30 VSS 0.00887783f $X=0.306 $Y=0.036
c48 29 VSS 0.00446007f $X=0.234 $Y=0.036
c49 28 VSS 0.00700532f $X=0.432 $Y=0.036
c50 24 VSS 0.00988214f $X=0.216 $Y=0.036
c51 21 VSS 0.00782805f $X=0.558 $Y=0.036
c52 19 VSS 0.00107488f $X=0.538 $Y=0.2025
c53 15 VSS 0.00275365f $X=0.432 $Y=0.2025
c54 11 VSS 6.18295e-19 $X=0.449 $Y=0.2025
c55 9 VSS 4.53057e-19 $X=0.43 $Y=0.0675
c56 1 VSS 5.72268e-19 $X=0.233 $Y=0.0675
r57 51 52 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.171 $X2=0.567 $Y2=0.18
r58 49 50 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.063 $X2=0.567 $Y2=0.095
r59 48 51 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.127 $X2=0.567 $Y2=0.171
r60 48 50 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.127 $X2=0.567 $Y2=0.095
r61 46 52 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.567 $Y2=0.18
r62 45 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.045 $X2=0.567 $Y2=0.063
r63 43 44 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.198 $X2=0.5 $Y2=0.198
r64 41 44 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.198 $X2=0.5 $Y2=0.198
r65 37 43 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.198 $X2=0.468 $Y2=0.198
r66 35 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.198 $X2=0.567 $Y2=0.189
r67 35 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.198 $X2=0.54 $Y2=0.198
r68 33 34 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.513 $Y2=0.036
r69 31 32 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.036 $X2=0.396 $Y2=0.036
r70 30 31 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.338 $Y2=0.036
r71 29 30 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.306 $Y2=0.036
r72 27 33 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.468 $Y2=0.036
r73 27 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.396 $Y2=0.036
r74 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r75 23 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.234 $Y2=0.036
r76 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r77 21 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.036 $X2=0.567 $Y2=0.045
r78 21 34 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.513 $Y2=0.036
r79 19 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.198 $X2=0.54
+ $Y2=0.198
r80 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.538 $Y2=0.2025
r81 15 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.198 $X2=0.432
+ $Y2=0.198
r82 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r83 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r84 9 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r85 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.43 $Y2=0.0675
r86 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.216
+ $Y=0.0675 $X2=0.216 $Y2=0.036
r87 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r88 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends


* END of "./NOR3x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR3x1_ASAP7_75t_R  VSS VDD C B A Y
* 
* Y	Y
* A	A
* B	B
* C	C
M0 N_Y_M0_d N_C_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M1 VSS N_B_M1_g N_Y_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M2 N_Y_M2_d N_A_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M3 N_6_M3_d N_C_M3_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M4 N_6_M4_d N_C_M4_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M5 N_6_M5_d N_C_M5_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M6 N_7_M6_d N_B_M6_g N_6_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M7 N_7_M7_d N_B_M7_g N_6_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M8 N_7_M8_d N_B_M8_g N_6_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M9 N_Y_M9_d N_A_M9_g N_7_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M10 N_Y_M10_d N_A_M10_g N_7_M10_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M11 N_Y_M11_d N_A_M11_g N_7_M11_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
*
* 
* .include "NOR3x1_ASAP7_75t_R.pex.sp.NOR3X1_ASAP7_75T_R.pxi"
* BEGIN of "./NOR3x1_ASAP7_75t_R.pex.sp.NOR3X1_ASAP7_75T_R.pxi"
* File: NOR3x1_ASAP7_75t_R.pex.sp.NOR3X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:44:19 2017
* 
x_PM_NOR3X1_ASAP7_75T_R%C N_C_M3_g N_C_c_1_p N_C_M4_g N_C_M0_g N_C_c_4_p
+ N_C_M5_g C VSS PM_NOR3X1_ASAP7_75T_R%C
x_PM_NOR3X1_ASAP7_75T_R%B N_B_M1_g N_B_M6_g N_B_c_13_n N_B_M7_g N_B_c_14_n
+ N_B_M8_g B VSS PM_NOR3X1_ASAP7_75T_R%B
x_PM_NOR3X1_ASAP7_75T_R%A N_A_M2_g N_A_M9_g N_A_c_40_n N_A_M10_g N_A_c_41_n
+ N_A_M11_g A VSS PM_NOR3X1_ASAP7_75T_R%A
x_PM_NOR3X1_ASAP7_75T_R%6 N_6_M4_d N_6_M3_d N_6_c_68_n N_6_M6_s N_6_M5_d
+ N_6_c_80_p N_6_M8_s N_6_M7_s N_6_c_74_n N_6_c_69_n N_6_c_72_n N_6_c_84_p
+ N_6_c_89_p N_6_c_76_n N_6_c_78_n N_6_c_79_n VSS PM_NOR3X1_ASAP7_75T_R%6
x_PM_NOR3X1_ASAP7_75T_R%7 N_7_M7_d N_7_M6_d N_7_c_93_n N_7_M9_s N_7_M8_d
+ N_7_c_97_n N_7_M11_s N_7_M10_s N_7_c_99_n N_7_c_95_n N_7_c_96_n N_7_c_101_n
+ N_7_c_102_n VSS PM_NOR3X1_ASAP7_75T_R%7
x_PM_NOR3X1_ASAP7_75T_R%Y N_Y_M1_s N_Y_M0_d N_Y_M2_d N_Y_c_126_n N_Y_M10_d
+ N_Y_M9_d N_Y_c_128_n N_Y_M11_d N_Y_c_150_n N_Y_c_130_n N_Y_c_120_n N_Y_c_131_n
+ N_Y_c_144_n N_Y_c_121_n N_Y_c_124_n N_Y_c_125_n N_Y_c_133_n N_Y_c_136_n
+ N_Y_c_137_n N_Y_c_138_n N_Y_c_140_n Y N_Y_c_142_n VSS PM_NOR3X1_ASAP7_75T_R%Y
cc_1 N_C_c_1_p N_B_M1_g 2.71887e-19 $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_2 N_C_M0_g N_B_M1_g 0.00357042f $X=0.189 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_3 N_C_M0_g N_B_c_13_n 2.71887e-19 $X=0.189 $Y=0.0675 $X2=0.297 $Y2=0.135
cc_4 N_C_c_4_p N_B_c_14_n 0.00166313f $X=0.189 $Y=0.135 $X2=0.351 $Y2=0.135
cc_5 N_C_c_4_p N_6_M4_d 3.67575e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.0675
cc_6 N_C_c_4_p N_6_c_68_n 0.00203185f $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.135
cc_7 N_C_c_1_p N_6_c_69_n 3.91767e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_8 N_C_c_4_p N_6_c_69_n 0.00173937f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_9 C N_6_c_69_n 5.30913e-19 $X=0.069 $Y=0.133 $X2=0 $Y2=0
cc_10 N_C_M0_g N_6_c_72_n 4.87149e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_11 N_B_c_13_n N_A_M2_g 2.71887e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_12 N_B_c_14_n N_A_M2_g 0.00333077f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_13 N_B_c_14_n N_A_c_40_n 2.71887e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_14 N_B_c_14_n N_A_c_41_n 0.00152609f $X=0.351 $Y=0.135 $X2=0.189 $Y2=0.135
cc_15 B A 8.97702e-19 $X=0.296 $Y=0.133 $X2=0 $Y2=0
cc_16 N_B_c_14_n N_6_M8_s 3.67575e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_17 N_B_c_14_n N_6_c_74_n 0.00203185f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_18 B N_6_c_74_n 3.24853e-19 $X=0.296 $Y=0.133 $X2=0 $Y2=0
cc_19 N_B_M1_g N_6_c_76_n 3.62146e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_20 B N_6_c_76_n 0.00666344f $X=0.296 $Y=0.133 $X2=0 $Y2=0
cc_21 N_B_c_13_n N_6_c_78_n 2.53669e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_22 N_B_c_14_n N_6_c_79_n 4.94606e-19 $X=0.351 $Y=0.135 $X2=0.069 $Y2=0.133
cc_23 N_B_c_14_n N_7_M7_d 3.64199e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 N_B_c_14_n N_7_c_93_n 7.57503e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_25 B N_7_c_93_n 0.00135416f $X=0.296 $Y=0.133 $X2=0.081 $Y2=0.2025
cc_26 N_B_c_13_n N_7_c_95_n 2.38524e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_27 N_B_c_14_n N_7_c_96_n 6.41116e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_28 B N_Y_c_120_n 3.34873e-19 $X=0.296 $Y=0.133 $X2=0 $Y2=0
cc_29 N_B_M1_g N_Y_c_121_n 2.51775e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_B_c_13_n N_Y_c_121_n 2.38524e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_31 B N_Y_c_121_n 0.00668415f $X=0.296 $Y=0.133 $X2=0 $Y2=0
cc_32 N_B_c_14_n N_Y_c_124_n 4.93209e-19 $X=0.351 $Y=0.135 $X2=0.069 $Y2=0.133
cc_33 N_B_c_14_n N_Y_c_125_n 4.61191e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_34 A N_7_c_97_n 3.24853e-19 $X=0.459 $Y=0.133 $X2=0.135 $Y2=0.2025
cc_35 N_A_c_41_n N_7_M11_s 3.67193e-19 $X=0.513 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_36 N_A_c_41_n N_7_c_99_n 0.00203185f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_37 A N_7_c_99_n 3.24853e-19 $X=0.459 $Y=0.133 $X2=0 $Y2=0
cc_38 N_A_c_40_n N_7_c_101_n 2.38524e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_39 N_A_M2_g N_7_c_102_n 3.63745e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_40 A N_7_c_102_n 8.30022e-19 $X=0.459 $Y=0.133 $X2=0 $Y2=0
cc_41 A N_Y_c_126_n 2.44687e-19 $X=0.459 $Y=0.133 $X2=0 $Y2=0
cc_42 N_A_c_41_n N_Y_M10_d 3.58237e-19 $X=0.513 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_43 N_A_c_41_n N_Y_c_128_n 7.57503e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_44 A N_Y_c_128_n 0.00143134f $X=0.459 $Y=0.133 $X2=0 $Y2=0
cc_45 N_A_c_41_n N_Y_c_130_n 2.70934e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_46 N_A_c_41_n N_Y_c_131_n 7.57503e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_47 A N_Y_c_131_n 0.00247906f $X=0.459 $Y=0.133 $X2=0 $Y2=0
cc_48 N_A_M2_g N_Y_c_133_n 2.48462e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_49 N_A_c_40_n N_Y_c_133_n 2.35211e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_50 A N_Y_c_133_n 0.00665787f $X=0.459 $Y=0.133 $X2=0 $Y2=0
cc_51 N_A_c_41_n N_Y_c_136_n 7.51301e-19 $X=0.513 $Y=0.135 $X2=0.07 $Y2=0.135
cc_52 N_A_c_41_n N_Y_c_137_n 4.944e-19 $X=0.513 $Y=0.135 $X2=0.07 $Y2=0.135
cc_53 N_A_c_40_n N_Y_c_138_n 2.53669e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_54 A N_Y_c_138_n 0.00442312f $X=0.459 $Y=0.133 $X2=0 $Y2=0
cc_55 N_A_c_41_n N_Y_c_140_n 8.63627e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.135
cc_56 A Y 0.00102249f $X=0.459 $Y=0.133 $X2=0 $Y2=0
cc_57 A N_Y_c_142_n 0.00102249f $X=0.459 $Y=0.133 $X2=0 $Y2=0
cc_58 N_6_c_80_p N_7_c_93_n 0.00332785f $X=0.216 $Y=0.2025 $X2=0.081 $Y2=0.2025
cc_59 N_6_c_74_n N_7_c_93_n 0.0036466f $X=0.324 $Y=0.2025 $X2=0.081 $Y2=0.2025
cc_60 N_6_c_78_n N_7_c_93_n 0.00238995f $X=0.306 $Y=0.198 $X2=0.081 $Y2=0.2025
cc_61 N_6_c_74_n N_7_c_97_n 0.00350779f $X=0.324 $Y=0.2025 $X2=0.135 $Y2=0.2025
cc_62 N_6_c_84_p N_7_c_97_n 4.49606e-19 $X=0.324 $Y=0.198 $X2=0.135 $Y2=0.2025
cc_63 N_6_c_80_p N_7_c_95_n 4.49606e-19 $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_64 N_6_c_74_n N_7_c_95_n 0.00250914f $X=0.324 $Y=0.2025 $X2=0 $Y2=0
cc_65 N_6_c_78_n N_7_c_95_n 0.00702445f $X=0.306 $Y=0.198 $X2=0 $Y2=0
cc_66 N_6_c_80_p N_Y_c_120_n 0.00138157f $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_67 N_6_c_89_p N_Y_c_144_n 2.34741e-19 $X=0.234 $Y=0.198 $X2=0 $Y2=0
cc_68 N_6_c_79_n N_Y_c_124_n 2.34741e-19 $X=0.315 $Y=0.198 $X2=0.069 $Y2=0.133
cc_69 N_6_c_84_p N_Y_c_138_n 3.04405e-19 $X=0.324 $Y=0.198 $X2=0 $Y2=0
cc_70 N_7_c_97_n N_Y_c_128_n 0.00342927f $X=0.378 $Y=0.2025 $X2=0.351 $Y2=0.135
cc_71 N_7_c_99_n N_Y_c_128_n 0.0036466f $X=0.486 $Y=0.2025 $X2=0.351 $Y2=0.135
cc_72 N_7_c_101_n N_Y_c_128_n 0.00250914f $X=0.486 $Y=0.234 $X2=0.351 $Y2=0.135
cc_73 N_7_c_99_n N_Y_c_150_n 0.00349481f $X=0.486 $Y=0.2025 $X2=0.351 $Y2=0.2025
cc_74 N_7_c_101_n N_Y_c_150_n 3.09693e-19 $X=0.486 $Y=0.234 $X2=0.351 $Y2=0.2025
cc_75 N_7_c_97_n N_Y_c_138_n 4.51951e-19 $X=0.378 $Y=0.2025 $X2=0 $Y2=0
cc_76 N_7_c_101_n N_Y_c_138_n 0.00704516f $X=0.486 $Y=0.234 $X2=0 $Y2=0
cc_77 N_7_c_99_n N_Y_c_140_n 0.00233206f $X=0.486 $Y=0.2025 $X2=0 $Y2=0

* END of "./NOR3x1_ASAP7_75t_R.pex.sp.NOR3X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR3x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:44:42 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR3x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR3x2_ASAP7_75t_R.pex.sp.pex"
* File: NOR3x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:44:42 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR3X2_ASAP7_75T_R%A 2 5 8 11 14 17 19 22 27 30 33 36 39 49 52 54 61
+ 66 VSS
c70 66 VSS 0.00274836f $X=0.894 $Y=0.135
c71 61 VSS 0.00247844f $X=0.183 $Y=0.135
c72 54 VSS 0.00171206f $X=0.894 $Y=0.081
c73 52 VSS 0.0251808f $X=0.894 $Y=0.078
c74 49 VSS 0.00182484f $X=0.183 $Y=0.081
c75 36 VSS 0.074344f $X=0.999 $Y=0.135
c76 30 VSS 0.0649556f $X=0.945 $Y=0.135
c77 22 VSS 0.0621952f $X=0.891 $Y=0.0675
c78 17 VSS 0.00595222f $X=0.189 $Y=0.135
c79 14 VSS 0.0623361f $X=0.189 $Y=0.0675
c80 8 VSS 0.0649686f $X=0.135 $Y=0.135
c81 2 VSS 0.0684308f $X=0.081 $Y=0.135
r82 54 66 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.894
+ $Y=0.081 $X2=0.894 $Y2=0.135
r83 52 54 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.894 $Y=0.081 $X2=0.894
+ $Y2=0.081
r84 49 61 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.183
+ $Y=0.081 $X2=0.183 $Y2=0.135
r85 48 52 48.2778 $w=1.8e-08 $l=7.11e-07 $layer=M2 $thickness=3.6e-08 $X=0.183
+ $Y=0.081 $X2=0.894 $Y2=0.081
r86 48 49 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.183 $Y=0.081 $X2=0.183
+ $Y2=0.081
r87 36 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.999
+ $Y=0.135 $X2=0.999 $Y2=0.2025
r88 30 36 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.945 $Y=0.135
+ $X2=0.999 $Y2=0.135
r89 30 33 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.945
+ $Y=0.135 $X2=0.945 $Y2=0.2025
r90 25 30 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.891 $Y=0.135
+ $X2=0.945 $Y2=0.135
r91 25 66 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.894 $Y=0.135 $X2=0.894
+ $Y2=0.135
r92 25 27 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.135 $X2=0.891 $Y2=0.2025
r93 22 25 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.891
+ $Y=0.0675 $X2=0.891 $Y2=0.135
r94 17 61 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.183 $Y=0.135 $X2=0.183
+ $Y2=0.135
r95 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r96 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r97 8 17 48 $w=2e-08 $l=4.8e-08 $layer=LIG $thickness=5e-08 $X=0.135 $Y=0.135
+ $X2=0.183 $Y2=0.135
r98 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r99 2 8 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081 $Y=0.135
+ $X2=0.135 $Y2=0.135
r100 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
.ends

.subckt PM_NOR3X2_ASAP7_75T_R%B 2 5 8 11 14 17 19 22 27 30 33 36 39 43 44 45 49
+ 50 51 52 55 57 58 VSS
c74 58 VSS 3.98855e-19 $X=0.734 $Y=0.1205
c75 57 VSS 0.00128427f $X=0.734 $Y=0.106
c76 55 VSS 9.44712e-19 $X=0.734 $Y=0.135
c77 52 VSS 3.49249e-19 $X=0.565 $Y=0.072
c78 51 VSS 0.00481358f $X=0.547 $Y=0.072
c79 50 VSS 9.15736e-19 $X=0.356 $Y=0.072
c80 49 VSS 0.0051315f $X=0.725 $Y=0.072
c81 45 VSS 3.69184e-19 $X=0.347 $Y=0.1195
c82 44 VSS 0.00127181f $X=0.347 $Y=0.106
c83 43 VSS 8.81025e-19 $X=0.348 $Y=0.133
c84 36 VSS 0.0706331f $X=0.837 $Y=0.135
c85 30 VSS 0.0640963f $X=0.783 $Y=0.135
c86 22 VSS 0.0630165f $X=0.729 $Y=0.0675
c87 17 VSS 0.00834409f $X=0.351 $Y=0.135
c88 14 VSS 0.0629776f $X=0.351 $Y=0.0675
c89 8 VSS 0.0640813f $X=0.297 $Y=0.135
c90 2 VSS 0.0622537f $X=0.243 $Y=0.135
r91 57 58 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.734
+ $Y=0.106 $X2=0.734 $Y2=0.1205
r92 55 58 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.734
+ $Y=0.135 $X2=0.734 $Y2=0.1205
r93 53 57 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.734
+ $Y=0.081 $X2=0.734 $Y2=0.106
r94 51 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.547
+ $Y=0.072 $X2=0.565 $Y2=0.072
r95 50 51 12.9691 $w=1.8e-08 $l=1.91e-07 $layer=M1 $thickness=3.6e-08 $X=0.356
+ $Y=0.072 $X2=0.547 $Y2=0.072
r96 49 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.725 $Y=0.072 $X2=0.734 $Y2=0.081
r97 49 52 10.8642 $w=1.8e-08 $l=1.6e-07 $layer=M1 $thickness=3.6e-08 $X=0.725
+ $Y=0.072 $X2=0.565 $Y2=0.072
r98 44 45 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.347
+ $Y=0.106 $X2=0.347 $Y2=0.1195
r99 43 45 0.916667 $w=1.8e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.347
+ $Y=0.133 $X2=0.347 $Y2=0.1195
r100 41 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.347 $Y=0.081 $X2=0.356 $Y2=0.072
r101 41 44 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.347
+ $Y=0.081 $X2=0.347 $Y2=0.106
r102 36 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.837 $Y=0.135 $X2=0.837 $Y2=0.2025
r103 30 36 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.783 $Y=0.135
+ $X2=0.837 $Y2=0.135
r104 30 33 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.135 $X2=0.783 $Y2=0.2025
r105 25 30 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729 $Y=0.135
+ $X2=0.783 $Y2=0.135
r106 25 55 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.734 $Y=0.135 $X2=0.734
+ $Y2=0.135
r107 25 27 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.135 $X2=0.729 $Y2=0.2025
r108 22 25 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.135
r109 17 43 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.347 $Y=0.135 $X2=0.347
+ $Y2=0.135
r110 17 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r111 14 17 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r112 8 17 50 $w=2e-08 $l=5e-08 $layer=LIG $thickness=5e-08 $X=0.297 $Y=0.135
+ $X2=0.347 $Y2=0.135
r113 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r114 2 8 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243 $Y=0.135
+ $X2=0.297 $Y2=0.135
r115 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
.ends

.subckt PM_NOR3X2_ASAP7_75T_R%C 2 7 10 13 16 19 22 25 28 31 34 37 39 42 VSS
c41 42 VSS 0.00152202f $X=0.555 $Y=0.133
c42 37 VSS 0.0203793f $X=0.675 $Y=0.135
c43 34 VSS 0.062961f $X=0.675 $Y=0.0675
c44 28 VSS 0.0644377f $X=0.621 $Y=0.135
c45 22 VSS 0.0653595f $X=0.567 $Y=0.135
c46 16 VSS 0.06505f $X=0.513 $Y=0.135
c47 10 VSS 0.0644495f $X=0.459 $Y=0.135
c48 2 VSS 0.0629441f $X=0.405 $Y=0.0675
r49 42 45 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.556 $Y=0.135 $X2=0.556
+ $Y2=0.135
r50 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.2025
r51 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0675 $X2=0.675 $Y2=0.135
r52 28 37 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621 $Y=0.135
+ $X2=0.675 $Y2=0.135
r53 28 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r54 22 28 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.567 $Y=0.135
+ $X2=0.621 $Y2=0.135
r55 22 45 11 $w=2e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.567 $Y=0.135
+ $X2=0.556 $Y2=0.135
r56 22 25 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r57 16 45 43 $w=2e-08 $l=4.3e-08 $layer=LIG $thickness=5e-08 $X=0.513 $Y=0.135
+ $X2=0.556 $Y2=0.135
r58 16 19 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r59 10 16 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459 $Y=0.135
+ $X2=0.513 $Y2=0.135
r60 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r61 5 10 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405 $Y=0.135
+ $X2=0.459 $Y2=0.135
r62 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r63 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_NOR3X2_ASAP7_75T_R%6 1 2 5 6 7 10 11 12 15 23 24 25 28 30 31 VSS
c27 31 VSS 0.00267306f $X=0.29 $Y=0.234
c28 30 VSS 0.00383338f $X=0.256 $Y=0.234
c29 28 VSS 0.00453277f $X=0.324 $Y=0.234
c30 26 VSS 3.19325e-19 $X=0.2135 $Y=0.234
c31 25 VSS 0.00193913f $X=0.211 $Y=0.234
c32 24 VSS 0.00129872f $X=0.192 $Y=0.234
c33 23 VSS 0.00695592f $X=0.176 $Y=0.234
c34 15 VSS 0.00475672f $X=0.324 $Y=0.2025
c35 11 VSS 7.17878e-19 $X=0.341 $Y=0.2025
c36 10 VSS 0.00347287f $X=0.216 $Y=0.2025
c37 6 VSS 5.38922e-19 $X=0.233 $Y=0.2025
c38 5 VSS 0.00269882f $X=0.108 $Y=0.2025
c39 1 VSS 6.4978e-19 $X=0.125 $Y=0.2025
r40 30 31 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.234 $X2=0.29 $Y2=0.234
r41 28 31 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.29 $Y2=0.234
r42 25 26 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.211
+ $Y=0.234 $X2=0.2135 $Y2=0.234
r43 24 25 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.192
+ $Y=0.234 $X2=0.211 $Y2=0.234
r44 23 24 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.176
+ $Y=0.234 $X2=0.192 $Y2=0.234
r45 21 30 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.256 $Y2=0.234
r46 21 26 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.2135 $Y2=0.234
r47 17 23 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.176 $Y2=0.234
r48 15 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r49 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r50 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r51 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r52 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r53 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r54 5 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r55 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.2025 $X2=0.108 $Y2=0.2025
r56 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.108 $Y2=0.2025
.ends

.subckt PM_NOR3X2_ASAP7_75T_R%7 1 2 5 6 7 10 11 12 15 16 17 20 21 22 25 26 27 30
+ 38 39 43 48 49 53 54 56 59 61 VSS
c53 61 VSS 2.78809e-19 $X=0.7765 $Y=0.198
c54 59 VSS 5.17444e-19 $X=0.742 $Y=0.198
c55 58 VSS 0.00203085f $X=0.725 $Y=0.198
c56 56 VSS 2.97451e-19 $X=0.81 $Y=0.198
c57 54 VSS 7.11849e-19 $X=0.682 $Y=0.198
c58 53 VSS 0.0106025f $X=0.662 $Y=0.198
c59 49 VSS 0.00240114f $X=0.565 $Y=0.198
c60 48 VSS 0.00978135f $X=0.547 $Y=0.198
c61 44 VSS 0.0051489f $X=0.452 $Y=0.198
c62 43 VSS 0.00262736f $X=0.418 $Y=0.198
c63 39 VSS 5.46526e-19 $X=0.356 $Y=0.198
c64 38 VSS 5.72503e-19 $X=0.338 $Y=0.198
c65 30 VSS 0.0027527f $X=0.81 $Y=0.2025
c66 26 VSS 5.75435e-19 $X=0.827 $Y=0.2025
c67 25 VSS 0.00438161f $X=0.702 $Y=0.2025
c68 21 VSS 6.69874e-19 $X=0.719 $Y=0.2025
c69 20 VSS 0.0125184f $X=0.594 $Y=0.2025
c70 16 VSS 6.05897e-19 $X=0.611 $Y=0.2025
c71 15 VSS 0.0124222f $X=0.486 $Y=0.2025
c72 11 VSS 6.05897e-19 $X=0.503 $Y=0.2025
c73 10 VSS 0.00438003f $X=0.378 $Y=0.2025
c74 6 VSS 6.69874e-19 $X=0.395 $Y=0.2025
c75 5 VSS 0.00274973f $X=0.27 $Y=0.2025
c76 1 VSS 5.76015e-19 $X=0.287 $Y=0.2025
r77 60 61 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.743
+ $Y=0.198 $X2=0.7765 $Y2=0.198
r78 59 60 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.742
+ $Y=0.198 $X2=0.743 $Y2=0.198
r79 58 59 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.725
+ $Y=0.198 $X2=0.742 $Y2=0.198
r80 56 61 2.27469 $w=1.8e-08 $l=3.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.198 $X2=0.7765 $Y2=0.198
r81 53 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.662
+ $Y=0.198 $X2=0.682 $Y2=0.198
r82 51 58 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.198 $X2=0.725 $Y2=0.198
r83 51 54 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.198 $X2=0.682 $Y2=0.198
r84 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.547
+ $Y=0.198 $X2=0.565 $Y2=0.198
r85 46 53 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.198 $X2=0.662 $Y2=0.198
r86 46 49 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.198 $X2=0.565 $Y2=0.198
r87 43 44 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.198 $X2=0.452 $Y2=0.198
r88 41 48 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.198 $X2=0.547 $Y2=0.198
r89 41 44 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.198 $X2=0.452 $Y2=0.198
r90 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.198 $X2=0.356 $Y2=0.198
r91 36 43 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.198 $X2=0.418 $Y2=0.198
r92 36 39 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.198 $X2=0.356 $Y2=0.198
r93 32 38 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.198 $X2=0.338 $Y2=0.198
r94 30 56 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.198 $X2=0.81
+ $Y2=0.198
r95 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.2025 $X2=0.81 $Y2=0.2025
r96 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.827 $Y=0.2025 $X2=0.81 $Y2=0.2025
r97 25 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.198 $X2=0.702
+ $Y2=0.198
r98 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2025 $X2=0.702 $Y2=0.2025
r99 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.2025 $X2=0.702 $Y2=0.2025
r100 20 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.198
+ $X2=0.594 $Y2=0.198
r101 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2025 $X2=0.594 $Y2=0.2025
r102 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2025 $X2=0.594 $Y2=0.2025
r103 15 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.198
+ $X2=0.486 $Y2=0.198
r104 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.486 $Y2=0.2025
r105 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.2025 $X2=0.486 $Y2=0.2025
r106 10 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.198
+ $X2=0.378 $Y2=0.198
r107 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r108 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r109 5 32 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.198 $X2=0.27
+ $Y2=0.198
r110 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r111 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
.ends

.subckt PM_NOR3X2_ASAP7_75T_R%8 1 2 5 6 7 10 11 12 15 23 24 26 30 VSS
c26 31 VSS 1.63466e-19 $X=0.904 $Y=0.234
c27 30 VSS 0.00140149f $X=0.903 $Y=0.234
c28 29 VSS 0.00181697f $X=0.885 $Y=0.234
c29 28 VSS 0.00201427f $X=0.866 $Y=0.234
c30 26 VSS 0.00696456f $X=0.972 $Y=0.234
c31 24 VSS 0.00181142f $X=0.844 $Y=0.234
c32 23 VSS 0.00715189f $X=0.824 $Y=0.234
c33 15 VSS 0.00269882f $X=0.972 $Y=0.2025
c34 11 VSS 6.48198e-19 $X=0.989 $Y=0.2025
c35 10 VSS 0.00341054f $X=0.864 $Y=0.2025
c36 6 VSS 5.38922e-19 $X=0.881 $Y=0.2025
c37 5 VSS 0.00472107f $X=0.756 $Y=0.2025
c38 1 VSS 7.13675e-19 $X=0.773 $Y=0.2025
r39 30 31 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.903
+ $Y=0.234 $X2=0.904 $Y2=0.234
r40 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.885
+ $Y=0.234 $X2=0.903 $Y2=0.234
r41 28 29 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.866
+ $Y=0.234 $X2=0.885 $Y2=0.234
r42 26 31 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.972
+ $Y=0.234 $X2=0.904 $Y2=0.234
r43 23 24 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.824
+ $Y=0.234 $X2=0.844 $Y2=0.234
r44 21 28 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.866 $Y2=0.234
r45 21 24 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.864
+ $Y=0.234 $X2=0.844 $Y2=0.234
r46 17 23 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.824 $Y2=0.234
r47 15 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.234 $X2=0.972
+ $Y2=0.234
r48 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.2025 $X2=0.972 $Y2=0.2025
r49 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.989 $Y=0.2025 $X2=0.972 $Y2=0.2025
r50 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.864 $Y=0.234 $X2=0.864
+ $Y2=0.234
r51 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.847 $Y=0.2025 $X2=0.864 $Y2=0.2025
r52 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.881 $Y=0.2025 $X2=0.864 $Y2=0.2025
r53 5 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234 $X2=0.756
+ $Y2=0.234
r54 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.2025 $X2=0.756 $Y2=0.2025
r55 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.2025 $X2=0.756 $Y2=0.2025
.ends

.subckt PM_NOR3X2_ASAP7_75T_R%Y 1 6 7 11 12 16 21 24 26 27 30 31 32 35 36 39 44
+ 45 49 52 53 54 55 56 59 62 63 64 65 66 68 74 76 77 88 89 93 95 VSS
c77 97 VSS 6.6224e-20 $X=1.053 $Y=0.164
c78 95 VSS 0.00172644f $X=1.053 $Y=0.095
c79 94 VSS 9.47077e-19 $X=1.053 $Y=0.063
c80 93 VSS 0.00353169f $X=1.052 $Y=0.127
c81 91 VSS 0.00101778f $X=1.053 $Y=0.189
c82 89 VSS 7.12898e-19 $X=1.006 $Y=0.198
c83 88 VSS 6.13025e-19 $X=0.986 $Y=0.198
c84 80 VSS 0.00405642f $X=1.044 $Y=0.198
c85 77 VSS 3.04498e-19 $X=0.128 $Y=0.198
c86 76 VSS 0.00279066f $X=0.094 $Y=0.198
c87 74 VSS 4.5381e-19 $X=0.162 $Y=0.198
c88 69 VSS 0.0019505f $X=0.036 $Y=0.198
c89 68 VSS 6.76809e-19 $X=0.911 $Y=0.036
c90 66 VSS 0.00423963f $X=0.903 $Y=0.036
c91 65 VSS 0.00578947f $X=0.866 $Y=0.036
c92 64 VSS 0.0103422f $X=0.824 $Y=0.036
c93 63 VSS 0.0385756f $X=0.743 $Y=0.036
c94 62 VSS 0.00686016f $X=0.918 $Y=0.036
c95 59 VSS 0.0105087f $X=0.702 $Y=0.036
c96 56 VSS 0.0103888f $X=0.338 $Y=0.036
c97 55 VSS 0.00631091f $X=0.256 $Y=0.036
c98 54 VSS 0.00404191f $X=0.211 $Y=0.036
c99 53 VSS 0.0126481f $X=0.174 $Y=0.036
c100 52 VSS 0.0106828f $X=0.378 $Y=0.036
c101 49 VSS 0.00716926f $X=0.162 $Y=0.036
c102 46 VSS 0.00354522f $X=0.036 $Y=0.036
c103 45 VSS 0.0156892f $X=1.044 $Y=0.036
c104 44 VSS 0.00534065f $X=0.027 $Y=0.164
c105 43 VSS 9.47077e-19 $X=0.027 $Y=0.063
c106 42 VSS 0.00101778f $X=0.027 $Y=0.189
c107 39 VSS 0.00107488f $X=1.024 $Y=0.2025
c108 35 VSS 0.0027527f $X=0.918 $Y=0.2025
c109 31 VSS 5.9588e-19 $X=0.935 $Y=0.2025
c110 30 VSS 0.00278521f $X=0.162 $Y=0.2025
c111 26 VSS 6.95677e-19 $X=0.179 $Y=0.2025
c112 24 VSS 7.39942e-19 $X=0.056 $Y=0.2025
c113 21 VSS 3.34937e-19 $X=0.071 $Y=0.2025
c114 19 VSS 6.29922e-19 $X=0.916 $Y=0.0675
c115 11 VSS 5.97768e-19 $X=0.719 $Y=0.0675
c116 6 VSS 5.97768e-19 $X=0.395 $Y=0.0675
c117 1 VSS 5.4394e-19 $X=0.179 $Y=0.0675
r118 96 97 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.162 $X2=1.053 $Y2=0.164
r119 94 95 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.063 $X2=1.053 $Y2=0.095
r120 93 96 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.127 $X2=1.053 $Y2=0.162
r121 93 95 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.127 $X2=1.053 $Y2=0.095
r122 91 97 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.189 $X2=1.053 $Y2=0.164
r123 90 94 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.045 $X2=1.053 $Y2=0.063
r124 88 89 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.986
+ $Y=0.198 $X2=1.006 $Y2=0.198
r125 86 89 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=1.026
+ $Y=0.198 $X2=1.006 $Y2=0.198
r126 82 88 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.198 $X2=0.986 $Y2=0.198
r127 80 91 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.198 $X2=1.053 $Y2=0.189
r128 80 86 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.198 $X2=1.026 $Y2=0.198
r129 76 77 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.198 $X2=0.128 $Y2=0.198
r130 74 77 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.198 $X2=0.128 $Y2=0.198
r131 71 76 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.198 $X2=0.094 $Y2=0.198
r132 69 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.198 $X2=0.054 $Y2=0.198
r133 67 68 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.904
+ $Y=0.036 $X2=0.911 $Y2=0.036
r134 66 67 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.903
+ $Y=0.036 $X2=0.904 $Y2=0.036
r135 65 66 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.866
+ $Y=0.036 $X2=0.903 $Y2=0.036
r136 64 65 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.824
+ $Y=0.036 $X2=0.866 $Y2=0.036
r137 63 64 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.743
+ $Y=0.036 $X2=0.824 $Y2=0.036
r138 61 68 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.918
+ $Y=0.036 $X2=0.911 $Y2=0.036
r139 61 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.036
+ $X2=0.918 $Y2=0.036
r140 58 63 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.036 $X2=0.743 $Y2=0.036
r141 58 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.036
+ $X2=0.702 $Y2=0.036
r142 55 56 5.5679 $w=1.8e-08 $l=8.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.036 $X2=0.338 $Y2=0.036
r143 54 55 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.211
+ $Y=0.036 $X2=0.256 $Y2=0.036
r144 53 54 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.174
+ $Y=0.036 $X2=0.211 $Y2=0.036
r145 51 58 22 $w=1.8e-08 $l=3.24e-07 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.702 $Y2=0.036
r146 51 56 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.338 $Y2=0.036
r147 51 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036
+ $X2=0.378 $Y2=0.036
r148 48 53 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.174 $Y2=0.036
r149 48 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r150 46 48 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.162 $Y2=0.036
r151 45 90 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.036 $X2=1.053 $Y2=0.045
r152 45 61 8.55556 $w=1.8e-08 $l=1.26e-07 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=0.918 $Y2=0.036
r153 43 44 6.85802 $w=1.8e-08 $l=1.01e-07 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.063 $X2=0.027 $Y2=0.164
r154 42 69 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.189 $X2=0.036 $Y2=0.198
r155 42 44 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.189 $X2=0.027 $Y2=0.164
r156 41 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r157 41 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.063
r158 39 86 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=1.026 $Y=0.198
+ $X2=1.026 $Y2=0.198
r159 36 39 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=1.009 $Y=0.2025 $X2=1.024 $Y2=0.2025
r160 35 82 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.918 $Y=0.198
+ $X2=0.918 $Y2=0.198
r161 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.2025 $X2=0.918 $Y2=0.2025
r162 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.935 $Y=0.2025 $X2=0.918 $Y2=0.2025
r163 30 74 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.198
+ $X2=0.162 $Y2=0.198
r164 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r165 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r166 24 71 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.198
+ $X2=0.054 $Y2=0.198
r167 21 24 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r168 19 62 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.918 $Y=0.0675 $X2=0.918 $Y2=0.036
r169 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.901 $Y=0.0675 $X2=0.916 $Y2=0.0675
r170 15 59 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.702 $Y=0.0675 $X2=0.702 $Y2=0.036
r171 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.0675 $X2=0.702 $Y2=0.0675
r172 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.0675 $X2=0.702 $Y2=0.0675
r173 10 52 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.378 $Y=0.0675 $X2=0.378 $Y2=0.036
r174 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.378 $Y2=0.0675
r175 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.0675 $X2=0.378 $Y2=0.0675
r176 4 49 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r177 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.164 $Y2=0.0675
.ends


* END of "./NOR3x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR3x2_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 VSS N_A_M0_g N_Y_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M1 N_Y_M1_d N_B_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M2 VSS N_C_M2_g N_Y_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M3 VSS N_C_M3_g N_Y_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665 $Y=0.027
M4 N_Y_M4_d N_B_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M5 VSS N_A_M5_g N_Y_M5_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.881 $Y=0.027
M6 N_Y_M6_d N_A_M6_g N_6_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 N_Y_M7_d N_A_M7_g N_6_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 N_Y_M8_d N_A_M8_g N_6_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 N_6_M9_d N_B_M9_g N_7_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 N_6_M10_d N_B_M10_g N_7_M10_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_6_M11_d N_B_M11_g N_7_M11_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M12 VDD N_C_M12_g N_7_M12_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M13 VDD N_C_M13_g N_7_M13_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M14 VDD N_C_M14_g N_7_M14_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M15 VDD N_C_M15_g N_7_M15_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M16 VDD N_C_M16_g N_7_M16_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M17 VDD N_C_M17_g N_7_M17_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
M18 N_8_M18_d N_B_M18_g N_7_M18_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M19 N_8_M19_d N_B_M19_g N_7_M19_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
M20 N_8_M20_d N_B_M20_g N_7_M20_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.827
+ $Y=0.162
M21 N_Y_M21_d N_A_M21_g N_8_M21_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.881
+ $Y=0.162
M22 N_Y_M22_d N_A_M22_g N_8_M22_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.162
M23 N_Y_M23_d N_A_M23_g N_8_M23_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
*
* 
* .include "NOR3x2_ASAP7_75t_R.pex.sp.NOR3X2_ASAP7_75T_R.pxi"
* BEGIN of "./NOR3x2_ASAP7_75t_R.pex.sp.NOR3X2_ASAP7_75T_R.pxi"
* File: NOR3x2_ASAP7_75t_R.pex.sp.NOR3X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:44:42 2017
* 
x_PM_NOR3X2_ASAP7_75T_R%A N_A_c_48_p N_A_M6_g N_A_c_1_p N_A_M7_g N_A_M0_g
+ N_A_c_4_p N_A_M8_g N_A_M5_g N_A_M21_g N_A_c_8_p N_A_M22_g N_A_c_9_p N_A_M23_g
+ N_A_c_41_p A N_A_c_57_p N_A_c_12_p N_A_c_18_p VSS PM_NOR3X2_ASAP7_75T_R%A
x_PM_NOR3X2_ASAP7_75T_R%B N_B_c_71_n N_B_M9_g N_B_c_73_n N_B_M10_g N_B_M1_g
+ N_B_c_74_n N_B_M11_g N_B_M4_g N_B_M18_g N_B_c_76_n N_B_M19_g N_B_c_77_n
+ N_B_M20_g B N_B_c_81_n N_B_c_106_p N_B_c_83_n N_B_c_84_n N_B_c_85_n N_B_c_86_n
+ N_B_c_126_p N_B_c_87_n N_B_c_108_p VSS PM_NOR3X2_ASAP7_75T_R%B
x_PM_NOR3X2_ASAP7_75T_R%C N_C_M2_g N_C_M12_g N_C_c_150_n N_C_M13_g N_C_c_152_n
+ N_C_M14_g N_C_c_153_n N_C_M15_g N_C_c_154_n N_C_M16_g N_C_M3_g N_C_c_145_n
+ N_C_M17_g C VSS PM_NOR3X2_ASAP7_75T_R%C
x_PM_NOR3X2_ASAP7_75T_R%6 N_6_M7_s N_6_M6_s N_6_c_187_n N_6_M9_d N_6_M8_s
+ N_6_c_197_p N_6_M11_d N_6_M10_d N_6_c_193_n N_6_c_188_n N_6_c_189_n
+ N_6_c_191_n N_6_c_194_n N_6_c_195_n N_6_c_199_p VSS PM_NOR3X2_ASAP7_75T_R%6
x_PM_NOR3X2_ASAP7_75T_R%7 N_7_M10_s N_7_M9_s N_7_c_217_n N_7_M12_s N_7_M11_s
+ N_7_c_246_n N_7_M14_s N_7_M13_s N_7_c_231_n N_7_M16_s N_7_M15_s N_7_c_233_n
+ N_7_M18_s N_7_M17_s N_7_c_251_p N_7_M20_s N_7_M19_s N_7_c_219_n N_7_c_213_n
+ N_7_c_222_n N_7_c_214_n N_7_c_236_n N_7_c_238_n N_7_c_225_n N_7_c_242_n
+ N_7_c_226_n N_7_c_227_n N_7_c_215_n VSS PM_NOR3X2_ASAP7_75T_R%7
x_PM_NOR3X2_ASAP7_75T_R%8 N_8_M19_d N_8_M18_d N_8_c_273_n N_8_M21_s N_8_M20_d
+ N_8_c_279_n N_8_M23_s N_8_M22_s N_8_c_267_n N_8_c_274_n N_8_c_268_n
+ N_8_c_269_n N_8_c_270_n VSS PM_NOR3X2_ASAP7_75T_R%8
x_PM_NOR3X2_ASAP7_75T_R%Y N_Y_M0_s N_Y_M2_s N_Y_M1_d N_Y_M4_d N_Y_M3_s N_Y_M5_s
+ N_Y_M6_d N_Y_c_346_n N_Y_M8_d N_Y_M7_d N_Y_c_293_n N_Y_M22_d N_Y_M21_d
+ N_Y_c_295_n N_Y_M23_d N_Y_c_364_n N_Y_c_296_n N_Y_c_298_n N_Y_c_300_n
+ N_Y_c_303_n N_Y_c_304_n N_Y_c_307_n N_Y_c_309_n N_Y_c_331_n N_Y_c_310_n
+ N_Y_c_311_n N_Y_c_334_n N_Y_c_314_n N_Y_c_339_n N_Y_c_315_n N_Y_c_317_n
+ N_Y_c_318_n N_Y_c_319_n N_Y_c_352_n N_Y_c_321_n N_Y_c_323_n Y N_Y_c_326_n VSS
+ PM_NOR3X2_ASAP7_75T_R%Y
cc_1 N_A_c_1_p N_B_c_71_n 2.71887e-19 $X=0.135 $Y=0.135 $X2=0.243 $Y2=0.135
cc_2 N_A_M0_g N_B_c_71_n 0.00333077f $X=0.189 $Y=0.0675 $X2=0.243 $Y2=0.135
cc_3 N_A_M0_g N_B_c_73_n 2.71887e-19 $X=0.189 $Y=0.0675 $X2=0.297 $Y2=0.135
cc_4 N_A_c_4_p N_B_c_74_n 0.00148959f $X=0.189 $Y=0.135 $X2=0.351 $Y2=0.135
cc_5 A N_B_c_74_n 0.00167219f $X=0.894 $Y=0.078 $X2=0.351 $Y2=0.135
cc_6 N_A_M5_g N_B_c_76_n 2.71887e-19 $X=0.891 $Y=0.0675 $X2=0.783 $Y2=0.135
cc_7 N_A_M5_g N_B_c_77_n 0.00333077f $X=0.891 $Y=0.0675 $X2=0.837 $Y2=0.135
cc_8 N_A_c_8_p N_B_c_77_n 2.71887e-19 $X=0.945 $Y=0.135 $X2=0.837 $Y2=0.135
cc_9 N_A_c_9_p N_B_c_77_n 0.00147123f $X=0.999 $Y=0.135 $X2=0.837 $Y2=0.135
cc_10 A N_B_c_77_n 0.00167219f $X=0.894 $Y=0.078 $X2=0.837 $Y2=0.135
cc_11 A N_B_c_81_n 6.70023e-19 $X=0.894 $Y=0.078 $X2=0.347 $Y2=0.106
cc_12 N_A_c_12_p N_B_c_81_n 7.06357e-19 $X=0.183 $Y=0.135 $X2=0.347 $Y2=0.106
cc_13 A N_B_c_83_n 0.00498306f $X=0.894 $Y=0.078 $X2=0.725 $Y2=0.072
cc_14 A N_B_c_84_n 6.61822e-19 $X=0.894 $Y=0.078 $X2=0.356 $Y2=0.072
cc_15 A N_B_c_85_n 0.00522817f $X=0.894 $Y=0.078 $X2=0.547 $Y2=0.072
cc_16 A N_B_c_86_n 4.52398e-19 $X=0.894 $Y=0.078 $X2=0.565 $Y2=0.072
cc_17 A N_B_c_87_n 6.68469e-19 $X=0.894 $Y=0.078 $X2=0.734 $Y2=0.106
cc_18 N_A_c_18_p N_B_c_87_n 7.19714e-19 $X=0.894 $Y=0.135 $X2=0.734 $Y2=0.106
cc_19 A N_C_c_145_n 0.00401629f $X=0.894 $Y=0.078 $X2=0 $Y2=0
cc_20 A C 3.78779e-19 $X=0.894 $Y=0.078 $X2=0.347 $Y2=0.133
cc_21 N_A_c_4_p N_6_M7_s 3.67193e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.135
cc_22 N_A_c_4_p N_6_c_187_n 0.00203185f $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.2025
cc_23 N_A_c_1_p N_6_c_188_n 2.65027e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_24 N_A_M0_g N_6_c_189_n 2.58643e-19 $X=0.189 $Y=0.0675 $X2=0.729 $Y2=0.135
cc_25 N_A_c_12_p N_6_c_189_n 4.7743e-19 $X=0.183 $Y=0.135 $X2=0.729 $Y2=0.135
cc_26 A N_6_c_191_n 5.9683e-19 $X=0.894 $Y=0.078 $X2=0.729 $Y2=0.135
cc_27 A N_7_c_213_n 9.00135e-19 $X=0.894 $Y=0.078 $X2=0.837 $Y2=0.2025
cc_28 A N_7_c_214_n 0.00374227f $X=0.894 $Y=0.078 $X2=0.348 $Y2=0.133
cc_29 A N_7_c_215_n 8.86139e-19 $X=0.894 $Y=0.078 $X2=0.243 $Y2=0.135
cc_30 N_A_c_9_p N_8_M23_s 3.67193e-19 $X=0.999 $Y=0.135 $X2=0.297 $Y2=0.2025
cc_31 N_A_c_9_p N_8_c_267_n 0.00203185f $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_32 A N_8_c_268_n 5.67277e-19 $X=0.894 $Y=0.078 $X2=0.729 $Y2=0.135
cc_33 N_A_c_8_p N_8_c_269_n 2.65027e-19 $X=0.945 $Y=0.135 $X2=0.729 $Y2=0.2025
cc_34 N_A_M5_g N_8_c_270_n 3.11408e-19 $X=0.891 $Y=0.0675 $X2=0.783 $Y2=0.135
cc_35 N_A_c_18_p N_8_c_270_n 4.96853e-19 $X=0.894 $Y=0.135 $X2=0.783 $Y2=0.135
cc_36 N_A_c_4_p N_Y_M8_d 3.39222e-19 $X=0.189 $Y=0.135 $X2=0.729 $Y2=0.2025
cc_37 N_A_c_4_p N_Y_c_293_n 7.57503e-19 $X=0.189 $Y=0.135 $X2=0.783 $Y2=0.135
cc_38 N_A_c_9_p N_Y_M22_d 3.56132e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_39 N_A_c_9_p N_Y_c_295_n 7.57503e-19 $X=0.999 $Y=0.135 $X2=0.837 $Y2=0.135
cc_40 N_A_c_4_p N_Y_c_296_n 3.56528e-19 $X=0.189 $Y=0.135 $X2=0.347 $Y2=0.106
cc_41 N_A_c_41_p N_Y_c_296_n 0.00101083f $X=0.183 $Y=0.081 $X2=0.347 $Y2=0.106
cc_42 N_A_c_8_p N_Y_c_298_n 4.62055e-19 $X=0.945 $Y=0.135 $X2=0.347 $Y2=0.1195
cc_43 N_A_c_9_p N_Y_c_298_n 5.55762e-19 $X=0.999 $Y=0.135 $X2=0.347 $Y2=0.1195
cc_44 N_A_c_4_p N_Y_c_300_n 7.57503e-19 $X=0.189 $Y=0.135 $X2=0.725 $Y2=0.072
cc_45 N_A_c_41_p N_Y_c_300_n 7.78109e-19 $X=0.183 $Y=0.081 $X2=0.725 $Y2=0.072
cc_46 A N_Y_c_300_n 2.39784e-19 $X=0.894 $Y=0.078 $X2=0.725 $Y2=0.072
cc_47 A N_Y_c_303_n 3.68996e-19 $X=0.894 $Y=0.078 $X2=0.565 $Y2=0.072
cc_48 N_A_c_48_p N_Y_c_304_n 5.55762e-19 $X=0.081 $Y=0.135 $X2=0.734 $Y2=0.081
cc_49 N_A_c_1_p N_Y_c_304_n 4.62055e-19 $X=0.135 $Y=0.135 $X2=0.734 $Y2=0.081
cc_50 N_A_c_4_p N_Y_c_304_n 8.58361e-19 $X=0.189 $Y=0.135 $X2=0.734 $Y2=0.081
cc_51 N_A_M0_g N_Y_c_307_n 2.63908e-19 $X=0.189 $Y=0.0675 $X2=0.734 $Y2=0.135
cc_52 N_A_c_41_p N_Y_c_307_n 0.00371636f $X=0.183 $Y=0.081 $X2=0.734 $Y2=0.135
cc_53 A N_Y_c_309_n 0.00228933f $X=0.894 $Y=0.078 $X2=0.734 $Y2=0.135
cc_54 A N_Y_c_310_n 3.68996e-19 $X=0.894 $Y=0.078 $X2=0 $Y2=0
cc_55 N_A_c_9_p N_Y_c_311_n 7.57503e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_56 A N_Y_c_311_n 2.84578e-19 $X=0.894 $Y=0.078 $X2=0 $Y2=0
cc_57 N_A_c_57_p N_Y_c_311_n 0.00136727f $X=0.894 $Y=0.081 $X2=0 $Y2=0
cc_58 A N_Y_c_314_n 0.00223503f $X=0.894 $Y=0.078 $X2=0.347 $Y2=0.135
cc_59 N_A_M5_g N_Y_c_315_n 2.5731e-19 $X=0.891 $Y=0.0675 $X2=0.729 $Y2=0.135
cc_60 N_A_c_57_p N_Y_c_315_n 0.00373008f $X=0.894 $Y=0.081 $X2=0.729 $Y2=0.135
cc_61 N_A_c_9_p N_Y_c_317_n 8.88792e-19 $X=0.999 $Y=0.135 $X2=0.783 $Y2=0.135
cc_62 N_A_c_1_p N_Y_c_318_n 3.34178e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_63 N_A_c_48_p N_Y_c_319_n 4.944e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_64 N_A_c_4_p N_Y_c_319_n 0.0015591f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_65 N_A_c_8_p N_Y_c_321_n 3.99019e-19 $X=0.945 $Y=0.135 $X2=0 $Y2=0
cc_66 N_A_c_9_p N_Y_c_321_n 0.00158095f $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_67 N_A_c_9_p N_Y_c_323_n 4.2024e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_68 N_A_c_9_p Y 3.57243e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_69 N_A_c_18_p Y 4.73012e-19 $X=0.894 $Y=0.135 $X2=0 $Y2=0
cc_70 N_A_c_57_p N_Y_c_326_n 4.73012e-19 $X=0.894 $Y=0.081 $X2=0 $Y2=0
cc_71 N_B_c_73_n N_C_M2_g 2.71887e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_72 N_B_M1_g N_C_M2_g 0.00357042f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_73 N_B_c_85_n N_C_M2_g 4.95866e-19 $X=0.547 $Y=0.072 $X2=0.081 $Y2=0.135
cc_74 N_B_M1_g N_C_c_150_n 2.71887e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.2025
cc_75 N_B_c_85_n N_C_c_150_n 4.95866e-19 $X=0.547 $Y=0.072 $X2=0.135 $Y2=0.2025
cc_76 N_B_c_85_n N_C_c_152_n 6.8328e-19 $X=0.547 $Y=0.072 $X2=0.189 $Y2=0.135
cc_77 N_B_c_83_n N_C_c_153_n 4.01427e-19 $X=0.725 $Y=0.072 $X2=0.891 $Y2=0.0675
cc_78 N_B_M4_g N_C_c_154_n 2.71887e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_79 N_B_c_83_n N_C_c_154_n 4.95866e-19 $X=0.725 $Y=0.072 $X2=0 $Y2=0
cc_80 N_B_M4_g N_C_M3_g 0.00357042f $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_81 N_B_c_76_n N_C_M3_g 2.71887e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_82 N_B_c_83_n N_C_M3_g 4.95866e-19 $X=0.725 $Y=0.072 $X2=0 $Y2=0
cc_83 N_B_c_74_n N_C_c_145_n 0.00150454f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_84 N_B_c_77_n N_C_c_145_n 0.00151103f $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_85 B N_C_c_145_n 4.22126e-19 $X=0.348 $Y=0.133 $X2=0 $Y2=0
cc_86 N_B_c_83_n N_C_c_145_n 0.00162478f $X=0.725 $Y=0.072 $X2=0 $Y2=0
cc_87 N_B_c_85_n N_C_c_145_n 0.00196905f $X=0.547 $Y=0.072 $X2=0 $Y2=0
cc_88 N_B_c_106_p C 4.99572e-19 $X=0.347 $Y=0.1195 $X2=0 $Y2=0
cc_89 N_B_c_86_n C 0.00109049f $X=0.565 $Y=0.072 $X2=0 $Y2=0
cc_90 N_B_c_108_p C 5.1368e-19 $X=0.734 $Y=0.1205 $X2=0 $Y2=0
cc_91 N_B_c_74_n N_6_M11_d 3.5041e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_92 N_B_c_74_n N_6_c_193_n 7.57503e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_93 N_B_c_73_n N_6_c_194_n 2.2196e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_94 N_B_c_71_n N_6_c_195_n 4.61191e-19 $X=0.243 $Y=0.135 $X2=0.945 $Y2=0.135
cc_95 N_B_c_74_n N_6_c_195_n 2.20764e-19 $X=0.351 $Y=0.135 $X2=0.945 $Y2=0.135
cc_96 N_B_c_74_n N_7_M10_s 3.67575e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_97 N_B_c_74_n N_7_c_217_n 0.00203185f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_98 N_B_c_77_n N_7_M20_s 3.67575e-19 $X=0.837 $Y=0.135 $X2=0.891 $Y2=0.2025
cc_99 N_B_c_77_n N_7_c_219_n 0.00203185f $X=0.837 $Y=0.135 $X2=0.945 $Y2=0.135
cc_100 N_B_c_73_n N_7_c_213_n 4.01136e-19 $X=0.297 $Y=0.135 $X2=0.999 $Y2=0.2025
cc_101 N_B_c_74_n N_7_c_213_n 0.00106723f $X=0.351 $Y=0.135 $X2=0.999 $Y2=0.2025
cc_102 N_B_M1_g N_7_c_222_n 3.02555e-19 $X=0.351 $Y=0.0675 $X2=0.999 $Y2=0.2025
cc_103 B N_7_c_222_n 0.00123688f $X=0.348 $Y=0.133 $X2=0.999 $Y2=0.2025
cc_104 N_B_c_85_n N_7_c_214_n 9.87157e-19 $X=0.547 $Y=0.072 $X2=0 $Y2=0
cc_105 N_B_c_83_n N_7_c_225_n 9.87157e-19 $X=0.725 $Y=0.072 $X2=0.894 $Y2=0.081
cc_106 N_B_c_76_n N_7_c_226_n 3.10881e-19 $X=0.783 $Y=0.135 $X2=0.081 $Y2=0.135
cc_107 N_B_M4_g N_7_c_227_n 2.82384e-19 $X=0.729 $Y=0.0675 $X2=0.183 $Y2=0.135
cc_108 N_B_c_126_p N_7_c_227_n 0.0012042f $X=0.734 $Y=0.135 $X2=0.183 $Y2=0.135
cc_109 N_B_c_77_n N_7_c_215_n 0.00105285f $X=0.837 $Y=0.135 $X2=0.183 $Y2=0.135
cc_110 N_B_c_77_n N_8_M19_d 3.44816e-19 $X=0.837 $Y=0.135 $X2=0.081 $Y2=0.135
cc_111 N_B_c_77_n N_8_c_273_n 7.57503e-19 $X=0.837 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_112 N_B_c_76_n N_8_c_274_n 2.65027e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_113 N_B_c_77_n N_8_c_268_n 6.1263e-19 $X=0.837 $Y=0.135 $X2=0.891 $Y2=0.135
cc_114 N_B_c_81_n N_Y_c_303_n 5.88358e-19 $X=0.347 $Y=0.106 $X2=0.894 $Y2=0.078
cc_115 N_B_c_85_n N_Y_c_303_n 0.00186448f $X=0.547 $Y=0.072 $X2=0.894 $Y2=0.078
cc_116 N_B_c_71_n N_Y_c_309_n 4.58673e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_117 N_B_c_74_n N_Y_c_309_n 6.40192e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_118 N_B_c_73_n N_Y_c_331_n 4.62489e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_119 N_B_c_83_n N_Y_c_310_n 0.00218056f $X=0.725 $Y=0.072 $X2=0.183 $Y2=0.135
cc_120 N_B_c_87_n N_Y_c_310_n 5.803e-19 $X=0.734 $Y=0.106 $X2=0.183 $Y2=0.135
cc_121 N_B_M1_g N_Y_c_334_n 2.5731e-19 $X=0.351 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_122 N_B_M4_g N_Y_c_334_n 2.63908e-19 $X=0.729 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_123 N_B_c_84_n N_Y_c_334_n 0.0328697f $X=0.356 $Y=0.072 $X2=0.891 $Y2=0.135
cc_124 N_B_c_76_n N_Y_c_314_n 4.62489e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_125 N_B_c_77_n N_Y_c_314_n 6.30157e-19 $X=0.837 $Y=0.135 $X2=0 $Y2=0
cc_126 N_B_c_77_n N_Y_c_339_n 4.58673e-19 $X=0.837 $Y=0.135 $X2=0.894 $Y2=0.135
cc_127 N_C_c_145_n N_7_M14_s 3.67193e-19 $X=0.675 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_128 N_C_c_145_n N_7_c_231_n 0.00203185f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_129 N_C_c_145_n N_7_M16_s 3.67193e-19 $X=0.675 $Y=0.135 $X2=0.189 $Y2=0.135
cc_130 N_C_c_145_n N_7_c_233_n 0.00203185f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_131 N_C_M2_g N_7_c_214_n 4.98189e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_132 N_C_c_145_n N_7_c_214_n 0.00203644f $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_133 N_C_c_150_n N_7_c_236_n 3.37351e-19 $X=0.459 $Y=0.135 $X2=0.183 $Y2=0.081
cc_134 N_C_c_152_n N_7_c_236_n 4.02808e-19 $X=0.513 $Y=0.135 $X2=0.183 $Y2=0.081
cc_135 C N_7_c_238_n 0.00115485f $X=0.555 $Y=0.133 $X2=0.183 $Y2=0.081
cc_136 N_C_c_153_n N_7_c_225_n 2.3665e-19 $X=0.567 $Y=0.135 $X2=0.894 $Y2=0.081
cc_137 N_C_c_154_n N_7_c_225_n 4.02808e-19 $X=0.621 $Y=0.135 $X2=0.894 $Y2=0.081
cc_138 N_C_c_145_n N_7_c_225_n 0.00140374f $X=0.675 $Y=0.135 $X2=0.894 $Y2=0.081
cc_139 N_C_M3_g N_7_c_242_n 4.23461e-19 $X=0.675 $Y=0.0675 $X2=0.894 $Y2=0.081
cc_140 N_C_M2_g N_Y_c_334_n 2.63908e-19 $X=0.405 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_141 N_C_c_150_n N_Y_c_334_n 2.63908e-19 $X=0.459 $Y=0.135 $X2=0.891 $Y2=0.135
cc_142 N_C_c_152_n N_Y_c_334_n 3.57615e-19 $X=0.513 $Y=0.135 $X2=0.891 $Y2=0.135
cc_143 N_C_c_153_n N_Y_c_334_n 3.57615e-19 $X=0.567 $Y=0.135 $X2=0.891 $Y2=0.135
cc_144 N_C_c_154_n N_Y_c_334_n 2.63908e-19 $X=0.621 $Y=0.135 $X2=0.891 $Y2=0.135
cc_145 N_C_M3_g N_Y_c_334_n 2.63908e-19 $X=0.675 $Y=0.0675 $X2=0.891 $Y2=0.135
cc_146 N_6_c_197_p N_7_c_217_n 0.003312f $X=0.216 $Y=0.2025 $X2=0.081 $Y2=0.2025
cc_147 N_6_c_193_n N_7_c_217_n 0.00352905f $X=0.324 $Y=0.2025 $X2=0.081
+ $Y2=0.2025
cc_148 N_6_c_199_p N_7_c_217_n 0.00250914f $X=0.29 $Y=0.234 $X2=0.081 $Y2=0.2025
cc_149 N_6_c_193_n N_7_c_246_n 0.00317152f $X=0.324 $Y=0.2025 $X2=0.135
+ $Y2=0.2025
cc_150 N_6_c_194_n N_7_c_246_n 4.49606e-19 $X=0.324 $Y=0.234 $X2=0.135
+ $Y2=0.2025
cc_151 N_6_c_197_p N_7_c_213_n 4.51268e-19 $X=0.216 $Y=0.2025 $X2=0.999
+ $Y2=0.2025
cc_152 N_6_c_193_n N_7_c_213_n 0.00233206f $X=0.324 $Y=0.2025 $X2=0.999
+ $Y2=0.2025
cc_153 N_6_c_199_p N_7_c_213_n 0.00704495f $X=0.29 $Y=0.234 $X2=0.999 $Y2=0.2025
cc_154 N_6_c_187_n N_Y_c_346_n 0.00337028f $X=0.108 $Y=0.2025 $X2=0.891
+ $Y2=0.135
cc_155 N_6_c_188_n N_Y_c_346_n 3.09693e-19 $X=0.176 $Y=0.234 $X2=0.891 $Y2=0.135
cc_156 N_6_c_187_n N_Y_c_293_n 0.00352892f $X=0.108 $Y=0.2025 $X2=0.945
+ $Y2=0.135
cc_157 N_6_c_197_p N_Y_c_293_n 0.00332044f $X=0.216 $Y=0.2025 $X2=0.945
+ $Y2=0.135
cc_158 N_6_c_188_n N_Y_c_293_n 0.00250914f $X=0.176 $Y=0.234 $X2=0.945 $Y2=0.135
cc_159 N_6_c_197_p N_Y_c_318_n 4.48103e-19 $X=0.216 $Y=0.2025 $X2=0.894
+ $Y2=0.135
cc_160 N_6_c_187_n N_Y_c_352_n 0.00233206f $X=0.108 $Y=0.2025 $X2=0 $Y2=0
cc_161 N_6_c_188_n N_Y_c_352_n 0.00702934f $X=0.176 $Y=0.234 $X2=0 $Y2=0
cc_162 N_7_c_251_p N_8_c_273_n 0.00317169f $X=0.702 $Y=0.2025 $X2=0.081
+ $Y2=0.2025
cc_163 N_7_c_219_n N_8_c_273_n 0.00352901f $X=0.81 $Y=0.2025 $X2=0.081
+ $Y2=0.2025
cc_164 N_7_c_215_n N_8_c_273_n 0.00233206f $X=0.7765 $Y=0.198 $X2=0.081
+ $Y2=0.2025
cc_165 N_7_c_219_n N_8_c_279_n 0.00328787f $X=0.81 $Y=0.2025 $X2=0.135
+ $Y2=0.2025
cc_166 N_7_c_226_n N_8_c_279_n 4.51268e-19 $X=0.81 $Y=0.198 $X2=0.135 $Y2=0.2025
cc_167 N_7_c_251_p N_8_c_274_n 4.49606e-19 $X=0.702 $Y=0.2025 $X2=0 $Y2=0
cc_168 N_7_c_219_n N_8_c_274_n 0.00250914f $X=0.81 $Y=0.2025 $X2=0 $Y2=0
cc_169 N_7_c_215_n N_8_c_274_n 0.00697856f $X=0.7765 $Y=0.198 $X2=0 $Y2=0
cc_170 N_7_c_246_n N_Y_c_303_n 0.00158656f $X=0.378 $Y=0.2025 $X2=0.894
+ $Y2=0.078
cc_171 N_7_c_213_n N_Y_c_331_n 4.01913e-19 $X=0.338 $Y=0.198 $X2=0.081 $Y2=0.135
cc_172 N_7_c_251_p N_Y_c_310_n 0.0015999f $X=0.702 $Y=0.2025 $X2=0.183 $Y2=0.135
cc_173 N_7_c_214_n N_Y_c_334_n 4.01913e-19 $X=0.418 $Y=0.198 $X2=0.891 $Y2=0.135
cc_174 N_7_c_215_n N_Y_c_314_n 4.01913e-19 $X=0.7765 $Y=0.198 $X2=0 $Y2=0
cc_175 N_7_c_213_n N_Y_c_318_n 3.18557e-19 $X=0.338 $Y=0.198 $X2=0.894 $Y2=0.135
cc_176 N_7_c_226_n N_Y_c_321_n 3.18557e-19 $X=0.81 $Y=0.198 $X2=0 $Y2=0
cc_177 N_8_c_279_n N_Y_c_295_n 0.00328789f $X=0.864 $Y=0.2025 $X2=0.999
+ $Y2=0.135
cc_178 N_8_c_267_n N_Y_c_295_n 0.00350515f $X=0.972 $Y=0.2025 $X2=0.999
+ $Y2=0.135
cc_179 N_8_c_269_n N_Y_c_295_n 0.00249187f $X=0.972 $Y=0.234 $X2=0.999 $Y2=0.135
cc_180 N_8_c_267_n N_Y_c_364_n 0.00337028f $X=0.972 $Y=0.2025 $X2=0.999
+ $Y2=0.2025
cc_181 N_8_c_269_n N_Y_c_364_n 3.09693e-19 $X=0.972 $Y=0.234 $X2=0.999
+ $Y2=0.2025
cc_182 N_8_c_279_n N_Y_c_321_n 4.48103e-19 $X=0.864 $Y=0.2025 $X2=0 $Y2=0
cc_183 N_8_c_267_n N_Y_c_321_n 0.00233206f $X=0.972 $Y=0.2025 $X2=0 $Y2=0
cc_184 N_8_c_269_n N_Y_c_321_n 0.00704501f $X=0.972 $Y=0.234 $X2=0 $Y2=0

* END of "./NOR3x2_ASAP7_75t_R.pex.sp.NOR3X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR3xp33_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:45:04 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR3xp33_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR3xp33_ASAP7_75t_R.pex.sp.pex"
* File: NOR3xp33_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:45:04 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR3XP33_ASAP7_75T_R%A 2 5 7 10 VSS
c9 10 VSS 0.00149021f $X=0.083 $Y=0.133
c10 5 VSS 0.0016745f $X=0.081 $Y=0.135
c11 2 VSS 0.0649376f $X=0.081 $Y=0.054
r12 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r14 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NOR3XP33_ASAP7_75T_R%B 2 5 7 11 VSS
c12 11 VSS 0.00596567f $X=0.136 $Y=0.133
c13 5 VSS 0.00116826f $X=0.135 $Y=0.135
c14 2 VSS 0.0601197f $X=0.135 $Y=0.054
r15 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r17 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_NOR3XP33_ASAP7_75T_R%C 2 7 11 14 VSS
c5 14 VSS 0.00522154f $X=0.2 $Y=0.135
c6 11 VSS 0.0144657f $X=0.202 $Y=0.133
c7 2 VSS 0.0639038f $X=0.189 $Y=0.054
r8 11 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.2 $Y=0.135 $X2=0.2
+ $Y2=0.135
r9 5 14 11 $w=2e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.189 $Y=0.135
+ $X2=0.2 $Y2=0.135
r10 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r11 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_NOR3XP33_ASAP7_75T_R%Y 1 4 6 7 10 11 14 19 21 33 35 42 VSS
c11 45 VSS 9.40634e-19 $X=0.045 $Y=0.234
c12 44 VSS 0.0032947f $X=0.036 $Y=0.234
c13 42 VSS 0.00287833f $X=0.054 $Y=0.234
c14 36 VSS 0.00103857f $X=0.153 $Y=0.036
c15 35 VSS 0.00142296f $X=0.144 $Y=0.036
c16 34 VSS 0.00632432f $X=0.126 $Y=0.036
c17 33 VSS 0.00142296f $X=0.09 $Y=0.036
c18 32 VSS 4.19006e-19 $X=0.072 $Y=0.036
c19 31 VSS 0.00321919f $X=0.068 $Y=0.036
c20 29 VSS 0.00358469f $X=0.162 $Y=0.036
c21 24 VSS 0.00335462f $X=0.036 $Y=0.036
c22 23 VSS 5.62956e-19 $X=0.027 $Y=0.2125
c23 21 VSS 0.00125275f $X=0.027 $Y=0.0985
c24 20 VSS 8.11244e-19 $X=0.027 $Y=0.07
c25 19 VSS 0.00448957f $X=0.028 $Y=0.127
c26 17 VSS 5.45722e-19 $X=0.027 $Y=0.225
c27 14 VSS 0.00224295f $X=0.056 $Y=0.2025
c28 11 VSS 3.02808e-19 $X=0.071 $Y=0.2025
c29 10 VSS 0.0075021f $X=0.162 $Y=0.054
c30 6 VSS 5.65078e-19 $X=0.179 $Y=0.054
c31 4 VSS 0.00549622f $X=0.056 $Y=0.054
c32 1 VSS 2.53241e-19 $X=0.071 $Y=0.054
r33 44 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.045 $Y2=0.234
r34 42 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.045 $Y2=0.234
r35 39 44 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.036 $Y2=0.234
r36 35 36 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.153 $Y2=0.036
r37 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r38 33 34 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.126 $Y2=0.036
r39 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r40 31 32 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.068
+ $Y=0.036 $X2=0.072 $Y2=0.036
r41 29 36 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.153 $Y2=0.036
r42 26 31 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.068 $Y2=0.036
r43 24 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.054 $Y2=0.036
r44 22 23 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.2 $X2=0.027 $Y2=0.2125
r45 20 21 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.0985
r46 19 22 4.95679 $w=1.8e-08 $l=7.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.127 $X2=0.027 $Y2=0.2
r47 19 21 1.93519 $w=1.8e-08 $l=2.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.127 $X2=0.027 $Y2=0.0985
r48 17 39 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.234
r49 17 23 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.2125
r50 16 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r51 16 20 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r52 14 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r53 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r54 10 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r55 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.162 $Y2=0.054
r56 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.054 $X2=0.162 $Y2=0.054
r57 4 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r58 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.054 $X2=0.056 $Y2=0.054
.ends

.subckt PM_NOR3XP33_ASAP7_75T_R%7 1 2 VSS
c0 1 VSS 0.00221026f $X=0.125 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends

.subckt PM_NOR3XP33_ASAP7_75T_R%8 1 2 VSS
c1 1 VSS 0.00199907f $X=0.179 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends


* END of "./NOR3xp33_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR3xp33_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 VSS N_A_M0_g N_Y_M0_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_B_M1_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_C_M2_g N_Y_M2_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 N_7_M3_d N_A_M3_g N_Y_M3_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M4 N_8_M4_d N_B_M4_g N_7_M4_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M5 VDD N_C_M5_g N_8_M5_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
*
* 
* .include "NOR3xp33_ASAP7_75t_R.pex.sp.NOR3XP33_ASAP7_75T_R.pxi"
* BEGIN of "./NOR3xp33_ASAP7_75t_R.pex.sp.NOR3XP33_ASAP7_75T_R.pxi"
* File: NOR3xp33_ASAP7_75t_R.pex.sp.NOR3XP33_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:45:04 2017
* 
x_PM_NOR3XP33_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M3_g A VSS
+ PM_NOR3XP33_ASAP7_75T_R%A
x_PM_NOR3XP33_ASAP7_75T_R%B N_B_M1_g N_B_c_11_n N_B_M4_g B VSS
+ PM_NOR3XP33_ASAP7_75T_R%B
x_PM_NOR3XP33_ASAP7_75T_R%C N_C_M2_g N_C_M5_g C N_C_c_25_n VSS
+ PM_NOR3XP33_ASAP7_75T_R%C
x_PM_NOR3XP33_ASAP7_75T_R%Y N_Y_M0_s N_Y_c_27_n N_Y_M2_s N_Y_M1_d N_Y_c_32_n
+ N_Y_M3_s N_Y_c_28_n Y N_Y_c_29_n N_Y_c_30_n N_Y_c_34_n N_Y_c_36_n VSS
+ PM_NOR3XP33_ASAP7_75T_R%Y
x_PM_NOR3XP33_ASAP7_75T_R%7 N_7_M4_s N_7_M3_d VSS PM_NOR3XP33_ASAP7_75T_R%7
x_PM_NOR3XP33_ASAP7_75T_R%8 N_8_M5_s N_8_M4_d VSS PM_NOR3XP33_ASAP7_75T_R%8
cc_1 N_A_M0_g N_B_M1_g 0.00327995f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A_c_2_p N_B_c_11_n 8.52536e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A B 0.00618453f $X=0.083 $Y=0.133 $X2=0.136 $Y2=0.133
cc_4 N_A_M0_g N_C_M2_g 2.66145e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 A N_Y_c_27_n 3.31541e-19 $X=0.083 $Y=0.133 $X2=0.135 $Y2=0.135
cc_6 A N_Y_c_28_n 0.0013295f $X=0.083 $Y=0.133 $X2=0.135 $Y2=0.135
cc_7 A N_Y_c_29_n 0.00547852f $X=0.083 $Y=0.133 $X2=0 $Y2=0
cc_8 N_A_M0_g N_Y_c_30_n 2.57255e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_9 A N_Y_c_30_n 0.00123619f $X=0.083 $Y=0.133 $X2=0 $Y2=0
cc_10 N_B_M1_g N_C_M2_g 0.00344695f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_11 B C 0.00690454f $X=0.136 $Y=0.133 $X2=0 $Y2=0
cc_12 N_B_c_11_n N_C_c_25_n 9.17588e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_13 B N_Y_c_32_n 3.55402e-19 $X=0.136 $Y=0.133 $X2=0.083 $Y2=0.133
cc_14 B N_Y_c_28_n 6.83303e-19 $X=0.136 $Y=0.133 $X2=0 $Y2=0
cc_15 N_B_M1_g N_Y_c_34_n 2.57255e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_16 B N_Y_c_34_n 0.00123985f $X=0.136 $Y=0.133 $X2=0 $Y2=0
cc_17 B N_Y_c_36_n 7.1001e-19 $X=0.136 $Y=0.133 $X2=0 $Y2=0
cc_18 B N_8_M5_s 3.84149e-19 $X=0.136 $Y=0.133 $X2=0.081 $Y2=0.054
cc_19 C N_Y_c_32_n 2.68871e-19 $X=0.202 $Y=0.133 $X2=0.083 $Y2=0.133

* END of "./NOR3xp33_ASAP7_75t_R.pex.sp.NOR3XP33_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR4xp25_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:45:27 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR4xp25_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR4xp25_ASAP7_75t_R.pex.sp.pex"
* File: NOR4xp25_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:45:27 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR4XP25_ASAP7_75T_R%D 2 5 7 15 VSS
c8 15 VSS 0.022281f $X=0.081 $Y=0.132
c9 5 VSS 0.00296916f $X=0.081 $Y=0.135
c10 2 VSS 0.0646435f $X=0.081 $Y=0.054
r11 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r12 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r13 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NOR4XP25_ASAP7_75T_R%C 2 5 7 10 VSS
c10 10 VSS 0.00301312f $X=0.135 $Y=0.132
c11 5 VSS 0.00183837f $X=0.135 $Y=0.135
c12 2 VSS 0.0597098f $X=0.135 $Y=0.054
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r15 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_NOR4XP25_ASAP7_75T_R%B 2 5 7 10 VSS
c13 10 VSS 0.00210298f $X=0.189 $Y=0.132
c14 5 VSS 0.00106871f $X=0.189 $Y=0.135
c15 2 VSS 0.0600389f $X=0.189 $Y=0.054
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
.ends

.subckt PM_NOR4XP25_ASAP7_75T_R%A 2 5 7 10 VSS
c9 10 VSS 0.00165342f $X=0.243 $Y=0.132
c10 5 VSS 0.00225849f $X=0.243 $Y=0.135
c11 2 VSS 0.0653596f $X=0.243 $Y=0.054
r12 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r14 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_NOR4XP25_ASAP7_75T_R%Y 1 4 6 7 10 11 14 16 19 29 30 32 37 39 45 49 55
+ VSS
c18 55 VSS 0.00396291f $X=0.288 $Y=0.234
c19 54 VSS 0.00278493f $X=0.297 $Y=0.234
c20 49 VSS 4.30865e-19 $X=0.297 $Y=0.2125
c21 47 VSS 2.31784e-19 $X=0.297 $Y=0.07
c22 46 VSS 5.7946e-19 $X=0.297 $Y=0.063
c23 45 VSS 0.00568545f $X=0.297 $Y=0.124
c24 43 VSS 8.62726e-19 $X=0.297 $Y=0.225
c25 41 VSS 6.8347e-19 $X=0.263 $Y=0.036
c26 40 VSS 3.38363e-19 $X=0.256 $Y=0.036
c27 39 VSS 0.00146362f $X=0.252 $Y=0.036
c28 38 VSS 0.00631478f $X=0.234 $Y=0.036
c29 37 VSS 0.00146362f $X=0.198 $Y=0.036
c30 36 VSS 0.00377397f $X=0.18 $Y=0.036
c31 32 VSS 0.00146362f $X=0.144 $Y=0.036
c32 31 VSS 0.00575705f $X=0.126 $Y=0.036
c33 30 VSS 0.00322775f $X=0.095 $Y=0.036
c34 29 VSS 0.0024767f $X=0.057 $Y=0.036
c35 21 VSS 0.00591782f $X=0.288 $Y=0.036
c36 19 VSS 0.00261811f $X=0.268 $Y=0.2025
c37 14 VSS 0.00574816f $X=0.268 $Y=0.054
c38 10 VSS 0.0079209f $X=0.162 $Y=0.054
c39 6 VSS 5.3314e-19 $X=0.179 $Y=0.054
c40 4 VSS 0.0058471f $X=0.056 $Y=0.054
c41 1 VSS 4.80622e-19 $X=0.071 $Y=0.054
r42 55 56 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.2925 $Y2=0.234
r43 54 56 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.234 $X2=0.2925 $Y2=0.234
r44 51 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.288 $Y2=0.234
r45 48 49 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.2 $X2=0.297 $Y2=0.2125
r46 46 47 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.063 $X2=0.297 $Y2=0.07
r47 45 48 5.16049 $w=1.8e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.124 $X2=0.297 $Y2=0.2
r48 45 47 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.124 $X2=0.297 $Y2=0.07
r49 43 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.234
r50 43 49 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.2125
r51 42 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.063
r52 40 41 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.036 $X2=0.263 $Y2=0.036
r53 39 40 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.256 $Y2=0.036
r54 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r55 37 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.234 $Y2=0.036
r56 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r57 34 41 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.263 $Y2=0.036
r58 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r59 30 31 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.036 $X2=0.126 $Y2=0.036
r60 29 30 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.057
+ $Y=0.036 $X2=0.095 $Y2=0.036
r61 27 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r62 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.144 $Y2=0.036
r63 23 29 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.057 $Y2=0.036
r64 21 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r65 21 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.27 $Y2=0.036
r66 19 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r67 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.268 $Y2=0.2025
r68 14 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r69 11 14 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.054 $X2=0.268 $Y2=0.054
r70 10 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r71 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.162 $Y2=0.054
r72 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.054 $X2=0.162 $Y2=0.054
r73 4 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r74 1 4 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.054 $X2=0.056 $Y2=0.054
.ends

.subckt PM_NOR4XP25_ASAP7_75T_R%8 1 2 VSS
c0 1 VSS 0.00233476f $X=0.125 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends

.subckt PM_NOR4XP25_ASAP7_75T_R%9 1 2 VSS
c0 1 VSS 0.00228146f $X=0.179 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends

.subckt PM_NOR4XP25_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00228146f $X=0.233 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.199 $Y2=0.2025
.ends


* END of "./NOR4xp25_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR4xp25_ASAP7_75t_R  VSS VDD D C B A Y
* 
* Y	Y
* A	A
* B	B
* C	C
* D	D
M0 VSS N_D_M0_g N_Y_M0_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_C_M1_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_B_M2_g N_Y_M2_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_A_M3_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 N_8_M4_d N_D_M4_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M5 N_9_M5_d N_C_M5_g N_8_M5_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 N_10_M6_d N_B_M6_g N_9_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M7 N_Y_M7_d N_A_M7_g N_10_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
*
* 
* .include "NOR4xp25_ASAP7_75t_R.pex.sp.NOR4XP25_ASAP7_75T_R.pxi"
* BEGIN of "./NOR4xp25_ASAP7_75t_R.pex.sp.NOR4XP25_ASAP7_75T_R.pxi"
* File: NOR4xp25_ASAP7_75t_R.pex.sp.NOR4XP25_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:45:27 2017
* 
x_PM_NOR4XP25_ASAP7_75T_R%D N_D_M0_g N_D_c_2_p N_D_M4_g D VSS
+ PM_NOR4XP25_ASAP7_75T_R%D
x_PM_NOR4XP25_ASAP7_75T_R%C N_C_M1_g N_C_c_10_n N_C_M5_g C VSS
+ PM_NOR4XP25_ASAP7_75T_R%C
x_PM_NOR4XP25_ASAP7_75T_R%B N_B_M2_g N_B_c_21_n N_B_M6_g B VSS
+ PM_NOR4XP25_ASAP7_75T_R%B
x_PM_NOR4XP25_ASAP7_75T_R%A N_A_M3_g N_A_c_34_n N_A_M7_g A VSS
+ PM_NOR4XP25_ASAP7_75T_R%A
x_PM_NOR4XP25_ASAP7_75T_R%Y N_Y_M0_s N_Y_c_41_n N_Y_M2_s N_Y_M1_d N_Y_c_45_n
+ N_Y_M3_d N_Y_c_54_n N_Y_M7_d N_Y_c_49_n N_Y_c_42_n N_Y_c_43_n N_Y_c_46_n
+ N_Y_c_50_n N_Y_c_56_n Y N_Y_c_52_n N_Y_c_53_n VSS PM_NOR4XP25_ASAP7_75T_R%Y
x_PM_NOR4XP25_ASAP7_75T_R%8 N_8_M5_s N_8_M4_d VSS PM_NOR4XP25_ASAP7_75T_R%8
x_PM_NOR4XP25_ASAP7_75T_R%9 N_9_M6_s N_9_M5_d VSS PM_NOR4XP25_ASAP7_75T_R%9
x_PM_NOR4XP25_ASAP7_75T_R%10 N_10_M7_s N_10_M6_d VSS PM_NOR4XP25_ASAP7_75T_R%10
cc_1 N_D_M0_g N_C_M1_g 0.0032073f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_D_c_2_p N_C_c_10_n 0.00101358f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 D C 0.00294793f $X=0.081 $Y=0.132 $X2=0.135 $Y2=0.132
cc_4 N_D_M0_g N_B_M2_g 2.66145e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 D N_Y_c_41_n 0.00208467f $X=0.081 $Y=0.132 $X2=0.135 $Y2=0.135
cc_6 D N_Y_c_42_n 0.00194715f $X=0.081 $Y=0.132 $X2=0 $Y2=0
cc_7 N_D_M0_g N_Y_c_43_n 4.31632e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_8 D N_Y_c_43_n 3.65373e-19 $X=0.081 $Y=0.132 $X2=0 $Y2=0
cc_9 N_C_M1_g N_B_M2_g 0.0035196f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_10 N_C_c_10_n N_B_c_21_n 7.51247e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_11 C B 0.00814915f $X=0.135 $Y=0.132 $X2=0 $Y2=0
cc_12 N_C_M1_g N_A_M3_g 2.71887e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_13 C N_Y_c_45_n 3.24828e-19 $X=0.135 $Y=0.132 $X2=0 $Y2=0
cc_14 N_C_M1_g N_Y_c_46_n 2.64924e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_15 C N_Y_c_46_n 0.00125705f $X=0.135 $Y=0.132 $X2=0 $Y2=0
cc_16 N_B_M2_g N_A_M3_g 0.00333077f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_17 N_B_c_21_n N_A_c_34_n 7.51046e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_18 B A 0.00620922f $X=0.189 $Y=0.132 $X2=0 $Y2=0
cc_19 B N_Y_c_45_n 3.31541e-19 $X=0.189 $Y=0.132 $X2=0 $Y2=0
cc_20 B N_Y_c_49_n 4.68998e-19 $X=0.189 $Y=0.132 $X2=0.081 $Y2=0.135
cc_21 N_B_M2_g N_Y_c_50_n 2.64606e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_22 B N_Y_c_50_n 0.0012569f $X=0.189 $Y=0.132 $X2=0 $Y2=0
cc_23 B N_Y_c_52_n 2.69891e-19 $X=0.189 $Y=0.132 $X2=0 $Y2=0
cc_24 B N_Y_c_53_n 4.44922e-19 $X=0.189 $Y=0.132 $X2=0 $Y2=0
cc_25 A N_Y_c_54_n 3.31541e-19 $X=0.243 $Y=0.132 $X2=0.135 $Y2=0.135
cc_26 A N_Y_c_49_n 0.0013295f $X=0.243 $Y=0.132 $X2=0 $Y2=0
cc_27 N_A_M3_g N_Y_c_56_n 2.64924e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_28 A N_Y_c_56_n 0.00125383f $X=0.243 $Y=0.132 $X2=0 $Y2=0
cc_29 A Y 0.00549499f $X=0.243 $Y=0.132 $X2=0 $Y2=0

* END of "./NOR4xp25_ASAP7_75t_R.pex.sp.NOR4XP25_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR4xp75_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:45:49 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR4xp75_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR4xp75_ASAP7_75t_R.pex.sp.pex"
* File: NOR4xp75_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:45:49 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR4XP75_ASAP7_75T_R%D 2 7 10 15 18 21 23 41 VSS
c16 41 VSS 0.0313986f $X=0.081 $Y=0.138
c17 21 VSS 0.0109493f $X=0.189 $Y=0.135
c18 18 VSS 0.0622597f $X=0.189 $Y=0.054
c19 10 VSS 0.0638991f $X=0.135 $Y=0.054
c20 2 VSS 0.0646334f $X=0.081 $Y=0.054
r21 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r22 18 21 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.135
r23 13 21 60 $w=1.8e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135 $Y=0.135
+ $X2=0.189 $Y2=0.135
r24 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r25 10 13 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
r26 5 13 60 $w=1.8e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081 $Y=0.135
+ $X2=0.135 $Y2=0.135
r27 5 41 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r28 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r29 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_NOR4XP75_ASAP7_75T_R%C 2 7 10 15 18 21 23 33 VSS
c35 33 VSS 0.00488597f $X=0.3 $Y=0.138
c36 21 VSS 0.00619913f $X=0.351 $Y=0.135
c37 18 VSS 0.0624063f $X=0.351 $Y=0.054
c38 10 VSS 0.0636165f $X=0.297 $Y=0.054
c39 2 VSS 0.0620301f $X=0.243 $Y=0.054
r40 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r41 18 21 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.054 $X2=0.351 $Y2=0.135
r42 13 21 60 $w=1.8e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297 $Y=0.135
+ $X2=0.351 $Y2=0.135
r43 13 33 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r44 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r45 10 13 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.135
r46 5 13 60 $w=1.8e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243 $Y=0.135
+ $X2=0.297 $Y2=0.135
r47 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r48 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
.ends

.subckt PM_NOR4XP75_ASAP7_75T_R%B 2 7 10 15 18 21 23 30 VSS
c34 30 VSS 0.00265592f $X=0.521 $Y=0.138
c35 21 VSS 0.00647082f $X=0.513 $Y=0.135
c36 18 VSS 0.0621861f $X=0.513 $Y=0.054
c37 10 VSS 0.0640813f $X=0.459 $Y=0.054
c38 2 VSS 0.0623945f $X=0.405 $Y=0.054
r39 21 30 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r40 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r41 18 21 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.054 $X2=0.513 $Y2=0.135
r42 13 21 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459 $Y=0.135
+ $X2=0.513 $Y2=0.135
r43 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r44 10 13 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.054 $X2=0.459 $Y2=0.135
r45 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405 $Y=0.135
+ $X2=0.459 $Y2=0.135
r46 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r47 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.054 $X2=0.405 $Y2=0.135
.ends

.subckt PM_NOR4XP75_ASAP7_75T_R%A 2 7 10 15 18 21 23 29 VSS
c27 29 VSS 0.00150073f $X=0.621 $Y=0.138
c28 21 VSS 0.00700146f $X=0.675 $Y=0.135
c29 18 VSS 0.066303f $X=0.675 $Y=0.054
c30 10 VSS 0.0636276f $X=0.621 $Y=0.054
c31 2 VSS 0.0627233f $X=0.567 $Y=0.054
r32 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.2025
r33 18 21 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.054 $X2=0.675 $Y2=0.135
r34 13 21 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621 $Y=0.135
+ $X2=0.675 $Y2=0.135
r35 13 29 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r36 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r37 10 13 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.054 $X2=0.621 $Y2=0.135
r38 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.567 $Y=0.135
+ $X2=0.621 $Y2=0.135
r39 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r40 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.054 $X2=0.567 $Y2=0.135
.ends

.subckt PM_NOR4XP75_ASAP7_75T_R%7 1 2 5 6 7 10 11 12 15 17 25 26 28 31 VSS
c28 31 VSS 0.0024855f $X=0.256 $Y=0.234
c29 30 VSS 9.70579e-19 $X=0.225 $Y=0.234
c30 28 VSS 0.00708487f $X=0.324 $Y=0.234
c31 26 VSS 3.3597e-19 $X=0.2115 $Y=0.234
c32 25 VSS 0.0118841f $X=0.207 $Y=0.234
c33 17 VSS 0.00160315f $X=0.108 $Y=0.234
c34 15 VSS 0.00283956f $X=0.324 $Y=0.2025
c35 11 VSS 6.1922e-19 $X=0.341 $Y=0.2025
c36 10 VSS 0.00618448f $X=0.216 $Y=0.2025
c37 6 VSS 6.20841e-19 $X=0.233 $Y=0.2025
c38 5 VSS 0.00903596f $X=0.108 $Y=0.2025
c39 1 VSS 5.24403e-19 $X=0.125 $Y=0.2025
r40 30 31 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.234 $X2=0.256 $Y2=0.234
r41 28 31 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.256 $Y2=0.234
r42 25 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.234 $X2=0.2115 $Y2=0.234
r43 23 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.225 $Y2=0.234
r44 23 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.2115 $Y2=0.234
r45 17 25 6.72222 $w=1.8e-08 $l=9.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.207 $Y2=0.234
r46 15 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r47 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r48 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r49 10 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r50 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r51 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r52 5 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r53 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.2025 $X2=0.108 $Y2=0.2025
r54 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.108 $Y2=0.2025
.ends

.subckt PM_NOR4XP75_ASAP7_75T_R%8 1 2 5 6 7 10 11 12 15 23 24 26 28 29 VSS
c31 29 VSS 3.56711e-19 $X=0.4485 $Y=0.198
c32 28 VSS 0.00305582f $X=0.412 $Y=0.198
c33 26 VSS 4.07927e-19 $X=0.485 $Y=0.198
c34 24 VSS 3.19402e-19 $X=0.34 $Y=0.198
c35 23 VSS 8.46035e-21 $X=0.306 $Y=0.198
c36 15 VSS 0.00387497f $X=0.486 $Y=0.2025
c37 11 VSS 5.71502e-19 $X=0.503 $Y=0.2025
c38 10 VSS 0.00180298f $X=0.378 $Y=0.2025
c39 6 VSS 7.40637e-19 $X=0.395 $Y=0.2025
c40 5 VSS 0.00353193f $X=0.27 $Y=0.2025
c41 1 VSS 6.21322e-19 $X=0.287 $Y=0.2025
r42 28 29 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.412
+ $Y=0.198 $X2=0.4485 $Y2=0.198
r43 26 29 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.485
+ $Y=0.198 $X2=0.4485 $Y2=0.198
r44 23 24 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.198 $X2=0.34 $Y2=0.198
r45 21 28 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.198 $X2=0.412 $Y2=0.198
r46 21 24 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.198 $X2=0.34 $Y2=0.198
r47 17 23 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.198 $X2=0.306 $Y2=0.198
r48 15 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.485 $Y=0.198 $X2=0.485
+ $Y2=0.198
r49 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.486 $Y2=0.2025
r50 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.2025 $X2=0.486 $Y2=0.2025
r51 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.198 $X2=0.378
+ $Y2=0.198
r52 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r53 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r54 5 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.198 $X2=0.27
+ $Y2=0.198
r55 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.2025 $X2=0.27 $Y2=0.2025
r56 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.27 $Y2=0.2025
.ends

.subckt PM_NOR4XP75_ASAP7_75T_R%9 1 2 5 6 7 10 11 12 15 23 25 26 28 31 VSS
c33 31 VSS 0.00288066f $X=0.58 $Y=0.234
c34 30 VSS 9.70579e-19 $X=0.549 $Y=0.234
c35 28 VSS 0.00738141f $X=0.648 $Y=0.234
c36 26 VSS 3.3597e-19 $X=0.5355 $Y=0.234
c37 25 VSS 0.00212432f $X=0.531 $Y=0.234
c38 24 VSS 6.07508e-19 $X=0.504 $Y=0.234
c39 23 VSS 0.00739746f $X=0.499 $Y=0.234
c40 15 VSS 0.00276854f $X=0.648 $Y=0.2025
c41 11 VSS 6.30433e-19 $X=0.665 $Y=0.2025
c42 10 VSS 0.00216821f $X=0.54 $Y=0.2025
c43 6 VSS 6.20841e-19 $X=0.557 $Y=0.2025
c44 5 VSS 0.00283848f $X=0.432 $Y=0.2025
c45 1 VSS 6.25349e-19 $X=0.449 $Y=0.2025
r46 30 31 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.549
+ $Y=0.234 $X2=0.58 $Y2=0.234
r47 28 31 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.58 $Y2=0.234
r48 25 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.531
+ $Y=0.234 $X2=0.5355 $Y2=0.234
r49 24 25 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.531 $Y2=0.234
r50 23 24 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.499
+ $Y=0.234 $X2=0.504 $Y2=0.234
r51 21 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.549 $Y2=0.234
r52 21 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.5355 $Y2=0.234
r53 17 23 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.499 $Y2=0.234
r54 15 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234 $X2=0.648
+ $Y2=0.234
r55 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.648 $Y2=0.2025
r56 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.648 $Y2=0.2025
r57 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r58 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r59 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r60 5 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r61 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.2025 $X2=0.432 $Y2=0.2025
r62 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.449
+ $Y=0.2025 $X2=0.432 $Y2=0.2025
.ends

.subckt PM_NOR4XP75_ASAP7_75T_R%Y 1 2 5 6 7 10 11 12 15 16 17 20 21 22 25 26 27
+ 30 31 32 35 36 39 41 43 51 52 56 57 64 66 67 72 74 83 84 85 86 90 92 VSS
c58 94 VSS 5.54434e-19 $X=0.729 $Y=0.1765
c59 92 VSS 0.00205494f $X=0.729 $Y=0.108
c60 91 VSS 0.00131846f $X=0.729 $Y=0.07
c61 90 VSS 0.00288705f $X=0.732 $Y=0.146
c62 88 VSS 6.07272e-19 $X=0.729 $Y=0.189
c63 86 VSS 6.39993e-19 $X=0.6845 $Y=0.198
c64 85 VSS 3.43772e-19 $X=0.666 $Y=0.198
c65 84 VSS 8.46035e-21 $X=0.63 $Y=0.198
c66 83 VSS 3.77963e-19 $X=0.612 $Y=0.198
c67 75 VSS 0.00367873f $X=0.72 $Y=0.198
c68 74 VSS 0.00146362f $X=0.63 $Y=0.036
c69 73 VSS 0.00501797f $X=0.612 $Y=0.036
c70 72 VSS 0.00285554f $X=0.58 $Y=0.036
c71 71 VSS 0.00172044f $X=0.549 $Y=0.036
c72 67 VSS 8.32314e-19 $X=0.531 $Y=0.036
c73 66 VSS 0.00142296f $X=0.522 $Y=0.036
c74 65 VSS 5.34627e-19 $X=0.504 $Y=0.036
c75 64 VSS 0.0214141f $X=0.499 $Y=0.036
c76 57 VSS 0.00146362f $X=0.306 $Y=0.036
c77 56 VSS 0.00900134f $X=0.288 $Y=0.036
c78 52 VSS 4.42399e-19 $X=0.2115 $Y=0.036
c79 51 VSS 0.0117964f $X=0.207 $Y=0.036
c80 43 VSS 0.00128823f $X=0.108 $Y=0.036
c81 41 VSS 0.0134649f $X=0.72 $Y=0.036
c82 39 VSS 0.00220041f $X=0.7 $Y=0.2025
c83 35 VSS 0.00395433f $X=0.594 $Y=0.2025
c84 31 VSS 5.7545e-19 $X=0.611 $Y=0.2025
c85 30 VSS 0.00824104f $X=0.648 $Y=0.054
c86 26 VSS 5.3314e-19 $X=0.665 $Y=0.054
c87 25 VSS 0.00775062f $X=0.54 $Y=0.054
c88 21 VSS 5.3314e-19 $X=0.557 $Y=0.054
c89 20 VSS 0.00774743f $X=0.432 $Y=0.054
c90 16 VSS 5.3314e-19 $X=0.449 $Y=0.054
c91 15 VSS 0.00820645f $X=0.324 $Y=0.054
c92 11 VSS 5.3314e-19 $X=0.341 $Y=0.054
c93 10 VSS 0.0073284f $X=0.216 $Y=0.054
c94 6 VSS 5.3314e-19 $X=0.233 $Y=0.054
c95 5 VSS 0.00750643f $X=0.108 $Y=0.054
c96 1 VSS 5.5175e-19 $X=0.125 $Y=0.054
r97 93 94 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.164 $X2=0.729 $Y2=0.1765
r98 91 92 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.07 $X2=0.729 $Y2=0.108
r99 90 93 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.146 $X2=0.729 $Y2=0.164
r100 90 92 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.146 $X2=0.729 $Y2=0.108
r101 88 94 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.189 $X2=0.729 $Y2=0.1765
r102 87 91 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.729
+ $Y=0.045 $X2=0.729 $Y2=0.07
r103 85 86 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.666
+ $Y=0.198 $X2=0.6845 $Y2=0.198
r104 84 85 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.198 $X2=0.666 $Y2=0.198
r105 83 84 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.198 $X2=0.63 $Y2=0.198
r106 81 86 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.703
+ $Y=0.198 $X2=0.6845 $Y2=0.198
r107 77 83 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.198 $X2=0.612 $Y2=0.198
r108 75 88 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.198 $X2=0.729 $Y2=0.189
r109 75 81 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.198 $X2=0.703 $Y2=0.198
r110 73 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.63 $Y2=0.036
r111 72 73 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.58
+ $Y=0.036 $X2=0.612 $Y2=0.036
r112 71 72 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.549
+ $Y=0.036 $X2=0.58 $Y2=0.036
r113 69 74 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.63 $Y2=0.036
r114 66 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.531 $Y2=0.036
r115 65 66 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.522 $Y2=0.036
r116 64 65 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.499
+ $Y=0.036 $X2=0.504 $Y2=0.036
r117 62 71 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.549 $Y2=0.036
r118 62 67 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.531 $Y2=0.036
r119 59 64 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.499 $Y2=0.036
r120 56 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r121 54 59 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r122 54 57 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.306 $Y2=0.036
r123 51 52 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.036 $X2=0.2115 $Y2=0.036
r124 49 56 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.288 $Y2=0.036
r125 49 52 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.2115 $Y2=0.036
r126 43 51 6.72222 $w=1.8e-08 $l=9.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.207 $Y2=0.036
r127 41 87 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.72 $Y=0.036 $X2=0.729 $Y2=0.045
r128 41 69 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.036 $X2=0.648 $Y2=0.036
r129 39 81 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.703 $Y=0.198
+ $X2=0.703 $Y2=0.198
r130 36 39 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.2025 $X2=0.7 $Y2=0.2025
r131 35 77 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.198
+ $X2=0.594 $Y2=0.198
r132 32 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2025 $X2=0.594 $Y2=0.2025
r133 31 35 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2025 $X2=0.594 $Y2=0.2025
r134 30 69 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036
+ $X2=0.648 $Y2=0.036
r135 27 30 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.054 $X2=0.648 $Y2=0.054
r136 26 30 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.054 $X2=0.648 $Y2=0.054
r137 25 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r138 22 25 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.054 $X2=0.54 $Y2=0.054
r139 21 25 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.054 $X2=0.54 $Y2=0.054
r140 20 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r141 17 20 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.054 $X2=0.432 $Y2=0.054
r142 16 20 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.054 $X2=0.432 $Y2=0.054
r143 15 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r144 12 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.054 $X2=0.324 $Y2=0.054
r145 11 15 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.054 $X2=0.324 $Y2=0.054
r146 10 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r147 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.054 $X2=0.216 $Y2=0.054
r148 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.054 $X2=0.216 $Y2=0.054
r149 5 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r150 2 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.054 $X2=0.108 $Y2=0.054
r151 1 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.054 $X2=0.108 $Y2=0.054
.ends


* END of "./NOR4xp75_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR4xp75_ASAP7_75t_R  VSS VDD D C B A Y
* 
* Y	Y
* A	A
* B	B
* C	C
* D	D
M0 N_Y_M0_d N_D_M0_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_D_M1_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_D_M2_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 VSS N_C_M3_g N_Y_M3_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 VSS N_C_M4_g N_Y_M4_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287 $Y=0.027
M5 VSS N_C_M5_g N_Y_M5_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_B_M6_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_B_M7_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_B_M8_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.503 $Y=0.027
M9 VSS N_A_M9_g N_Y_M9_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.557 $Y=0.027
M10 VSS N_A_M10_g N_Y_M10_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.611
+ $Y=0.027
M11 VSS N_A_M11_g N_Y_M11_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.665
+ $Y=0.027
M12 N_7_M12_d N_D_M12_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M13 N_7_M13_d N_D_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M14 N_7_M14_d N_D_M14_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M15 N_8_M15_d N_C_M15_g N_7_M15_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M16 N_8_M16_d N_C_M16_g N_7_M16_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M17 N_8_M17_d N_C_M17_g N_7_M17_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M18 N_9_M18_d N_B_M18_g N_8_M18_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M19 N_9_M19_d N_B_M19_g N_8_M19_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M20 N_9_M20_d N_B_M20_g N_8_M20_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M21 N_Y_M21_d N_A_M21_g N_9_M21_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M22 N_Y_M22_d N_A_M22_g N_9_M22_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M23 N_Y_M23_d N_A_M23_g N_9_M23_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
*
* 
* .include "NOR4xp75_ASAP7_75t_R.pex.sp.NOR4XP75_ASAP7_75T_R.pxi"
* BEGIN of "./NOR4xp75_ASAP7_75t_R.pex.sp.NOR4XP75_ASAP7_75T_R.pxi"
* File: NOR4xp75_ASAP7_75t_R.pex.sp.NOR4XP75_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:45:49 2017
* 
x_PM_NOR4XP75_ASAP7_75T_R%D N_D_M0_g N_D_M12_g N_D_M1_g N_D_M13_g N_D_M2_g
+ N_D_c_4_p N_D_M14_g D VSS PM_NOR4XP75_ASAP7_75T_R%D
x_PM_NOR4XP75_ASAP7_75T_R%C N_C_M3_g N_C_M15_g N_C_M4_g N_C_M16_g N_C_M5_g
+ N_C_c_20_n N_C_M17_g C VSS PM_NOR4XP75_ASAP7_75T_R%C
x_PM_NOR4XP75_ASAP7_75T_R%B N_B_M6_g N_B_M18_g N_B_M7_g N_B_M19_g N_B_M8_g
+ N_B_c_55_n N_B_M20_g B VSS PM_NOR4XP75_ASAP7_75T_R%B
x_PM_NOR4XP75_ASAP7_75T_R%A N_A_M9_g N_A_M21_g N_A_M10_g N_A_M22_g N_A_M11_g
+ N_A_c_89_n N_A_M23_g A VSS PM_NOR4XP75_ASAP7_75T_R%A
x_PM_NOR4XP75_ASAP7_75T_R%7 N_7_M13_d N_7_M12_d N_7_c_114_n N_7_M15_s N_7_M14_d
+ N_7_c_119_n N_7_M17_s N_7_M16_s N_7_c_121_n N_7_c_115_n N_7_c_117_n
+ N_7_c_123_n N_7_c_124_n N_7_c_125_n VSS PM_NOR4XP75_ASAP7_75T_R%7
x_PM_NOR4XP75_ASAP7_75T_R%8 N_8_M16_d N_8_M15_d N_8_c_142_n N_8_M18_s N_8_M17_d
+ N_8_c_158_n N_8_M20_s N_8_M19_s N_8_c_149_n N_8_c_144_n N_8_c_146_n
+ N_8_c_151_n N_8_c_147_n N_8_c_165_p VSS PM_NOR4XP75_ASAP7_75T_R%8
x_PM_NOR4XP75_ASAP7_75T_R%9 N_9_M19_d N_9_M18_d N_9_c_173_n N_9_M21_s N_9_M20_d
+ N_9_c_174_n N_9_M23_s N_9_M22_s N_9_c_181_n N_9_c_175_n N_9_c_177_n
+ N_9_c_179_n N_9_c_182_n N_9_c_183_n VSS PM_NOR4XP75_ASAP7_75T_R%9
x_PM_NOR4XP75_ASAP7_75T_R%Y N_Y_M1_d N_Y_M0_d N_Y_c_205_n N_Y_M3_s N_Y_M2_d
+ N_Y_c_247_n N_Y_M5_s N_Y_M4_s N_Y_c_210_n N_Y_M7_d N_Y_M6_d N_Y_c_220_n
+ N_Y_M9_s N_Y_M8_d N_Y_c_221_n N_Y_M11_s N_Y_M10_s N_Y_c_229_n N_Y_M22_d
+ N_Y_M21_d N_Y_c_232_n N_Y_M23_d N_Y_c_258_n N_Y_c_233_n N_Y_c_206_n
+ N_Y_c_208_n N_Y_c_212_n N_Y_c_213_n N_Y_c_216_n N_Y_c_218_n N_Y_c_225_n
+ N_Y_c_227_n N_Y_c_235_n N_Y_c_237_n N_Y_c_228_n N_Y_c_240_n N_Y_c_242_n
+ N_Y_c_243_n Y N_Y_c_245_n VSS PM_NOR4XP75_ASAP7_75T_R%Y
cc_1 N_D_M1_g N_C_M3_g 2.31381e-19 $X=0.135 $Y=0.054 $X2=0.243 $Y2=0.054
cc_2 N_D_M2_g N_C_M3_g 0.00344695f $X=0.189 $Y=0.054 $X2=0.243 $Y2=0.054
cc_3 N_D_M2_g N_C_M4_g 2.66145e-19 $X=0.189 $Y=0.054 $X2=0.297 $Y2=0.054
cc_4 N_D_c_4_p N_C_c_20_n 0.00139993f $X=0.189 $Y=0.135 $X2=0.351 $Y2=0.135
cc_5 D C 2.42911e-19 $X=0.081 $Y=0.138 $X2=0.3 $Y2=0.138
cc_6 N_D_c_4_p N_7_M13_d 3.47207e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.054
cc_7 N_D_c_4_p N_7_c_114_n 8.23937e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.135
cc_8 N_D_c_4_p N_7_c_115_n 0.00129866f $X=0.189 $Y=0.135 $X2=0.351 $Y2=0.054
cc_9 D N_7_c_115_n 7.8813e-19 $X=0.081 $Y=0.138 $X2=0.351 $Y2=0.054
cc_10 N_D_M1_g N_7_c_117_n 4.637e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_11 N_D_M2_g N_7_c_117_n 4.637e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_12 N_D_c_4_p N_Y_c_205_n 3.69297e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.135
cc_13 N_D_c_4_p N_Y_c_206_n 0.00126095f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_14 D N_Y_c_206_n 7.47007e-19 $X=0.081 $Y=0.138 $X2=0 $Y2=0
cc_15 N_D_M1_g N_Y_c_208_n 4.637e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_16 N_D_M2_g N_Y_c_208_n 4.637e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_17 N_C_M4_g N_B_M6_g 2.71887e-19 $X=0.297 $Y=0.054 $X2=0.081 $Y2=0.054
cc_18 N_C_M5_g N_B_M6_g 0.00333077f $X=0.351 $Y=0.054 $X2=0.081 $Y2=0.054
cc_19 N_C_M5_g N_B_M7_g 2.71887e-19 $X=0.351 $Y=0.054 $X2=0.135 $Y2=0.054
cc_20 N_C_c_20_n N_B_c_55_n 0.00136412f $X=0.351 $Y=0.135 $X2=0.189 $Y2=0.135
cc_21 C B 6.03898e-19 $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_22 C N_7_c_119_n 0.00300227f $X=0.3 $Y=0.138 $X2=0.135 $Y2=0.054
cc_23 N_C_c_20_n N_7_M17_s 3.53818e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_24 N_C_c_20_n N_7_c_121_n 8.23937e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_25 C N_7_c_121_n 2.5649e-19 $X=0.3 $Y=0.138 $X2=0.135 $Y2=0.2025
cc_26 C N_7_c_123_n 0.00101769f $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_27 N_C_M4_g N_7_c_124_n 2.38737e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_28 N_C_M3_g N_7_c_125_n 3.88389e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_29 C N_7_c_125_n 9.37582e-19 $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_30 N_C_c_20_n N_8_M16_d 3.46366e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.054
cc_31 N_C_c_20_n N_8_c_142_n 8.23937e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_32 C N_8_c_142_n 0.00158145f $X=0.3 $Y=0.138 $X2=0.081 $Y2=0.135
cc_33 N_C_M4_g N_8_c_144_n 2.60457e-19 $X=0.297 $Y=0.054 $X2=0.189 $Y2=0.2025
cc_34 C N_8_c_144_n 0.00445699f $X=0.3 $Y=0.138 $X2=0.189 $Y2=0.2025
cc_35 N_C_c_20_n N_8_c_146_n 8.71744e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_36 N_C_M5_g N_8_c_147_n 4.99916e-19 $X=0.351 $Y=0.054 $X2=0 $Y2=0
cc_37 N_C_c_20_n N_Y_c_210_n 3.69297e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_38 C N_Y_c_210_n 3.86867e-19 $X=0.3 $Y=0.138 $X2=0.135 $Y2=0.2025
cc_39 C N_Y_c_212_n 5.24578e-19 $X=0.3 $Y=0.138 $X2=0.135 $Y2=0.135
cc_40 N_C_M3_g N_Y_c_213_n 4.5519e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_41 N_C_c_20_n N_Y_c_213_n 6.79963e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_42 C N_Y_c_213_n 5.24578e-19 $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_43 N_C_M4_g N_Y_c_216_n 2.64924e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_44 C N_Y_c_216_n 0.00124933f $X=0.3 $Y=0.138 $X2=0 $Y2=0
cc_45 N_C_M5_g N_Y_c_218_n 4.67322e-19 $X=0.351 $Y=0.054 $X2=0 $Y2=0
cc_46 N_C_c_20_n N_Y_c_218_n 5.37353e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_47 N_B_M7_g N_A_M9_g 2.71887e-19 $X=0.459 $Y=0.054 $X2=0.081 $Y2=0.054
cc_48 N_B_M8_g N_A_M9_g 0.00357042f $X=0.513 $Y=0.054 $X2=0.081 $Y2=0.054
cc_49 N_B_M8_g N_A_M10_g 2.71887e-19 $X=0.513 $Y=0.054 $X2=0.135 $Y2=0.054
cc_50 N_B_c_55_n N_A_c_89_n 0.00121234f $X=0.513 $Y=0.135 $X2=0.189 $Y2=0.135
cc_51 B A 0.00192004f $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_52 N_B_c_55_n N_8_M20_s 3.67702e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_53 N_B_c_55_n N_8_c_149_n 8.69026e-19 $X=0.513 $Y=0.135 $X2=0.135 $Y2=0.2025
cc_54 B N_8_c_149_n 2.62694e-19 $X=0.521 $Y=0.138 $X2=0.135 $Y2=0.2025
cc_55 N_B_M7_g N_8_c_151_n 4.0114e-19 $X=0.459 $Y=0.054 $X2=0 $Y2=0
cc_56 B N_8_c_151_n 4.95077e-19 $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_57 N_B_M6_g N_8_c_147_n 4.15837e-19 $X=0.405 $Y=0.054 $X2=0 $Y2=0
cc_58 N_B_c_55_n N_8_c_147_n 0.00156237f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_59 N_B_c_55_n N_9_M19_d 3.67193e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.054
cc_60 N_B_c_55_n N_9_c_173_n 8.69026e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.135
cc_61 B N_9_c_174_n 0.00274961f $X=0.521 $Y=0.138 $X2=0.135 $Y2=0.054
cc_62 N_B_M6_g N_9_c_175_n 2.16933e-19 $X=0.405 $Y=0.054 $X2=0.189 $Y2=0.2025
cc_63 N_B_M7_g N_9_c_175_n 2.65027e-19 $X=0.459 $Y=0.054 $X2=0.189 $Y2=0.2025
cc_64 N_B_M8_g N_9_c_177_n 3.43821e-19 $X=0.513 $Y=0.054 $X2=0 $Y2=0
cc_65 B N_9_c_177_n 8.36482e-19 $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_66 B N_9_c_179_n 0.00101769f $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_67 N_B_c_55_n N_Y_c_220_n 3.75758e-19 $X=0.513 $Y=0.135 $X2=0.189 $Y2=0.135
cc_68 B N_Y_c_221_n 3.83412e-19 $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_69 N_B_M6_g N_Y_c_218_n 4.65034e-19 $X=0.405 $Y=0.054 $X2=0 $Y2=0
cc_70 N_B_M7_g N_Y_c_218_n 4.65034e-19 $X=0.459 $Y=0.054 $X2=0 $Y2=0
cc_71 N_B_c_55_n N_Y_c_218_n 0.00126591f $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_72 N_B_M8_g N_Y_c_225_n 2.57255e-19 $X=0.513 $Y=0.054 $X2=0 $Y2=0
cc_73 B N_Y_c_225_n 0.00123176f $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_74 B N_Y_c_227_n 4.04735e-19 $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_75 B N_Y_c_228_n 6.57587e-19 $X=0.521 $Y=0.138 $X2=0 $Y2=0
cc_76 N_A_c_89_n N_9_M23_s 3.67193e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_77 N_A_c_89_n N_9_c_181_n 8.69026e-19 $X=0.675 $Y=0.135 $X2=0.297 $Y2=0.2025
cc_78 N_A_M10_g N_9_c_182_n 2.38524e-19 $X=0.621 $Y=0.054 $X2=0 $Y2=0
cc_79 N_A_M9_g N_9_c_183_n 4.61191e-19 $X=0.567 $Y=0.054 $X2=0.297 $Y2=0.135
cc_80 N_A_c_89_n N_9_c_183_n 2.50471e-19 $X=0.675 $Y=0.135 $X2=0.297 $Y2=0.135
cc_81 N_A_c_89_n N_Y_c_229_n 3.75758e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_82 A N_Y_c_229_n 3.83412e-19 $X=0.621 $Y=0.138 $X2=0 $Y2=0
cc_83 N_A_c_89_n N_Y_M22_d 3.67575e-19 $X=0.675 $Y=0.135 $X2=0.297 $Y2=0.135
cc_84 N_A_c_89_n N_Y_c_232_n 8.69026e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_85 N_A_M11_g N_Y_c_233_n 4.38953e-19 $X=0.675 $Y=0.054 $X2=0 $Y2=0
cc_86 N_A_c_89_n N_Y_c_233_n 5.32086e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_87 N_A_M9_g N_Y_c_235_n 4.61191e-19 $X=0.567 $Y=0.054 $X2=0 $Y2=0
cc_88 N_A_c_89_n N_Y_c_235_n 7.74107e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_89 N_A_M10_g N_Y_c_237_n 2.64606e-19 $X=0.621 $Y=0.054 $X2=0 $Y2=0
cc_90 A N_Y_c_237_n 0.0012482f $X=0.621 $Y=0.138 $X2=0 $Y2=0
cc_91 N_A_c_89_n N_Y_c_228_n 4.94606e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_92 N_A_M10_g N_Y_c_240_n 2.77224e-19 $X=0.621 $Y=0.054 $X2=0 $Y2=0
cc_93 A N_Y_c_240_n 0.00123371f $X=0.621 $Y=0.138 $X2=0 $Y2=0
cc_94 N_A_c_89_n N_Y_c_242_n 8.61062e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_95 N_A_M11_g N_Y_c_243_n 4.5732e-19 $X=0.675 $Y=0.054 $X2=0 $Y2=0
cc_96 A Y 8.29246e-19 $X=0.621 $Y=0.138 $X2=0 $Y2=0
cc_97 A N_Y_c_245_n 8.29246e-19 $X=0.621 $Y=0.138 $X2=0 $Y2=0
cc_98 N_7_c_119_n N_8_c_142_n 0.00379429f $X=0.216 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_99 N_7_c_121_n N_8_c_142_n 0.00361461f $X=0.324 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_100 N_7_c_124_n N_8_c_142_n 0.00250918f $X=0.324 $Y=0.234 $X2=0.081 $Y2=0.135
cc_101 N_7_c_121_n N_8_c_158_n 0.0032677f $X=0.324 $Y=0.2025 $X2=0.135 $Y2=0.054
cc_102 N_7_c_124_n N_8_c_158_n 4.51105e-19 $X=0.324 $Y=0.234 $X2=0.135 $Y2=0.054
cc_103 N_7_c_119_n N_8_c_144_n 2.68768e-19 $X=0.216 $Y=0.2025 $X2=0.189
+ $Y2=0.2025
cc_104 N_7_c_124_n N_8_c_144_n 0.00723013f $X=0.324 $Y=0.234 $X2=0.189
+ $Y2=0.2025
cc_105 N_7_c_121_n N_8_c_146_n 0.00233206f $X=0.324 $Y=0.2025 $X2=0 $Y2=0
cc_106 N_7_c_124_n N_9_c_175_n 3.33393e-19 $X=0.324 $Y=0.234 $X2=0.189
+ $Y2=0.2025
cc_107 N_7_c_114_n N_Y_c_205_n 9.19308e-19 $X=0.108 $Y=0.2025 $X2=0.081
+ $Y2=0.135
cc_108 N_7_c_119_n N_Y_c_247_n 7.34324e-19 $X=0.216 $Y=0.2025 $X2=0.135
+ $Y2=0.054
cc_109 N_7_c_121_n N_Y_c_210_n 9.98826e-19 $X=0.324 $Y=0.2025 $X2=0.135
+ $Y2=0.2025
cc_110 N_7_c_115_n N_Y_c_206_n 2.27785e-19 $X=0.108 $Y=0.234 $X2=0 $Y2=0
cc_111 N_7_c_117_n N_Y_c_206_n 2.27785e-19 $X=0.207 $Y=0.234 $X2=0 $Y2=0
cc_112 N_8_c_158_n N_9_c_173_n 0.00317784f $X=0.378 $Y=0.2025 $X2=0.243
+ $Y2=0.135
cc_113 N_8_c_149_n N_9_c_173_n 0.00358852f $X=0.486 $Y=0.2025 $X2=0.243
+ $Y2=0.135
cc_114 N_8_c_165_p N_9_c_173_n 0.00233206f $X=0.4485 $Y=0.198 $X2=0.243
+ $Y2=0.135
cc_115 N_8_c_149_n N_9_c_174_n 0.00363127f $X=0.486 $Y=0.2025 $X2=0.297
+ $Y2=0.054
cc_116 N_8_c_151_n N_9_c_174_n 3.19711e-19 $X=0.485 $Y=0.198 $X2=0.297 $Y2=0.054
cc_117 N_8_c_158_n N_9_c_175_n 4.73069e-19 $X=0.378 $Y=0.2025 $X2=0.351
+ $Y2=0.2025
cc_118 N_8_c_149_n N_9_c_175_n 0.00250051f $X=0.486 $Y=0.2025 $X2=0.351
+ $Y2=0.2025
cc_119 N_8_c_165_p N_9_c_175_n 0.00744433f $X=0.4485 $Y=0.198 $X2=0.351
+ $Y2=0.2025
cc_120 N_8_c_146_n N_Y_c_218_n 0.00103693f $X=0.34 $Y=0.198 $X2=0 $Y2=0
cc_121 N_9_c_173_n N_Y_c_220_n 9.98826e-19 $X=0.432 $Y=0.2025 $X2=0.513
+ $Y2=0.135
cc_122 N_9_c_174_n N_Y_c_221_n 7.31912e-19 $X=0.54 $Y=0.2025 $X2=0 $Y2=0
cc_123 N_9_c_181_n N_Y_c_229_n 9.98826e-19 $X=0.648 $Y=0.2025 $X2=0.521
+ $Y2=0.138
cc_124 N_9_c_174_n N_Y_c_232_n 0.00362498f $X=0.54 $Y=0.2025 $X2=0.513 $Y2=0.135
cc_125 N_9_c_181_n N_Y_c_232_n 0.00348914f $X=0.648 $Y=0.2025 $X2=0.513
+ $Y2=0.135
cc_126 N_9_c_182_n N_Y_c_232_n 0.00250914f $X=0.648 $Y=0.234 $X2=0.513 $Y2=0.135
cc_127 N_9_c_181_n N_Y_c_258_n 0.00339247f $X=0.648 $Y=0.2025 $X2=0 $Y2=0
cc_128 N_9_c_182_n N_Y_c_258_n 2.9219e-19 $X=0.648 $Y=0.234 $X2=0 $Y2=0
cc_129 N_9_c_174_n N_Y_c_228_n 3.22784e-19 $X=0.54 $Y=0.2025 $X2=0 $Y2=0
cc_130 N_9_c_182_n N_Y_c_228_n 0.00739153f $X=0.648 $Y=0.234 $X2=0 $Y2=0
cc_131 N_9_c_181_n N_Y_c_242_n 0.00233206f $X=0.648 $Y=0.2025 $X2=0 $Y2=0

* END of "./NOR4xp75_ASAP7_75t_R.pex.sp.NOR4XP75_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: NOR5xp2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:46:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "NOR5xp2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./NOR5xp2_ASAP7_75t_R.pex.sp.pex"
* File: NOR5xp2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:46:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_NOR5XP2_ASAP7_75T_R%A 2 5 7 10 VSS
c11 10 VSS 0.00172965f $X=0.081 $Y=0.135
c12 5 VSS 0.00329644f $X=0.081 $Y=0.136
c13 2 VSS 0.0641893f $X=0.081 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.136 $X2=0.081
+ $Y2=0.136
r15 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.136 $X2=0.081 $Y2=0.2025
r16 2 5 307.213 $w=2e-08 $l=8.2e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.136
.ends

.subckt PM_NOR5XP2_ASAP7_75T_R%B 2 5 7 10 VSS
c13 10 VSS 0.00238574f $X=0.135 $Y=0.136
c14 5 VSS 0.0017057f $X=0.135 $Y=0.1355
c15 2 VSS 0.060473f $X=0.135 $Y=0.054
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.136 $X2=0.135
+ $Y2=0.136
r17 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.2025
r18 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.1355
.ends

.subckt PM_NOR5XP2_ASAP7_75T_R%C 2 5 7 10 VSS
c11 10 VSS 0.00220204f $X=0.189 $Y=0.135
c12 5 VSS 0.00160244f $X=0.189 $Y=0.1355
c13 2 VSS 0.0597904f $X=0.189 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.136 $X2=0.189
+ $Y2=0.136
r15 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1355 $X2=0.189 $Y2=0.2025
r16 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.1355
.ends

.subckt PM_NOR5XP2_ASAP7_75T_R%D 2 5 7 10 VSS
c10 10 VSS 0.00239098f $X=0.243 $Y=0.135
c11 5 VSS 0.0016285f $X=0.243 $Y=0.1355
c12 2 VSS 0.0597088f $X=0.243 $Y=0.054
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.136 $X2=0.243
+ $Y2=0.136
r14 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1355 $X2=0.243 $Y2=0.2025
r15 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.1355
.ends

.subckt PM_NOR5XP2_ASAP7_75T_R%E 2 5 7 10 VSS
c7 10 VSS 0.00562468f $X=0.297 $Y=0.135
c8 5 VSS 0.00255331f $X=0.297 $Y=0.1355
c9 2 VSS 0.0636337f $X=0.297 $Y=0.054
r10 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.136 $X2=0.297
+ $Y2=0.136
r11 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.1355 $X2=0.297 $Y2=0.2025
r12 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.1355
.ends

.subckt PM_NOR5XP2_ASAP7_75T_R%Y 1 2 5 6 7 10 11 14 16 19 24 26 28 33 35 41 43
+ 48 50 55 VSS
c22 58 VSS 8.89192e-19 $X=0.0455 $Y=0.234
c23 57 VSS 0.00360091f $X=0.037 $Y=0.234
c24 55 VSS 0.00319348f $X=0.054 $Y=0.234
c25 50 VSS 0.00146362f $X=0.306 $Y=0.036
c26 49 VSS 0.00631462f $X=0.288 $Y=0.036
c27 48 VSS 0.00146362f $X=0.252 $Y=0.036
c28 47 VSS 0.00377381f $X=0.234 $Y=0.036
c29 45 VSS 0.00496339f $X=0.324 $Y=0.036
c30 43 VSS 0.00146362f $X=0.198 $Y=0.036
c31 42 VSS 0.00631462f $X=0.18 $Y=0.036
c32 41 VSS 0.00146362f $X=0.144 $Y=0.036
c33 40 VSS 0.00284382f $X=0.126 $Y=0.036
c34 36 VSS 9.63895e-19 $X=0.099 $Y=0.036
c35 35 VSS 0.00142296f $X=0.09 $Y=0.036
c36 34 VSS 1.68773e-19 $X=0.072 $Y=0.036
c37 33 VSS 0.00513619f $X=0.07 $Y=0.036
c38 29 VSS 0.00369107f $X=0.037 $Y=0.036
c39 28 VSS 5.93854e-19 $X=0.027 $Y=0.2115
c40 26 VSS 0.00205605f $X=0.027 $Y=0.1055
c41 25 VSS 0.00170849f $X=0.027 $Y=0.07
c42 24 VSS 0.00468624f $X=0.025 $Y=0.141
c43 22 VSS 5.71859e-19 $X=0.027 $Y=0.225
c44 19 VSS 0.0033504f $X=0.056 $Y=0.2025
c45 16 VSS 4.49354e-19 $X=0.071 $Y=0.2025
c46 14 VSS 0.00613723f $X=0.322 $Y=0.054
c47 10 VSS 0.0079214f $X=0.216 $Y=0.054
c48 6 VSS 5.3314e-19 $X=0.233 $Y=0.054
c49 5 VSS 0.00790645f $X=0.108 $Y=0.054
c50 1 VSS 5.3314e-19 $X=0.125 $Y=0.054
r51 57 58 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.037
+ $Y=0.234 $X2=0.0455 $Y2=0.234
r52 55 58 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0455 $Y2=0.234
r53 52 57 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.037 $Y2=0.234
r54 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r55 48 49 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r56 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r57 45 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.306 $Y2=0.036
r58 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r59 41 42 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.18 $Y2=0.036
r60 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r61 38 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.234 $Y2=0.036
r62 38 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.198 $Y2=0.036
r63 35 36 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.099 $Y2=0.036
r64 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r65 33 34 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.07
+ $Y=0.036 $X2=0.072 $Y2=0.036
r66 31 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r67 31 36 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.099 $Y2=0.036
r68 29 33 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.037
+ $Y=0.036 $X2=0.07 $Y2=0.036
r69 27 28 0.804167 $w=2e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.198 $X2=0.027 $Y2=0.2115
r70 25 26 2.11466 $w=2e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.1055
r71 24 27 3.39537 $w=2e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.141 $X2=0.027 $Y2=0.198
r72 24 26 2.11466 $w=2e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.141 $X2=0.027 $Y2=0.1055
r73 22 52 0.00634181 $w=2e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.234
r74 22 28 0.804167 $w=2e-08 $l=1.35e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.2115
r75 21 29 0.685354 $w=2e-08 $l=1.3784e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.037 $Y2=0.036
r76 21 25 1.4892 $w=2e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r77 19 55 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r78 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r79 14 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r80 11 14 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.054 $X2=0.322 $Y2=0.054
r81 10 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r82 7 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.054 $X2=0.216 $Y2=0.054
r83 6 10 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.054 $X2=0.216 $Y2=0.054
r84 5 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r85 2 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.054 $X2=0.108 $Y2=0.054
r86 1 5 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.054 $X2=0.108 $Y2=0.054
.ends

.subckt PM_NOR5XP2_ASAP7_75T_R%9 1 2 VSS
c0 1 VSS 0.00228332f $X=0.125 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends

.subckt PM_NOR5XP2_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00228332f $X=0.179 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends

.subckt PM_NOR5XP2_ASAP7_75T_R%11 1 2 VSS
c0 1 VSS 0.00228332f $X=0.233 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.199 $Y2=0.2025
.ends

.subckt PM_NOR5XP2_ASAP7_75T_R%12 1 2 VSS
c0 1 VSS 0.00228332f $X=0.287 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.253 $Y2=0.2025
.ends


* END of "./NOR5xp2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt NOR5xp2_ASAP7_75t_R  VSS VDD A B C D E Y
* 
* Y	Y
* E	E
* D	D
* C	C
* B	B
* A	A
M0 N_Y_M0_d N_A_M0_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 VSS N_B_M1_g N_Y_M1_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_C_M2_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 VSS N_D_M3_g N_Y_M3_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_E_M4_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287 $Y=0.027
M5 N_9_M5_d N_A_M5_g N_Y_M5_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M6 N_10_M6_d N_B_M6_g N_9_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 N_11_M7_d N_C_M7_g N_10_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M8 N_12_M8_d N_D_M8_g N_11_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M9 VDD N_E_M9_g N_12_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
*
* 
* .include "NOR5xp2_ASAP7_75t_R.pex.sp.NOR5XP2_ASAP7_75T_R.pxi"
* BEGIN of "./NOR5xp2_ASAP7_75t_R.pex.sp.NOR5XP2_ASAP7_75T_R.pxi"
* File: NOR5xp2_ASAP7_75t_R.pex.sp.NOR5XP2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:46:11 2017
* 
x_PM_NOR5XP2_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M5_g A VSS
+ PM_NOR5XP2_ASAP7_75T_R%A
x_PM_NOR5XP2_ASAP7_75T_R%B N_B_M1_g N_B_c_13_n N_B_M6_g B VSS
+ PM_NOR5XP2_ASAP7_75T_R%B
x_PM_NOR5XP2_ASAP7_75T_R%C N_C_M2_g N_C_c_27_n N_C_M7_g C VSS
+ PM_NOR5XP2_ASAP7_75T_R%C
x_PM_NOR5XP2_ASAP7_75T_R%D N_D_M3_g N_D_c_38_n N_D_M8_g D VSS
+ PM_NOR5XP2_ASAP7_75T_R%D
x_PM_NOR5XP2_ASAP7_75T_R%E N_E_M4_g N_E_c_48_n N_E_M9_g E VSS
+ PM_NOR5XP2_ASAP7_75T_R%E
x_PM_NOR5XP2_ASAP7_75T_R%Y N_Y_M1_s N_Y_M0_d N_Y_c_53_n N_Y_M3_s N_Y_M2_d
+ N_Y_c_66_n N_Y_M4_d N_Y_c_72_n N_Y_M5_s N_Y_c_54_n Y N_Y_c_56_n N_Y_c_62_n
+ N_Y_c_57_n N_Y_c_58_n N_Y_c_63_n N_Y_c_67_n N_Y_c_70_n N_Y_c_73_n N_Y_c_65_n
+ VSS PM_NOR5XP2_ASAP7_75T_R%Y
x_PM_NOR5XP2_ASAP7_75T_R%9 N_9_M6_s N_9_M5_d VSS PM_NOR5XP2_ASAP7_75T_R%9
x_PM_NOR5XP2_ASAP7_75T_R%10 N_10_M7_s N_10_M6_d VSS PM_NOR5XP2_ASAP7_75T_R%10
x_PM_NOR5XP2_ASAP7_75T_R%11 N_11_M8_s N_11_M7_d VSS PM_NOR5XP2_ASAP7_75T_R%11
x_PM_NOR5XP2_ASAP7_75T_R%12 N_12_M9_s N_12_M8_d VSS PM_NOR5XP2_ASAP7_75T_R%12
cc_1 N_A_M0_g N_B_M1_g 0.00357042f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A_c_2_p N_B_c_13_n 7.98811e-19 $X=0.081 $Y=0.136 $X2=0.135 $Y2=0.1355
cc_3 A B 0.00611879f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.136
cc_4 N_A_M0_g N_C_M2_g 2.71887e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 A N_Y_c_53_n 3.31541e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.1355
cc_6 N_A_c_2_p N_Y_c_54_n 3.06446e-19 $X=0.081 $Y=0.136 $X2=0 $Y2=0
cc_7 A N_Y_c_54_n 0.00125785f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_8 A N_Y_c_56_n 0.00557682f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_A_c_2_p N_Y_c_57_n 2.36937e-19 $X=0.081 $Y=0.136 $X2=0 $Y2=0
cc_10 N_A_M0_g N_Y_c_58_n 2.57864e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_11 A N_Y_c_58_n 0.00123625f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_12 N_B_M1_g N_C_M2_g 0.00333077f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_13 N_B_c_13_n N_C_c_27_n 7.92653e-19 $X=0.135 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_14 B C 0.00817592f $X=0.135 $Y=0.136 $X2=0.081 $Y2=0.135
cc_15 N_B_M1_g N_D_M3_g 2.71887e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_16 B N_Y_c_53_n 3.31541e-19 $X=0.135 $Y=0.136 $X2=0.081 $Y2=0.136
cc_17 B N_Y_c_54_n 5.05783e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_18 B N_Y_c_62_n 2.96571e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_19 N_B_M1_g N_Y_c_63_n 2.64924e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_20 B N_Y_c_63_n 0.00125705f $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_21 B N_Y_c_65_n 4.62679e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_22 N_C_M2_g N_D_M3_g 0.0035196f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_23 N_C_c_27_n N_D_c_38_n 7.90494e-19 $X=0.189 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_24 C D 0.00819209f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_25 N_C_M2_g N_E_M4_g 2.66145e-19 $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_26 C N_Y_c_66_n 3.31541e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_27 N_C_M2_g N_Y_c_67_n 2.64924e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_28 C N_Y_c_67_n 0.00125705f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_29 N_D_M3_g N_E_M4_g 0.0032073f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_30 N_D_c_38_n N_E_c_48_n 8.31912e-19 $X=0.243 $Y=0.1355 $X2=0.135 $Y2=0.1355
cc_31 D E 0.00809651f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.136
cc_32 D N_Y_c_66_n 3.31541e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.136
cc_33 N_D_M3_g N_Y_c_70_n 2.64924e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_34 D N_Y_c_70_n 0.00125705f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_35 E N_Y_c_72_n 2.02161e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_36 N_E_M4_g N_Y_c_73_n 2.64924e-19 $X=0.297 $Y=0.054 $X2=0 $Y2=0
cc_37 E N_Y_c_73_n 0.00125705f $X=0.297 $Y=0.135 $X2=0 $Y2=0

* END of "./NOR5xp2_ASAP7_75t_R.pex.sp.NOR5XP2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: AND2x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 11:58:42 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AND2x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./AND2x2_ASAP7_75t_R.pex.sp.pex"
* File: AND2x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 11:58:42 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AND2X2_ASAP7_75T_R%B 2 5 7 23 VSS
c7 23 VSS 0.0158133f $X=0.073 $Y=0.133
c8 5 VSS 0.00454789f $X=0.081 $Y=0.1345
c9 2 VSS 0.0646732f $X=0.081 $Y=0.0675
r10 20 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.07 $Y=0.135 $X2=0.07
+ $Y2=0.135
r11 5 20 9.56522 $w=2.3e-08 $l=1.1e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1345 $X2=0.07 $Y2=0.1345
r12 5 7 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1345 $X2=0.081 $Y2=0.216
r13 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.1345
.ends

.subckt PM_AND2X2_ASAP7_75T_R%A 2 5 7 10 VSS
c17 10 VSS 0.00120225f $X=0.135 $Y=0.133
c18 5 VSS 0.00154473f $X=0.135 $Y=0.135
c19 2 VSS 0.0586444f $X=0.135 $Y=0.0675
r20 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r21 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r22 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AND2X2_ASAP7_75T_R%5 2 7 10 13 15 17 20 22 23 26 29 32 34 35 38 39 46
+ 48 49 50 52 53 54 58 60 VSS
c37 61 VSS 1.13166e-19 $X=0.1845 $Y=0.135
c38 60 VSS 1.73204e-19 $X=0.18 $Y=0.135
c39 58 VSS 5.7598e-19 $X=0.189 $Y=0.135
c40 54 VSS 3.97206e-19 $X=0.171 $Y=0.2
c41 53 VSS 0.00124019f $X=0.171 $Y=0.184
c42 52 VSS 6.48298e-19 $X=0.171 $Y=0.225
c43 50 VSS 3.97206e-19 $X=0.171 $Y=0.086
c44 49 VSS 6.19813e-19 $X=0.171 $Y=0.07
c45 48 VSS 0.00115863f $X=0.171 $Y=0.126
c46 46 VSS 0.00146362f $X=0.144 $Y=0.234
c47 45 VSS 0.00437783f $X=0.126 $Y=0.234
c48 40 VSS 0.00574629f $X=0.162 $Y=0.234
c49 39 VSS 0.00146362f $X=0.144 $Y=0.036
c50 38 VSS 0.00291865f $X=0.126 $Y=0.036
c51 37 VSS 0.00102009f $X=0.094 $Y=0.036
c52 36 VSS 0.00204372f $X=0.084 $Y=0.036
c53 35 VSS 0.00211324f $X=0.063 $Y=0.036
c54 34 VSS 0.00554029f $X=0.162 $Y=0.036
c55 31 VSS 2.30525e-19 $X=0.054 $Y=0.07
c56 29 VSS 1.03918e-19 $X=0.054 $Y=0.072
c57 26 VSS 0.00759416f $X=0.108 $Y=0.216
c58 22 VSS 5.65078e-19 $X=0.125 $Y=0.216
c59 20 VSS 0.00466594f $X=0.056 $Y=0.0675
c60 17 VSS 4.64427e-19 $X=0.071 $Y=0.0675
c61 13 VSS 0.00493701f $X=0.243 $Y=0.1345
c62 10 VSS 0.0639835f $X=0.243 $Y=0.0675
c63 2 VSS 0.0613324f $X=0.189 $Y=0.0675
r64 60 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.1845 $Y2=0.135
r65 58 61 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.135 $X2=0.1845 $Y2=0.135
r66 55 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.135 $X2=0.18 $Y2=0.135
r67 53 54 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.184 $X2=0.171 $Y2=0.2
r68 52 54 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.225 $X2=0.171 $Y2=0.2
r69 51 55 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.144 $X2=0.171 $Y2=0.135
r70 51 53 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.144 $X2=0.171 $Y2=0.184
r71 49 50 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.07 $X2=0.171 $Y2=0.086
r72 48 55 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.126 $X2=0.171 $Y2=0.135
r73 48 50 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.126 $X2=0.171 $Y2=0.086
r74 47 49 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.045 $X2=0.171 $Y2=0.07
r75 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r76 42 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r77 40 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.234 $X2=0.171 $Y2=0.225
r78 40 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.144 $Y2=0.234
r79 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r80 37 38 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.036 $X2=0.126 $Y2=0.036
r81 36 37 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.084
+ $Y=0.036 $X2=0.094 $Y2=0.036
r82 35 36 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.036 $X2=0.084 $Y2=0.036
r83 34 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.036 $X2=0.171 $Y2=0.045
r84 34 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.144 $Y2=0.036
r85 31 32 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.07 $X2=0.054 $Y2=0.071
r86 29 32 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.072 $X2=0.054 $Y2=0.071
r87 27 35 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.054 $Y=0.045 $X2=0.063 $Y2=0.036
r88 27 31 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.045 $X2=0.054 $Y2=0.07
r89 26 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r90 23 26 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.216 $X2=0.108 $Y2=0.216
r91 22 26 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.216 $X2=0.108 $Y2=0.216
r92 20 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.072 $X2=0.054
+ $Y2=0.072
r93 17 20 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r94 13 15 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1345 $X2=0.243 $Y2=0.2025
r95 10 13 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.1345
r96 5 13 46.9565 $w=2.3e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.1345 $X2=0.243 $Y2=0.1345
r97 5 58 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r98 5 7 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1345 $X2=0.189 $Y2=0.2025
r99 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.1345
.ends

.subckt PM_AND2X2_ASAP7_75T_R%Y 1 2 5 6 7 10 13 18 21 22 23 24 28 30 31 32 VSS
c18 34 VSS 0.00101302f $X=0.297 $Y=0.2045
c19 32 VSS 7.93583e-20 $X=0.297 $Y=0.14575
c20 31 VSS 7.74562e-19 $X=0.297 $Y=0.144
c21 30 VSS 0.00227931f $X=0.297 $Y=0.126
c22 29 VSS 0.00176873f $X=0.297 $Y=0.086
c23 28 VSS 0.00218466f $X=0.297 $Y=0.1475
c24 26 VSS 7.5805e-19 $X=0.297 $Y=0.225
c25 24 VSS 0.00212518f $X=0.225 $Y=0.234
c26 23 VSS 0.0112478f $X=0.288 $Y=0.234
c27 22 VSS 0.00212518f $X=0.225 $Y=0.036
c28 21 VSS 0.0112488f $X=0.288 $Y=0.036
c29 18 VSS 8.76752e-19 $X=0.216 $Y=0.198
c30 13 VSS 8.76752e-19 $X=0.216 $Y=0.072
c31 10 VSS 0.011152f $X=0.216 $Y=0.2025
c32 6 VSS 5.945e-19 $X=0.233 $Y=0.2025
c33 5 VSS 0.0108676f $X=0.216 $Y=0.0675
c34 1 VSS 5.945e-19 $X=0.233 $Y=0.0675
r35 33 34 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.184 $X2=0.297 $Y2=0.2045
r36 31 32 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.144 $X2=0.297 $Y2=0.14575
r37 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.144
r38 29 30 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.086 $X2=0.297 $Y2=0.126
r39 28 33 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1475 $X2=0.297 $Y2=0.184
r40 28 32 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1475 $X2=0.297 $Y2=0.14575
r41 26 34 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.2045
r42 25 29 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.086
r43 23 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.234 $X2=0.297 $Y2=0.225
r44 23 24 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.225 $Y2=0.234
r45 21 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r46 21 22 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.225 $Y2=0.036
r47 16 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.225 $X2=0.225 $Y2=0.234
r48 16 18 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.225 $X2=0.216 $Y2=0.198
r49 11 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.045 $X2=0.225 $Y2=0.036
r50 11 13 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.045 $X2=0.216 $Y2=0.072
r51 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r52 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r53 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r54 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072 $X2=0.216
+ $Y2=0.072
r55 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r56 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends

.subckt PM_AND2X2_ASAP7_75T_R%7 1 2 VSS
c1 1 VSS 0.0018307f $X=0.125 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends


* END of "./AND2x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt AND2x2_ASAP7_75t_R  VSS VDD B A Y
* 
* Y	Y
* A	A
* B	B
M0 N_7_M0_d N_B_M0_g N_5_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_A_M1_g N_7_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_5_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_5_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_5_M4_d N_B_M4_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M5 VDD N_A_M5_g N_5_M5_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
M6 N_Y_M6_d N_5_M6_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M7 N_Y_M7_d N_5_M7_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
*
* 
* .include "AND2x2_ASAP7_75t_R.pex.sp.AND2X2_ASAP7_75T_R.pxi"
* BEGIN of "./AND2x2_ASAP7_75t_R.pex.sp.AND2X2_ASAP7_75T_R.pxi"
* File: AND2x2_ASAP7_75t_R.pex.sp.AND2X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 11:58:42 2017
* 
x_PM_AND2X2_ASAP7_75T_R%B N_B_M0_g N_B_c_2_p N_B_M4_g B VSS
+ PM_AND2X2_ASAP7_75T_R%B
x_PM_AND2X2_ASAP7_75T_R%A N_A_M1_g N_A_c_9_n N_A_M5_g A VSS
+ PM_AND2X2_ASAP7_75T_R%A
x_PM_AND2X2_ASAP7_75T_R%5 N_5_M2_g N_5_M6_g N_5_M3_g N_5_c_31_n N_5_M7_g
+ N_5_M0_s N_5_c_26_n N_5_M5_s N_5_M4_d N_5_c_33_n N_5_c_27_n N_5_c_34_n
+ N_5_c_45_p N_5_c_28_n N_5_c_61_p N_5_c_35_n N_5_c_37_n N_5_c_39_n N_5_c_50_p
+ N_5_c_40_n N_5_c_56_p N_5_c_41_n N_5_c_52_p N_5_c_59_p N_5_c_42_n VSS
+ PM_AND2X2_ASAP7_75T_R%5
x_PM_AND2X2_ASAP7_75T_R%Y N_Y_M3_d N_Y_M2_d N_Y_c_63_n N_Y_M7_d N_Y_M6_d
+ N_Y_c_66_n N_Y_c_68_n N_Y_c_70_n N_Y_c_72_n N_Y_c_73_n N_Y_c_74_n N_Y_c_75_n Y
+ N_Y_c_76_n N_Y_c_78_n N_Y_c_79_n VSS PM_AND2X2_ASAP7_75T_R%Y
x_PM_AND2X2_ASAP7_75T_R%7 N_7_M1_s N_7_M0_d VSS PM_AND2X2_ASAP7_75T_R%7
cc_1 N_B_M0_g N_A_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_B_c_2_p N_A_c_9_n 0.00127799f $X=0.081 $Y=0.1345 $X2=0.135 $Y2=0.135
cc_3 B A 0.00188262f $X=0.073 $Y=0.133 $X2=0.135 $Y2=0.133
cc_4 N_B_M0_g N_5_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 B N_5_c_26_n 8.18408e-19 $X=0.073 $Y=0.133 $X2=0 $Y2=0
cc_6 B N_5_c_27_n 6.29493e-19 $X=0.073 $Y=0.133 $X2=0 $Y2=0
cc_7 B N_5_c_28_n 0.00447544f $X=0.073 $Y=0.133 $X2=0 $Y2=0
cc_8 N_A_M1_g N_5_M2_g 0.00284417f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_9 N_A_M1_g N_5_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_10 N_A_c_9_n N_5_c_31_n 0.00151388f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_11 A N_5_c_26_n 4.99565e-19 $X=0.135 $Y=0.133 $X2=0.07 $Y2=0.135
cc_12 A N_5_c_33_n 3.84694e-19 $X=0.135 $Y=0.133 $X2=0.07 $Y2=0.1345
cc_13 A N_5_c_34_n 4.32839e-19 $X=0.135 $Y=0.133 $X2=0 $Y2=0
cc_14 N_A_M1_g N_5_c_35_n 2.64276e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_15 A N_5_c_35_n 0.00125352f $X=0.135 $Y=0.133 $X2=0 $Y2=0
cc_16 N_A_M1_g N_5_c_37_n 2.64276e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_17 A N_5_c_37_n 0.00125352f $X=0.135 $Y=0.133 $X2=0 $Y2=0
cc_18 A N_5_c_39_n 0.00268918f $X=0.135 $Y=0.133 $X2=0 $Y2=0
cc_19 A N_5_c_40_n 0.00268918f $X=0.135 $Y=0.133 $X2=0 $Y2=0
cc_20 A N_5_c_41_n 0.00268918f $X=0.135 $Y=0.133 $X2=0 $Y2=0
cc_21 A N_5_c_42_n 0.00268918f $X=0.135 $Y=0.133 $X2=0 $Y2=0
cc_22 N_5_c_31_n N_Y_M3_d 3.89916e-19 $X=0.243 $Y=0.1345 $X2=0.081 $Y2=0.0675
cc_23 N_5_c_31_n N_Y_c_63_n 8.45347e-19 $X=0.243 $Y=0.1345 $X2=0.081 $Y2=0.1345
cc_24 N_5_c_45_p N_Y_c_63_n 0.00135217f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.1345
cc_25 N_5_c_31_n N_Y_M7_d 3.83395e-19 $X=0.243 $Y=0.1345 $X2=0.081 $Y2=0.216
cc_26 N_5_c_31_n N_Y_c_66_n 8.01479e-19 $X=0.243 $Y=0.1345 $X2=0 $Y2=0
cc_27 N_5_c_41_n N_Y_c_66_n 0.00135358f $X=0.171 $Y=0.184 $X2=0 $Y2=0
cc_28 N_5_c_31_n N_Y_c_68_n 2.51608e-19 $X=0.243 $Y=0.1345 $X2=0 $Y2=0
cc_29 N_5_c_50_p N_Y_c_68_n 0.0017671f $X=0.171 $Y=0.07 $X2=0 $Y2=0
cc_30 N_5_c_31_n N_Y_c_70_n 2.48871e-19 $X=0.243 $Y=0.1345 $X2=0 $Y2=0
cc_31 N_5_c_52_p N_Y_c_70_n 0.0017583f $X=0.171 $Y=0.2 $X2=0 $Y2=0
cc_32 N_5_M3_g N_Y_c_72_n 2.88603e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_33 N_5_c_45_p N_Y_c_73_n 0.0017671f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_34 N_5_M3_g N_Y_c_74_n 2.89885e-19 $X=0.243 $Y=0.0675 $X2=0.073 $Y2=0.133
cc_35 N_5_c_56_p N_Y_c_75_n 0.0017583f $X=0.171 $Y=0.225 $X2=0 $Y2=0
cc_36 N_5_c_31_n N_Y_c_76_n 5.21087e-19 $X=0.243 $Y=0.1345 $X2=0 $Y2=0
cc_37 N_5_c_39_n N_Y_c_76_n 3.97371e-19 $X=0.171 $Y=0.126 $X2=0 $Y2=0
cc_38 N_5_c_59_p N_Y_c_78_n 2.27943e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_39 N_5_c_41_n N_Y_c_79_n 4.03366e-19 $X=0.171 $Y=0.184 $X2=0 $Y2=0
cc_40 N_5_c_61_p N_7_M1_s 4.53269e-19 $X=0.126 $Y=0.036 $X2=0.081 $Y2=0.0675

* END of "./AND2x2_ASAP7_75t_R.pex.sp.AND2X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: AND2x4_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 11:59:04 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AND2x4_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./AND2x4_ASAP7_75t_R.pex.sp.pex"
* File: AND2x4_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 11:59:04 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AND2X4_ASAP7_75T_R%A 2 5 7 10 13 15 21 22 23 24 25 27 31 35 37 38 VSS
c27 38 VSS 0.00255655f $X=0.243 $Y=0.121
c28 37 VSS 8.45284e-19 $X=0.243 $Y=0.064
c29 35 VSS 2.3666e-19 $X=0.243 $Y=0.135
c30 32 VSS 0.00189145f $X=0.216 $Y=0.037
c31 31 VSS 0.00636831f $X=0.198 $Y=0.037
c32 30 VSS 0.00199175f $X=0.115 $Y=0.037
c33 29 VSS 3.03073e-19 $X=0.094 $Y=0.037
c34 28 VSS 0.0030786f $X=0.09 $Y=0.037
c35 27 VSS 0.00438018f $X=0.234 $Y=0.037
c36 25 VSS 0.00242134f $X=0.083 $Y=0.14
c37 24 VSS 3.59668e-19 $X=0.081 $Y=0.121
c38 23 VSS 0.0011834f $X=0.081 $Y=0.107
c39 22 VSS 9.44831e-19 $X=0.081 $Y=0.082
c40 21 VSS 8.45284e-19 $X=0.081 $Y=0.064
c41 13 VSS 9.42534e-19 $X=0.243 $Y=0.135
c42 10 VSS 0.059423f $X=0.243 $Y=0.0675
c43 5 VSS 0.00198216f $X=0.081 $Y=0.135
c44 2 VSS 0.0627695f $X=0.081 $Y=0.0675
r45 37 38 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.064 $X2=0.243 $Y2=0.121
r46 35 38 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.121
r47 33 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.046 $X2=0.243 $Y2=0.064
r48 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.037 $X2=0.216 $Y2=0.037
r49 30 31 5.6358 $w=1.8e-08 $l=8.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.115
+ $Y=0.037 $X2=0.198 $Y2=0.037
r50 29 30 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.037 $X2=0.115 $Y2=0.037
r51 28 29 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.037 $X2=0.094 $Y2=0.037
r52 27 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.037 $X2=0.243 $Y2=0.046
r53 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.037 $X2=0.216 $Y2=0.037
r54 24 25 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.121 $X2=0.081 $Y2=0.135
r55 23 24 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.107 $X2=0.081 $Y2=0.121
r56 22 23 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.082 $X2=0.081 $Y2=0.107
r57 21 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.064 $X2=0.081 $Y2=0.082
r58 17 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.046 $X2=0.09 $Y2=0.037
r59 17 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.046 $X2=0.081 $Y2=0.064
r60 13 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r61 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r62 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r63 5 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r64 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r65 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AND2X4_ASAP7_75T_R%B 2 7 10 13 15 18 22 VSS
c23 22 VSS 4.12915e-19 $X=0.135 $Y=0.152
c24 18 VSS 4.05597e-19 $X=0.135 $Y=0.135
c25 13 VSS 0.00443352f $X=0.189 $Y=0.135
c26 10 VSS 0.0626014f $X=0.189 $Y=0.0675
c27 2 VSS 0.0615487f $X=0.135 $Y=0.0675
r28 18 22 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.152
r29 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r30 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r31 5 13 60 $w=1.8e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135 $Y=0.135
+ $X2=0.189 $Y2=0.135
r32 5 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r33 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r34 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AND2X4_ASAP7_75T_R%5 2 7 10 15 18 23 26 29 31 33 34 37 38 39 42 43 44
+ 55 56 57 63 64 71 75 79 80 83 VSS
c49 86 VSS 6.58501e-19 $X=0.207 $Y=0.234
c50 85 VSS 0.00176786f $X=0.198 $Y=0.234
c51 83 VSS 0.00285708f $X=0.216 $Y=0.234
c52 80 VSS 4.93096e-19 $X=0.1885 $Y=0.191
c53 79 VSS 3.73908e-19 $X=0.297 $Y=0.166
c54 75 VSS 6.51961e-19 $X=0.297 $Y=0.135
c55 73 VSS 7.72048e-19 $X=0.297 $Y=0.182
c56 72 VSS 0.00254231f $X=0.27 $Y=0.191
c57 71 VSS 4.66176e-19 $X=0.252 $Y=0.191
c58 70 VSS 1.69914e-19 $X=0.234 $Y=0.191
c59 69 VSS 6.30164e-19 $X=0.231 $Y=0.191
c60 67 VSS 0.00194692f $X=0.288 $Y=0.191
c61 66 VSS 0.00121124f $X=0.189 $Y=0.225
c62 64 VSS 2.55645e-19 $X=0.189 $Y=0.15
c63 63 VSS 6.49295e-20 $X=0.189 $Y=0.107
c64 62 VSS 5.03482e-19 $X=0.189 $Y=0.182
c65 57 VSS 9.05837e-19 $X=0.18 $Y=0.073
c66 56 VSS 0.0053518f $X=0.179 $Y=0.234
c67 55 VSS 0.00142296f $X=0.144 $Y=0.234
c68 54 VSS 0.00105114f $X=0.126 $Y=0.234
c69 53 VSS 0.00346796f $X=0.115 $Y=0.234
c70 47 VSS 0.00906573f $X=0.216 $Y=0.216
c71 43 VSS 5.54432e-19 $X=0.233 $Y=0.216
c72 42 VSS 0.00827708f $X=0.108 $Y=0.216
c73 38 VSS 5.65078e-19 $X=0.125 $Y=0.216
c74 37 VSS 0.00481009f $X=0.162 $Y=0.0675
c75 33 VSS 7.28464e-19 $X=0.179 $Y=0.0675
c76 29 VSS 0.0144554f $X=0.459 $Y=0.135
c77 26 VSS 0.0645347f $X=0.459 $Y=0.0675
c78 18 VSS 0.0644226f $X=0.405 $Y=0.0675
c79 10 VSS 0.0642127f $X=0.351 $Y=0.0675
c80 2 VSS 0.061136f $X=0.297 $Y=0.0675
r81 85 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.207 $Y2=0.234
r82 83 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.207 $Y2=0.234
r83 81 85 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.198 $Y2=0.234
r84 78 79 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.15 $X2=0.297 $Y2=0.166
r85 75 78 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.15
r86 73 79 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.182 $X2=0.297 $Y2=0.166
r87 71 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.191 $X2=0.27 $Y2=0.191
r88 70 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.191 $X2=0.252 $Y2=0.191
r89 69 70 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.231
+ $Y=0.191 $X2=0.234 $Y2=0.191
r90 68 80 0.134501 $w=3.6e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.191 $X2=0.1885 $Y2=0.191
r91 68 69 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.191 $X2=0.231 $Y2=0.191
r92 67 73 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.191 $X2=0.297 $Y2=0.182
r93 67 72 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.191 $X2=0.27 $Y2=0.191
r94 66 81 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.234
r95 65 80 0.517544 $w=1.8e-08 $l=9.24662e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.2 $X2=0.1885 $Y2=0.191
r96 65 66 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.2 $X2=0.189 $Y2=0.225
r97 63 64 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.107 $X2=0.189 $Y2=0.15
r98 62 80 0.517544 $w=1.8e-08 $l=9.24662e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.182 $X2=0.1885 $Y2=0.191
r99 62 64 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.182 $X2=0.189 $Y2=0.15
r100 61 63 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.082 $X2=0.189 $Y2=0.107
r101 57 61 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.073 $X2=0.189 $Y2=0.082
r102 57 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.073 $X2=0.162 $Y2=0.073
r103 55 56 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.179 $Y2=0.234
r104 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r105 53 54 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.115
+ $Y=0.234 $X2=0.126 $Y2=0.234
r106 50 53 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.115 $Y2=0.234
r107 48 81 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.189 $Y2=0.234
r108 48 56 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.179 $Y2=0.234
r109 47 83 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r110 44 47 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.216 $X2=0.216 $Y2=0.216
r111 43 47 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.216 $X2=0.216 $Y2=0.216
r112 42 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r113 39 42 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.216 $X2=0.108 $Y2=0.216
r114 38 42 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.216 $X2=0.108 $Y2=0.216
r115 37 59 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.073
+ $X2=0.162 $Y2=0.073
r116 34 37 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r117 33 37 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r118 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r119 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r120 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r121 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r122 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r123 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r124 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r125 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r126 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r127 5 75 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r128 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r129 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AND2X4_ASAP7_75T_R%Y 1 2 6 7 11 12 15 16 17 20 21 24 28 29 40 42 VSS
c20 44 VSS 7.14098e-19 $X=0.513 $Y=0.2125
c21 42 VSS 8.03494e-19 $X=0.513 $Y=0.13425
c22 41 VSS 0.00497692f $X=0.513 $Y=0.121
c23 40 VSS 0.00419348f $X=0.5115 $Y=0.1475
c24 38 VSS 6.07272e-19 $X=0.513 $Y=0.225
c25 29 VSS 0.0266017f $X=0.504 $Y=0.234
c26 28 VSS 0.0092975f $X=0.432 $Y=0.036
c27 24 VSS 0.00913302f $X=0.324 $Y=0.036
c28 21 VSS 0.0265191f $X=0.504 $Y=0.036
c29 20 VSS 0.00929709f $X=0.432 $Y=0.2025
c30 16 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c31 15 VSS 0.010224f $X=0.324 $Y=0.2025
c32 11 VSS 5.72268e-19 $X=0.341 $Y=0.2025
c33 6 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c34 1 VSS 5.72268e-19 $X=0.341 $Y=0.0675
r35 43 44 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.2 $X2=0.513 $Y2=0.2125
r36 41 42 0.899691 $w=1.8e-08 $l=1.325e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.121 $X2=0.513 $Y2=0.13425
r37 40 43 3.56481 $w=1.8e-08 $l=5.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.1475 $X2=0.513 $Y2=0.2
r38 40 42 0.899691 $w=1.8e-08 $l=1.325e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.1475 $X2=0.513 $Y2=0.13425
r39 38 44 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.225 $X2=0.513 $Y2=0.2125
r40 37 41 5.16049 $w=1.8e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.045 $X2=0.513 $Y2=0.121
r41 31 35 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r42 29 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.234 $X2=0.513 $Y2=0.225
r43 29 35 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.432 $Y2=0.234
r44 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r45 23 27 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r46 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r47 21 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.504 $Y=0.036 $X2=0.513 $Y2=0.045
r48 21 27 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.432 $Y2=0.036
r49 20 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r50 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r51 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r52 15 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r53 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r54 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r55 10 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r56 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r57 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r58 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r59 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.324 $Y2=0.0675
r60 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.0675 $X2=0.324 $Y2=0.0675
.ends

.subckt PM_AND2X4_ASAP7_75T_R%7 1 2 VSS
c1 1 VSS 0.00241777f $X=0.125 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends

.subckt PM_AND2X4_ASAP7_75T_R%8 1 2 VSS
c0 1 VSS 0.00246714f $X=0.233 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.199 $Y2=0.0675
.ends


* END of "./AND2x4_ASAP7_75t_R.pex.sp.pex"
* 
.subckt AND2x4_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 VSS N_A_M0_g N_7_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_7_M1_d N_B_M1_g N_5_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_8_M2_d N_B_M2_g N_5_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_A_M3_g N_8_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_5_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_5_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_5_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_5_M7_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_5_M8_d N_A_M8_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M9 VDD N_B_M9_g N_5_M9_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
M10 VDD N_B_M10_g N_5_M10_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M11 N_5_M11_d N_A_M11_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M12 N_Y_M12_d N_5_M12_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M13 N_Y_M13_d N_5_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M14 N_Y_M14_d N_5_M14_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M15 N_Y_M15_d N_5_M15_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "AND2x4_ASAP7_75t_R.pex.sp.AND2X4_ASAP7_75T_R.pxi"
* BEGIN of "./AND2x4_ASAP7_75t_R.pex.sp.AND2X4_ASAP7_75T_R.pxi"
* File: AND2x4_ASAP7_75t_R.pex.sp.AND2X4_ASAP7_75T_R.pxi
* Created: Tue Sep  5 11:59:04 2017
* 
x_PM_AND2X4_ASAP7_75T_R%A N_A_M0_g N_A_c_7_p N_A_M8_g N_A_M3_g N_A_c_8_p
+ N_A_M11_g N_A_c_14_p N_A_c_19_p N_A_c_15_p N_A_c_9_p A N_A_c_27_p N_A_c_3_p
+ N_A_c_23_p N_A_c_17_p N_A_c_21_p VSS PM_AND2X4_ASAP7_75T_R%A
x_PM_AND2X4_ASAP7_75T_R%B N_B_M1_g N_B_M9_g N_B_M2_g N_B_c_34_n N_B_M10_g
+ N_B_c_36_n B VSS PM_AND2X4_ASAP7_75T_R%B
x_PM_AND2X4_ASAP7_75T_R%5 N_5_M4_g N_5_M12_g N_5_M5_g N_5_M13_g N_5_M6_g
+ N_5_M14_g N_5_M7_g N_5_c_53_n N_5_M15_g N_5_M2_s N_5_M1_s N_5_c_54_n N_5_M9_s
+ N_5_M8_d N_5_c_58_n N_5_M11_d N_5_M10_s N_5_c_71_n N_5_c_73_n N_5_c_59_n
+ N_5_c_62_n N_5_c_77_n N_5_c_64_n N_5_c_66_n N_5_c_84_p N_5_c_79_n N_5_c_97_p
+ VSS PM_AND2X4_ASAP7_75T_R%5
x_PM_AND2X4_ASAP7_75T_R%Y N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M6_d N_Y_M13_d
+ N_Y_M12_d N_Y_c_104_n N_Y_M15_d N_Y_M14_d N_Y_c_107_n N_Y_c_100_n N_Y_c_112_n
+ N_Y_c_113_n N_Y_c_114_n Y N_Y_c_119_n VSS PM_AND2X4_ASAP7_75T_R%Y
x_PM_AND2X4_ASAP7_75T_R%7 N_7_M1_d N_7_M0_s VSS PM_AND2X4_ASAP7_75T_R%7
x_PM_AND2X4_ASAP7_75T_R%8 N_8_M3_s N_8_M2_d VSS PM_AND2X4_ASAP7_75T_R%8
cc_1 N_A_M0_g N_B_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_M3_g N_B_M1_g 2.66145e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_3 N_A_c_3_p N_B_M1_g 2.41954e-19 $X=0.198 $Y=0.037 $X2=0.135 $Y2=0.0675
cc_4 N_A_M0_g N_B_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_5 N_A_M3_g N_B_M2_g 0.00343649f $X=0.243 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_6 N_A_c_3_p N_B_M2_g 2.38593e-19 $X=0.198 $Y=0.037 $X2=0.189 $Y2=0.0675
cc_7 N_A_c_7_p N_B_c_34_n 7.92842e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_8 N_A_c_8_p N_B_c_34_n 7.27564e-19 $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.135
cc_9 N_A_c_9_p N_B_c_36_n 0.00216743f $X=0.081 $Y=0.121 $X2=0.135 $Y2=0.135
cc_10 A B 0.00216743f $X=0.083 $Y=0.14 $X2=0.135 $Y2=0.152
cc_11 N_A_M3_g N_5_M4_g 0.00287344f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_12 N_A_M3_g N_5_M5_g 2.34385e-19 $X=0.243 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_13 N_A_c_8_p N_5_c_53_n 7.99973e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_14 N_A_c_14_p N_5_c_54_n 3.16725e-19 $X=0.081 $Y=0.064 $X2=0 $Y2=0
cc_15 N_A_c_15_p N_5_c_54_n 3.81105e-19 $X=0.081 $Y=0.107 $X2=0 $Y2=0
cc_16 N_A_c_3_p N_5_c_54_n 0.00275621f $X=0.198 $Y=0.037 $X2=0 $Y2=0
cc_17 N_A_c_17_p N_5_c_54_n 3.16725e-19 $X=0.243 $Y=0.064 $X2=0 $Y2=0
cc_18 A N_5_c_58_n 3.31541e-19 $X=0.083 $Y=0.14 $X2=0 $Y2=0
cc_19 N_A_c_19_p N_5_c_59_n 0.00124379f $X=0.081 $Y=0.082 $X2=0 $Y2=0
cc_20 N_A_c_3_p N_5_c_59_n 0.00767084f $X=0.198 $Y=0.037 $X2=0 $Y2=0
cc_21 N_A_c_21_p N_5_c_59_n 0.00191714f $X=0.243 $Y=0.121 $X2=0 $Y2=0
cc_22 N_A_c_15_p N_5_c_62_n 2.64182e-19 $X=0.081 $Y=0.107 $X2=0 $Y2=0
cc_23 N_A_c_23_p N_5_c_62_n 0.00191714f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_24 N_A_M3_g N_5_c_64_n 3.8173e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_25 N_A_c_23_p N_5_c_64_n 9.6052e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_26 N_A_c_23_p N_5_c_66_n 0.00122369f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_27 N_A_c_27_p N_Y_c_100_n 4.60508e-19 $X=0.234 $Y=0.037 $X2=0.135 $Y2=0.152
cc_28 N_B_M2_g N_5_M4_g 2.31381e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_29 N_B_c_34_n N_5_M2_s 3.53813e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.046
cc_30 N_B_c_34_n N_5_c_54_n 8.23937e-19 $X=0.189 $Y=0.135 $X2=0.243 $Y2=0.064
cc_31 B N_5_c_58_n 3.31541e-19 $X=0.135 $Y=0.152 $X2=0 $Y2=0
cc_32 N_B_M1_g N_5_c_71_n 2.57565e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_33 B N_5_c_71_n 0.00123074f $X=0.135 $Y=0.152 $X2=0 $Y2=0
cc_34 N_B_c_34_n N_5_c_73_n 5.63985e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_35 N_B_M1_g N_5_c_59_n 2.75912e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B_c_34_n N_5_c_59_n 6.27351e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_37 N_B_c_36_n N_5_c_59_n 0.00123355f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_38 N_B_c_34_n N_5_c_77_n 0.00202781f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_39 N_B_c_36_n N_5_c_77_n 0.00362836f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_40 B N_5_c_79_n 8.62553e-19 $X=0.135 $Y=0.152 $X2=0 $Y2=0
cc_41 N_5_c_53_n N_Y_M5_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_42 N_5_c_53_n N_Y_M7_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.216
cc_43 N_5_c_53_n N_Y_M13_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_44 N_5_c_53_n N_Y_c_104_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.216
cc_45 N_5_c_84_p N_Y_c_104_n 0.00134951f $X=0.297 $Y=0.166 $X2=0.243 $Y2=0.216
cc_46 N_5_c_53_n N_Y_M15_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_47 N_5_c_53_n N_Y_c_107_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.135
cc_48 N_5_M5_g N_Y_c_100_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.064
cc_49 N_5_M6_g N_Y_c_100_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.064
cc_50 N_5_M7_g N_Y_c_100_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.064
cc_51 N_5_c_53_n N_Y_c_100_n 0.00191346f $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.064
cc_52 N_5_c_53_n N_Y_c_112_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.121
cc_53 N_5_c_53_n N_Y_c_113_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.09 $Y2=0.037
cc_54 N_5_M5_g N_Y_c_114_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.094 $Y2=0.037
cc_55 N_5_M6_g N_Y_c_114_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0.094 $Y2=0.037
cc_56 N_5_M7_g N_Y_c_114_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.094 $Y2=0.037
cc_57 N_5_c_53_n N_Y_c_114_n 0.00191346f $X=0.459 $Y=0.135 $X2=0.094 $Y2=0.037
cc_58 N_5_c_97_p N_Y_c_114_n 3.03775e-19 $X=0.216 $Y=0.234 $X2=0.094 $Y2=0.037
cc_59 N_5_c_53_n N_Y_c_119_n 4.05816e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_60 N_5_c_59_n N_7_M1_d 2.13297e-19 $X=0.18 $Y=0.073 $X2=0.081 $Y2=0.0675

* END of "./AND2x4_ASAP7_75t_R.pex.sp.AND2X4_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: AND2x6_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 11:59:27 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AND2x6_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./AND2x6_ASAP7_75t_R.pex.sp.pex"
* File: AND2x6_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 11:59:27 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AND2X6_ASAP7_75T_R%A 2 5 7 10 13 15 21 22 23 24 25 27 31 35 37 38 VSS
c27 38 VSS 0.00255655f $X=0.243 $Y=0.121
c28 37 VSS 8.45284e-19 $X=0.243 $Y=0.064
c29 35 VSS 2.3666e-19 $X=0.243 $Y=0.135
c30 32 VSS 0.00189145f $X=0.216 $Y=0.037
c31 31 VSS 0.00636831f $X=0.198 $Y=0.037
c32 30 VSS 0.00199175f $X=0.115 $Y=0.037
c33 29 VSS 3.03073e-19 $X=0.094 $Y=0.037
c34 28 VSS 0.0030786f $X=0.09 $Y=0.037
c35 27 VSS 0.00438018f $X=0.234 $Y=0.037
c36 25 VSS 0.00242134f $X=0.083 $Y=0.14
c37 24 VSS 3.59668e-19 $X=0.081 $Y=0.121
c38 23 VSS 0.0011834f $X=0.081 $Y=0.107
c39 22 VSS 9.44831e-19 $X=0.081 $Y=0.082
c40 21 VSS 8.45284e-19 $X=0.081 $Y=0.064
c41 13 VSS 9.42534e-19 $X=0.243 $Y=0.135
c42 10 VSS 0.059423f $X=0.243 $Y=0.0675
c43 5 VSS 0.00198216f $X=0.081 $Y=0.135
c44 2 VSS 0.0627695f $X=0.081 $Y=0.0675
r45 37 38 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.064 $X2=0.243 $Y2=0.121
r46 35 38 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.121
r47 33 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.046 $X2=0.243 $Y2=0.064
r48 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.037 $X2=0.216 $Y2=0.037
r49 30 31 5.6358 $w=1.8e-08 $l=8.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.115
+ $Y=0.037 $X2=0.198 $Y2=0.037
r50 29 30 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.037 $X2=0.115 $Y2=0.037
r51 28 29 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.037 $X2=0.094 $Y2=0.037
r52 27 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.037 $X2=0.243 $Y2=0.046
r53 27 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.037 $X2=0.216 $Y2=0.037
r54 24 25 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.121 $X2=0.081 $Y2=0.135
r55 23 24 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.107 $X2=0.081 $Y2=0.121
r56 22 23 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.082 $X2=0.081 $Y2=0.107
r57 21 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.064 $X2=0.081 $Y2=0.082
r58 17 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.046 $X2=0.09 $Y2=0.037
r59 17 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.046 $X2=0.081 $Y2=0.064
r60 13 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r61 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.216
r62 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r63 5 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r64 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r65 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AND2X6_ASAP7_75T_R%B 2 7 10 13 15 18 22 VSS
c23 22 VSS 4.12915e-19 $X=0.135 $Y=0.152
c24 18 VSS 4.05597e-19 $X=0.135 $Y=0.135
c25 13 VSS 0.00443484f $X=0.189 $Y=0.135
c26 10 VSS 0.0626014f $X=0.189 $Y=0.0675
c27 2 VSS 0.0615487f $X=0.135 $Y=0.0675
r28 18 22 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.152
r29 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.216
r30 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r31 5 13 60 $w=1.8e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135 $Y=0.135
+ $X2=0.189 $Y2=0.135
r32 5 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r33 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r34 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AND2X6_ASAP7_75T_R%5 2 7 10 15 18 23 26 31 34 39 42 45 47 49 50 53 54
+ 55 58 59 60 71 72 73 79 80 87 91 95 96 99 VSS
c57 102 VSS 6.58501e-19 $X=0.207 $Y=0.234
c58 101 VSS 0.00176786f $X=0.198 $Y=0.234
c59 99 VSS 0.00285708f $X=0.216 $Y=0.234
c60 96 VSS 4.93096e-19 $X=0.1885 $Y=0.191
c61 95 VSS 5.11872e-19 $X=0.297 $Y=0.166
c62 91 VSS 5.49936e-19 $X=0.297 $Y=0.135
c63 89 VSS 6.27562e-19 $X=0.297 $Y=0.182
c64 88 VSS 0.00254231f $X=0.27 $Y=0.191
c65 87 VSS 4.66176e-19 $X=0.252 $Y=0.191
c66 86 VSS 1.69914e-19 $X=0.234 $Y=0.191
c67 85 VSS 6.30164e-19 $X=0.231 $Y=0.191
c68 83 VSS 0.00194692f $X=0.288 $Y=0.191
c69 82 VSS 0.00121124f $X=0.189 $Y=0.225
c70 80 VSS 2.55645e-19 $X=0.189 $Y=0.15
c71 79 VSS 6.49295e-20 $X=0.189 $Y=0.107
c72 78 VSS 5.03482e-19 $X=0.189 $Y=0.182
c73 73 VSS 9.05837e-19 $X=0.18 $Y=0.073
c74 72 VSS 0.0053518f $X=0.179 $Y=0.234
c75 71 VSS 0.00142296f $X=0.144 $Y=0.234
c76 70 VSS 0.00105114f $X=0.126 $Y=0.234
c77 69 VSS 0.00346796f $X=0.115 $Y=0.234
c78 63 VSS 0.00906573f $X=0.216 $Y=0.216
c79 59 VSS 5.54432e-19 $X=0.233 $Y=0.216
c80 58 VSS 0.00827708f $X=0.108 $Y=0.216
c81 54 VSS 5.65078e-19 $X=0.125 $Y=0.216
c82 53 VSS 0.00481009f $X=0.162 $Y=0.0675
c83 49 VSS 7.28464e-19 $X=0.179 $Y=0.0675
c84 45 VSS 0.0249841f $X=0.567 $Y=0.135
c85 42 VSS 0.0645347f $X=0.567 $Y=0.0675
c86 34 VSS 0.0644226f $X=0.513 $Y=0.0675
c87 26 VSS 0.0642127f $X=0.459 $Y=0.0675
c88 18 VSS 0.0642127f $X=0.405 $Y=0.0675
c89 10 VSS 0.0642127f $X=0.351 $Y=0.0675
c90 2 VSS 0.061136f $X=0.297 $Y=0.0675
r91 101 102 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.207 $Y2=0.234
r92 99 102 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.207 $Y2=0.234
r93 97 101 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.234 $X2=0.198 $Y2=0.234
r94 94 95 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.15 $X2=0.297 $Y2=0.166
r95 91 94 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.15
r96 89 95 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.182 $X2=0.297 $Y2=0.166
r97 87 88 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.191 $X2=0.27 $Y2=0.191
r98 86 87 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.191 $X2=0.252 $Y2=0.191
r99 85 86 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.231
+ $Y=0.191 $X2=0.234 $Y2=0.191
r100 84 96 0.134501 $w=3.6e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.191 $X2=0.1885 $Y2=0.191
r101 84 85 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.191 $X2=0.231 $Y2=0.191
r102 83 89 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.191 $X2=0.297 $Y2=0.182
r103 83 88 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.191 $X2=0.27 $Y2=0.191
r104 82 97 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.225 $X2=0.189 $Y2=0.234
r105 81 96 0.517544 $w=1.8e-08 $l=9.24662e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.2 $X2=0.1885 $Y2=0.191
r106 81 82 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.2 $X2=0.189 $Y2=0.225
r107 79 80 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.107 $X2=0.189 $Y2=0.15
r108 78 96 0.517544 $w=1.8e-08 $l=9.24662e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.182 $X2=0.1885 $Y2=0.191
r109 78 80 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.182 $X2=0.189 $Y2=0.15
r110 77 79 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.082 $X2=0.189 $Y2=0.107
r111 73 77 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.073 $X2=0.189 $Y2=0.082
r112 73 75 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.073 $X2=0.162 $Y2=0.073
r113 71 72 2.37654 $w=1.8e-08 $l=3.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.179 $Y2=0.234
r114 70 71 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r115 69 70 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.115
+ $Y=0.234 $X2=0.126 $Y2=0.234
r116 66 69 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.115 $Y2=0.234
r117 64 97 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.189 $Y2=0.234
r118 64 72 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.179 $Y2=0.234
r119 63 99 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r120 60 63 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.216 $X2=0.216 $Y2=0.216
r121 59 63 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.216 $X2=0.216 $Y2=0.216
r122 58 66 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r123 55 58 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.216 $X2=0.108 $Y2=0.216
r124 54 58 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.216 $X2=0.108 $Y2=0.216
r125 53 75 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.073
+ $X2=0.162 $Y2=0.073
r126 50 53 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r127 49 53 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r128 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.135 $X2=0.567 $Y2=0.2025
r129 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.0675 $X2=0.567 $Y2=0.135
r130 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r131 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r132 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r133 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r134 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r135 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r136 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r137 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r138 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r139 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r140 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r141 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r142 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r143 5 91 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r144 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r145 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AND2X6_ASAP7_75T_R%Y 1 2 6 7 11 12 16 17 20 21 22 25 26 27 30 31 34
+ 38 41 42 56 58 VSS
c28 60 VSS 7.14098e-19 $X=0.621 $Y=0.2125
c29 58 VSS 6.63487e-19 $X=0.621 $Y=0.13425
c30 57 VSS 0.00497692f $X=0.621 $Y=0.121
c31 56 VSS 0.00432017f $X=0.6195 $Y=0.1475
c32 54 VSS 6.07272e-19 $X=0.621 $Y=0.225
c33 42 VSS 0.0385606f $X=0.612 $Y=0.234
c34 41 VSS 0.00929752f $X=0.54 $Y=0.036
c35 38 VSS 0.00928951f $X=0.432 $Y=0.036
c36 34 VSS 0.00913304f $X=0.324 $Y=0.036
c37 31 VSS 0.0384777f $X=0.612 $Y=0.036
c38 30 VSS 0.00929752f $X=0.54 $Y=0.2025
c39 26 VSS 5.38922e-19 $X=0.557 $Y=0.2025
c40 25 VSS 0.0092891f $X=0.432 $Y=0.2025
c41 21 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c42 20 VSS 0.010224f $X=0.324 $Y=0.2025
c43 16 VSS 5.72268e-19 $X=0.341 $Y=0.2025
c44 11 VSS 5.38922e-19 $X=0.557 $Y=0.0675
c45 6 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c46 1 VSS 5.72268e-19 $X=0.341 $Y=0.0675
r47 59 60 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.2 $X2=0.621 $Y2=0.2125
r48 57 58 0.899691 $w=1.8e-08 $l=1.325e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.121 $X2=0.621 $Y2=0.13425
r49 56 59 3.56481 $w=1.8e-08 $l=5.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.1475 $X2=0.621 $Y2=0.2
r50 56 58 0.899691 $w=1.8e-08 $l=1.325e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.1475 $X2=0.621 $Y2=0.13425
r51 54 60 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.2125
r52 53 57 5.16049 $w=1.8e-08 $l=7.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.121
r53 48 51 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.54 $Y2=0.234
r54 44 48 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r55 42 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r56 42 51 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.54 $Y2=0.234
r57 40 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r58 37 40 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.54 $Y2=0.036
r59 37 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r60 33 37 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r61 33 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r62 31 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r63 31 40 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.54 $Y2=0.036
r64 30 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r65 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r66 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r67 25 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r68 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r69 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r70 20 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r71 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r72 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r73 15 41 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r74 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r75 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r76 10 38 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r77 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r78 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r79 5 34 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r80 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.324 $Y2=0.0675
r81 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.0675 $X2=0.324 $Y2=0.0675
.ends

.subckt PM_AND2X6_ASAP7_75T_R%7 1 2 VSS
c1 1 VSS 0.00241777f $X=0.125 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends

.subckt PM_AND2X6_ASAP7_75T_R%8 1 2 VSS
c0 1 VSS 0.00246714f $X=0.233 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.199 $Y2=0.0675
.ends


* END of "./AND2x6_ASAP7_75t_R.pex.sp.pex"
* 
.subckt AND2x6_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 VSS N_A_M0_g N_7_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_7_M1_d N_B_M1_g N_5_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_8_M2_d N_B_M2_g N_5_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_A_M3_g N_8_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_5_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_5_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_5_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_5_M7_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_5_M8_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_5_M9_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 N_5_M10_d N_A_M10_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M11 VDD N_B_M11_g N_5_M11_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M12 VDD N_B_M12_g N_5_M12_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179
+ $Y=0.189
M13 N_5_M13_d N_A_M13_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233
+ $Y=0.189
M14 N_Y_M14_d N_5_M14_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M15 N_Y_M15_d N_5_M15_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M16 N_Y_M16_d N_5_M16_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M17 N_Y_M17_d N_5_M17_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M18 N_Y_M18_d N_5_M18_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M19 N_Y_M19_d N_5_M19_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
*
* 
* .include "AND2x6_ASAP7_75t_R.pex.sp.AND2X6_ASAP7_75T_R.pxi"
* BEGIN of "./AND2x6_ASAP7_75t_R.pex.sp.AND2X6_ASAP7_75T_R.pxi"
* File: AND2x6_ASAP7_75t_R.pex.sp.AND2X6_ASAP7_75T_R.pxi
* Created: Tue Sep  5 11:59:27 2017
* 
x_PM_AND2X6_ASAP7_75T_R%A N_A_M0_g N_A_c_7_p N_A_M10_g N_A_M3_g N_A_c_8_p
+ N_A_M13_g N_A_c_14_p N_A_c_19_p N_A_c_15_p N_A_c_9_p A N_A_c_27_p N_A_c_3_p
+ N_A_c_23_p N_A_c_17_p N_A_c_21_p VSS PM_AND2X6_ASAP7_75T_R%A
x_PM_AND2X6_ASAP7_75T_R%B N_B_M1_g N_B_M11_g N_B_M2_g N_B_c_34_n N_B_M12_g
+ N_B_c_36_n B VSS PM_AND2X6_ASAP7_75T_R%B
x_PM_AND2X6_ASAP7_75T_R%5 N_5_M4_g N_5_M14_g N_5_M5_g N_5_M15_g N_5_M6_g
+ N_5_M16_g N_5_M7_g N_5_M17_g N_5_M8_g N_5_M18_g N_5_M9_g N_5_c_53_n N_5_M19_g
+ N_5_M2_s N_5_M1_s N_5_c_54_n N_5_M11_s N_5_M10_d N_5_c_58_n N_5_M13_d
+ N_5_M12_s N_5_c_71_n N_5_c_73_n N_5_c_59_n N_5_c_62_n N_5_c_77_n N_5_c_64_n
+ N_5_c_66_n N_5_c_85_p N_5_c_79_n N_5_c_105_p VSS PM_AND2X6_ASAP7_75T_R%5
x_PM_AND2X6_ASAP7_75T_R%Y N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M6_d N_Y_M9_d N_Y_M8_d
+ N_Y_M15_d N_Y_M14_d N_Y_c_113_n N_Y_M17_d N_Y_M16_d N_Y_c_116_n N_Y_M19_d
+ N_Y_M18_d N_Y_c_118_n N_Y_c_108_n N_Y_c_125_n N_Y_c_126_n N_Y_c_127_n
+ N_Y_c_128_n Y N_Y_c_135_n VSS PM_AND2X6_ASAP7_75T_R%Y
x_PM_AND2X6_ASAP7_75T_R%7 N_7_M1_d N_7_M0_s VSS PM_AND2X6_ASAP7_75T_R%7
x_PM_AND2X6_ASAP7_75T_R%8 N_8_M3_s N_8_M2_d VSS PM_AND2X6_ASAP7_75T_R%8
cc_1 N_A_M0_g N_B_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_M3_g N_B_M1_g 2.66145e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_3 N_A_c_3_p N_B_M1_g 2.41954e-19 $X=0.198 $Y=0.037 $X2=0.135 $Y2=0.0675
cc_4 N_A_M0_g N_B_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_5 N_A_M3_g N_B_M2_g 0.00343649f $X=0.243 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_6 N_A_c_3_p N_B_M2_g 2.38593e-19 $X=0.198 $Y=0.037 $X2=0.189 $Y2=0.0675
cc_7 N_A_c_7_p N_B_c_34_n 7.92842e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_8 N_A_c_8_p N_B_c_34_n 7.27564e-19 $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.135
cc_9 N_A_c_9_p N_B_c_36_n 0.00216743f $X=0.081 $Y=0.121 $X2=0.135 $Y2=0.135
cc_10 A B 0.00216743f $X=0.083 $Y=0.14 $X2=0.135 $Y2=0.152
cc_11 N_A_M3_g N_5_M4_g 0.00287344f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_12 N_A_M3_g N_5_M5_g 2.34385e-19 $X=0.243 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_13 N_A_c_8_p N_5_c_53_n 8.00951e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_14 N_A_c_14_p N_5_c_54_n 3.16725e-19 $X=0.081 $Y=0.064 $X2=0 $Y2=0
cc_15 N_A_c_15_p N_5_c_54_n 3.81105e-19 $X=0.081 $Y=0.107 $X2=0 $Y2=0
cc_16 N_A_c_3_p N_5_c_54_n 0.00275621f $X=0.198 $Y=0.037 $X2=0 $Y2=0
cc_17 N_A_c_17_p N_5_c_54_n 3.16725e-19 $X=0.243 $Y=0.064 $X2=0 $Y2=0
cc_18 A N_5_c_58_n 3.31541e-19 $X=0.083 $Y=0.14 $X2=0 $Y2=0
cc_19 N_A_c_19_p N_5_c_59_n 0.00124379f $X=0.081 $Y=0.082 $X2=0 $Y2=0
cc_20 N_A_c_3_p N_5_c_59_n 0.00767084f $X=0.198 $Y=0.037 $X2=0 $Y2=0
cc_21 N_A_c_21_p N_5_c_59_n 0.00191714f $X=0.243 $Y=0.121 $X2=0 $Y2=0
cc_22 N_A_c_15_p N_5_c_62_n 2.64182e-19 $X=0.081 $Y=0.107 $X2=0 $Y2=0
cc_23 N_A_c_23_p N_5_c_62_n 0.00191714f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_24 N_A_M3_g N_5_c_64_n 3.8173e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_25 N_A_c_23_p N_5_c_64_n 9.6052e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_26 N_A_c_23_p N_5_c_66_n 0.00122369f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_27 N_A_c_27_p N_Y_c_108_n 4.70766e-19 $X=0.234 $Y=0.037 $X2=0 $Y2=0
cc_28 N_B_M2_g N_5_M4_g 2.31381e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_29 N_B_c_34_n N_5_M2_s 3.53813e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_30 N_B_c_34_n N_5_c_54_n 8.23937e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_31 B N_5_c_58_n 3.31541e-19 $X=0.135 $Y=0.152 $X2=0 $Y2=0
cc_32 N_B_M1_g N_5_c_71_n 2.57565e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_33 B N_5_c_71_n 0.00123074f $X=0.135 $Y=0.152 $X2=0 $Y2=0
cc_34 N_B_c_34_n N_5_c_73_n 5.63985e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_35 N_B_M1_g N_5_c_59_n 2.75912e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B_c_34_n N_5_c_59_n 6.27351e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_37 N_B_c_36_n N_5_c_59_n 0.00123355f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_38 N_B_c_34_n N_5_c_77_n 0.00202781f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_39 N_B_c_36_n N_5_c_77_n 0.00362836f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_40 B N_5_c_79_n 8.62553e-19 $X=0.135 $Y=0.152 $X2=0 $Y2=0
cc_41 N_5_c_53_n N_Y_M5_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_42 N_5_c_53_n N_Y_M7_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.216
cc_43 N_5_c_53_n N_Y_M9_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_44 N_5_c_53_n N_Y_M15_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_45 N_5_c_53_n N_Y_c_113_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.135
cc_46 N_5_c_85_p N_Y_c_113_n 6.96092e-19 $X=0.297 $Y=0.166 $X2=0.081 $Y2=0.135
cc_47 N_5_c_53_n N_Y_M17_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.064
cc_48 N_5_c_53_n N_Y_c_116_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0.083 $Y2=0.14
cc_49 N_5_c_53_n N_Y_M19_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_50 N_5_c_53_n N_Y_c_118_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0.115 $Y2=0.037
cc_51 N_5_M5_g N_Y_c_108_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.198 $Y2=0.037
cc_52 N_5_M6_g N_Y_c_108_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0.198 $Y2=0.037
cc_53 N_5_M7_g N_Y_c_108_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.198 $Y2=0.037
cc_54 N_5_M8_g N_Y_c_108_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.198 $Y2=0.037
cc_55 N_5_M9_g N_Y_c_108_n 4.59284e-19 $X=0.567 $Y=0.0675 $X2=0.198 $Y2=0.037
cc_56 N_5_c_53_n N_Y_c_108_n 0.00327571f $X=0.567 $Y=0.135 $X2=0.198 $Y2=0.037
cc_57 N_5_c_53_n N_Y_c_125_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0.243 $Y2=0.135
cc_58 N_5_c_53_n N_Y_c_126_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0.243 $Y2=0.121
cc_59 N_5_c_53_n N_Y_c_127_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_60 N_5_M5_g N_Y_c_128_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_61 N_5_M6_g N_Y_c_128_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_62 N_5_M7_g N_Y_c_128_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_63 N_5_M8_g N_Y_c_128_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_5_M9_g N_Y_c_128_n 4.59284e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_65 N_5_c_53_n N_Y_c_128_n 0.00327571f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_66 N_5_c_105_p N_Y_c_128_n 3.10557e-19 $X=0.216 $Y=0.234 $X2=0 $Y2=0
cc_67 N_5_c_53_n N_Y_c_135_n 0.00101053f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_68 N_5_c_59_n N_7_M1_d 2.13297e-19 $X=0.18 $Y=0.073 $X2=0.081 $Y2=0.0675

* END of "./AND2x6_ASAP7_75t_R.pex.sp.AND2X6_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: AND3x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 11:59:49 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AND3x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./AND3x1_ASAP7_75t_R.pex.sp.pex"
* File: AND3x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 11:59:49 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AND3X1_ASAP7_75T_R%A 2 5 7 18 21 24 VSS
c11 24 VSS 0.0086019f $X=0.019 $Y=0.137
c12 21 VSS 5.05467e-19 $X=0.0605 $Y=0.135
c13 20 VSS 0.00132257f $X=0.04 $Y=0.135
c14 18 VSS 5.84838e-19 $X=0.081 $Y=0.135
c15 5 VSS 0.00271097f $X=0.081 $Y=0.135
c16 2 VSS 0.0654968f $X=0.081 $Y=0.0675
r17 20 21 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.135 $X2=0.0605 $Y2=0.135
r18 18 21 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0605 $Y2=0.135
r19 16 24 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r20 16 20 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.04 $Y2=0.135
r21 5 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AND3X1_ASAP7_75T_R%B 2 5 7 13 VSS
c14 13 VSS 0.00201056f $X=0.138 $Y=0.137
c15 5 VSS 0.00101978f $X=0.135 $Y=0.135
c16 2 VSS 0.0597337f $X=0.135 $Y=0.0675
r17 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AND3X1_ASAP7_75T_R%C 2 5 7 13 VSS
c12 13 VSS 0.00121916f $X=0.189 $Y=0.137
c13 5 VSS 0.00108616f $X=0.189 $Y=0.135
c14 2 VSS 0.0591532f $X=0.189 $Y=0.0675
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AND3X1_ASAP7_75T_R%6 2 5 7 9 14 17 19 20 23 24 27 29 30 31 32 33 43
+ 45 48 52 53 54 57 58 64 VSS
c33 67 VSS 1.83894e-19 $X=0.241 $Y=0.135
c34 66 VSS 1.75358e-19 $X=0.234 $Y=0.135
c35 64 VSS 6.45658e-19 $X=0.248 $Y=0.135
c36 60 VSS 2.09895e-19 $X=0.225 $Y=0.216
c37 59 VSS 2.94089e-19 $X=0.225 $Y=0.207
c38 58 VSS 3.99142e-19 $X=0.225 $Y=0.2
c39 57 VSS 0.00108888f $X=0.225 $Y=0.183
c40 56 VSS 1.99485e-19 $X=0.225 $Y=0.225
c41 54 VSS 7.72566e-19 $X=0.225 $Y=0.11
c42 53 VSS 5.51756e-19 $X=0.225 $Y=0.094
c43 52 VSS 3.26372e-19 $X=0.225 $Y=0.07
c44 51 VSS 3.86867e-19 $X=0.225 $Y=0.063
c45 50 VSS 1.92199e-19 $X=0.225 $Y=0.126
c46 48 VSS 0.00146362f $X=0.198 $Y=0.234
c47 47 VSS 0.00258369f $X=0.18 $Y=0.234
c48 46 VSS 8.80294e-19 $X=0.153 $Y=0.234
c49 45 VSS 0.00142296f $X=0.144 $Y=0.234
c50 44 VSS 0.00558198f $X=0.126 $Y=0.234
c51 43 VSS 0.00574452f $X=0.095 $Y=0.234
c52 35 VSS 0.00574187f $X=0.216 $Y=0.234
c53 34 VSS 0.00191122f $X=0.207 $Y=0.036
c54 33 VSS 0.00142296f $X=0.198 $Y=0.036
c55 32 VSS 0.00333444f $X=0.18 $Y=0.036
c56 31 VSS 0.00142296f $X=0.144 $Y=0.036
c57 30 VSS 0.00312666f $X=0.126 $Y=0.036
c58 29 VSS 0.00574452f $X=0.095 $Y=0.036
c59 27 VSS 0.00240442f $X=0.054 $Y=0.036
c60 24 VSS 0.00421964f $X=0.216 $Y=0.036
c61 23 VSS 0.0105167f $X=0.162 $Y=0.2025
c62 19 VSS 5.38922e-19 $X=0.179 $Y=0.2025
c63 17 VSS 0.00568611f $X=0.056 $Y=0.2025
c64 14 VSS 3.33606e-19 $X=0.071 $Y=0.2025
c65 9 VSS 3.33606e-19 $X=0.071 $Y=0.0675
c66 5 VSS 0.00413468f $X=0.243 $Y=0.135
c67 2 VSS 0.0653057f $X=0.243 $Y=0.0675
r68 66 67 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.241 $Y2=0.135
r69 64 67 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.135 $X2=0.241 $Y2=0.135
r70 61 66 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.135 $X2=0.234 $Y2=0.135
r71 59 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.207 $X2=0.225 $Y2=0.216
r72 58 59 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.2 $X2=0.225 $Y2=0.207
r73 57 58 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.183 $X2=0.225 $Y2=0.2
r74 56 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.225 $X2=0.225 $Y2=0.216
r75 55 61 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.144 $X2=0.225 $Y2=0.135
r76 55 57 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.144 $X2=0.225 $Y2=0.183
r77 53 54 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.094 $X2=0.225 $Y2=0.11
r78 52 53 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.07 $X2=0.225 $Y2=0.094
r79 51 52 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.063 $X2=0.225 $Y2=0.07
r80 50 61 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r81 50 54 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.11
r82 49 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.063
r83 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r84 45 46 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.153 $Y2=0.234
r85 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r86 43 44 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.234 $X2=0.126 $Y2=0.234
r87 41 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r88 41 46 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.153 $Y2=0.234
r89 37 43 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.095 $Y2=0.234
r90 35 56 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.234 $X2=0.225 $Y2=0.225
r91 35 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.198 $Y2=0.234
r92 33 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.207 $Y2=0.036
r93 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r94 31 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.18 $Y2=0.036
r95 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r96 29 30 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.036 $X2=0.126 $Y2=0.036
r97 26 29 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.095 $Y2=0.036
r98 26 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r99 24 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.036 $X2=0.225 $Y2=0.045
r100 24 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.207 $Y2=0.036
r101 23 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r102 20 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r103 19 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r104 17 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r105 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r106 12 27 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.054 $Y=0.0675 $X2=0.054 $Y2=0.036
r107 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r108 5 64 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.248 $Y=0.135 $X2=0.248
+ $Y2=0.135
r109 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r110 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AND3X1_ASAP7_75T_R%Y 1 6 9 11 14 19 20 21 22 31 VSS
c10 31 VSS 0.00429788f $X=0.27 $Y=0.215
c11 28 VSS 3.40666e-19 $X=0.288 $Y=0.085
c12 27 VSS 5.60077e-20 $X=0.279 $Y=0.085
c13 26 VSS 0.00155357f $X=0.297 $Y=0.085
c14 22 VSS 1.78524e-19 $X=0.27 $Y=0.085
c15 21 VSS 7.16262e-19 $X=0.297 $Y=0.144
c16 20 VSS 0.00116892f $X=0.297 $Y=0.126
c17 19 VSS 0.00145955f $X=0.298 $Y=0.1475
c18 14 VSS 0.00555681f $X=0.27 $Y=0.048
c19 11 VSS 0.00234334f $X=0.27 $Y=0.076
c20 9 VSS 0.00620109f $X=0.268 $Y=0.2025
c21 4 VSS 5.08721e-19 $X=0.268 $Y=0.0675
r22 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.085 $X2=0.288 $Y2=0.085
r23 26 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.085 $X2=0.288 $Y2=0.085
r24 22 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.085 $X2=0.279 $Y2=0.085
r25 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.144
r26 19 21 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1475 $X2=0.297 $Y2=0.144
r27 17 31 1.04762 $w=3.15e-08 $l=4.65833e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.297 $Y=0.183 $X2=0.27 $Y2=0.218
r28 17 19 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.183 $X2=0.297 $Y2=0.1475
r29 16 26 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.094 $X2=0.297 $Y2=0.085
r30 16 20 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.094 $X2=0.297 $Y2=0.126
r31 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.048 $X2=0.27
+ $Y2=0.048
r32 11 22 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.076 $X2=0.27 $Y2=0.085
r33 11 13 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.076 $X2=0.27 $Y2=0.048
r34 9 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.215 $X2=0.27
+ $Y2=0.215
r35 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.2025 $X2=0.268 $Y2=0.2025
r36 4 14 16.8304 $w=2.4e-08 $l=1.95e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.048
r37 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.268 $Y2=0.0675
.ends

.subckt PM_AND3X1_ASAP7_75T_R%8 1 2 VSS
c1 1 VSS 0.00187952f $X=0.125 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends

.subckt PM_AND3X1_ASAP7_75T_R%9 1 2 VSS
c1 1 VSS 0.00183233f $X=0.179 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.145 $Y2=0.0675
.ends


* END of "./AND3x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt AND3x1_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 N_8_M0_d N_A_M0_g N_6_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_9_M1_d N_B_M1_g N_8_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_C_M2_g N_9_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_6_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 VDD N_A_M4_g N_6_M4_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M5 N_6_M5_d N_B_M5_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M6 VDD N_C_M6_g N_6_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M7 N_Y_M7_d N_6_M7_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
*
* 
* .include "AND3x1_ASAP7_75t_R.pex.sp.AND3X1_ASAP7_75T_R.pxi"
* BEGIN of "./AND3x1_ASAP7_75t_R.pex.sp.AND3X1_ASAP7_75T_R.pxi"
* File: AND3x1_ASAP7_75t_R.pex.sp.AND3X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 11:59:49 2017
* 
x_PM_AND3X1_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M4_g N_A_c_3_p N_A_c_9_p A VSS
+ PM_AND3X1_ASAP7_75T_R%A
x_PM_AND3X1_ASAP7_75T_R%B N_B_M1_g N_B_c_13_n N_B_M5_g B VSS
+ PM_AND3X1_ASAP7_75T_R%B
x_PM_AND3X1_ASAP7_75T_R%C N_C_M2_g N_C_c_28_n N_C_M6_g C VSS
+ PM_AND3X1_ASAP7_75T_R%C
x_PM_AND3X1_ASAP7_75T_R%6 N_6_M3_g N_6_c_52_n N_6_M7_g N_6_M0_s N_6_M4_s
+ N_6_c_38_n N_6_M6_s N_6_M5_d N_6_c_45_n N_6_c_61_p N_6_c_39_n N_6_c_40_n
+ N_6_c_69_p N_6_c_47_n N_6_c_70_p N_6_c_54_n N_6_c_42_n N_6_c_49_n N_6_c_56_n
+ N_6_c_67_p N_6_c_58_n N_6_c_64_p N_6_c_60_p N_6_c_68_p N_6_c_66_p VSS
+ PM_AND3X1_ASAP7_75T_R%6
x_PM_AND3X1_ASAP7_75T_R%Y N_Y_M3_d N_Y_M7_d N_Y_c_71_n N_Y_c_73_n N_Y_c_74_n Y
+ N_Y_c_76_n N_Y_c_77_n N_Y_c_79_n N_Y_c_80_n VSS PM_AND3X1_ASAP7_75T_R%Y
x_PM_AND3X1_ASAP7_75T_R%8 N_8_M1_s N_8_M0_d VSS PM_AND3X1_ASAP7_75T_R%8
x_PM_AND3X1_ASAP7_75T_R%9 N_9_M2_s N_9_M1_d VSS PM_AND3X1_ASAP7_75T_R%9
cc_1 N_A_M0_g N_B_M1_g 0.00327995f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_13_n 0.0011545f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A_c_3_p B 8.88497e-19 $X=0.081 $Y=0.135 $X2=0.138 $Y2=0.137
cc_4 A B 0.00130308f $X=0.019 $Y=0.137 $X2=0.138 $Y2=0.137
cc_5 N_A_M0_g N_C_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 A N_6_c_38_n 0.0014314f $X=0.019 $Y=0.137 $X2=0 $Y2=0
cc_7 A N_6_c_39_n 0.00142969f $X=0.019 $Y=0.137 $X2=0 $Y2=0
cc_8 N_A_M0_g N_6_c_40_n 4.30157e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_9 N_A_c_9_p N_6_c_40_n 9.97533e-19 $X=0.0605 $Y=0.135 $X2=0 $Y2=0
cc_10 N_A_M0_g N_6_c_42_n 4.30157e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_11 N_A_c_9_p N_6_c_42_n 9.97533e-19 $X=0.0605 $Y=0.135 $X2=0 $Y2=0
cc_12 N_B_M1_g N_C_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_13 N_B_c_13_n N_C_c_28_n 8.10277e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 B C 0.00586278f $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_15 N_B_M1_g N_6_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 B N_6_c_45_n 0.00114532f $X=0.138 $Y=0.137 $X2=0.018 $Y2=0.135
cc_17 B N_6_c_39_n 0.00106987f $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_18 N_B_M1_g N_6_c_47_n 3.39249e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 B N_6_c_47_n 0.00123619f $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_20 N_B_M1_g N_6_c_49_n 2.57255e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_21 B N_6_c_49_n 0.00123619f $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_22 N_C_M2_g N_6_M3_g 0.00284417f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_23 N_C_c_28_n N_6_c_52_n 9.81903e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_24 C N_6_c_45_n 0.00114532f $X=0.189 $Y=0.137 $X2=0.018 $Y2=0.135
cc_25 N_C_M2_g N_6_c_54_n 2.57255e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 C N_6_c_54_n 0.00123619f $X=0.189 $Y=0.137 $X2=0 $Y2=0
cc_27 N_C_M2_g N_6_c_56_n 2.64606e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_28 C N_6_c_56_n 0.00125368f $X=0.189 $Y=0.137 $X2=0 $Y2=0
cc_29 C N_6_c_58_n 0.0107712f $X=0.189 $Y=0.137 $X2=0 $Y2=0
cc_30 N_6_c_45_n N_Y_c_71_n 3.22701e-19 $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_31 N_6_c_60_p N_Y_c_71_n 0.0012561f $X=0.225 $Y=0.183 $X2=0 $Y2=0
cc_32 N_6_c_61_p N_Y_c_73_n 0.00170995f $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_33 N_6_c_61_p N_Y_c_74_n 0.00121787f $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_34 N_6_c_60_p Y 9.92725e-19 $X=0.225 $Y=0.183 $X2=0.081 $Y2=0.135
cc_35 N_6_c_64_p N_Y_c_76_n 8.57213e-19 $X=0.225 $Y=0.11 $X2=0.04 $Y2=0.135
cc_36 N_6_c_52_n N_Y_c_77_n 4.07842e-19 $X=0.243 $Y=0.135 $X2=0.0605 $Y2=0.135
cc_37 N_6_c_66_p N_Y_c_77_n 0.00105712f $X=0.248 $Y=0.135 $X2=0.0605 $Y2=0.135
cc_38 N_6_c_67_p N_Y_c_79_n 0.00170995f $X=0.225 $Y=0.07 $X2=0 $Y2=0
cc_39 N_6_c_68_p N_Y_c_80_n 0.00303709f $X=0.225 $Y=0.2 $X2=0 $Y2=0
cc_40 N_6_c_69_p N_8_M1_s 3.03001e-19 $X=0.126 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_41 N_6_c_70_p N_9_M2_s 3.56327e-19 $X=0.18 $Y=0.036 $X2=0.081 $Y2=0.0675

* END of "./AND3x1_ASAP7_75t_R.pex.sp.AND3X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: AND3x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:00:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AND3x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./AND3x2_ASAP7_75t_R.pex.sp.pex"
* File: AND3x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:00:11 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AND3X2_ASAP7_75T_R%A 2 5 7 18 21 24 VSS
c11 24 VSS 0.00875606f $X=0.019 $Y=0.137
c12 21 VSS 5.05467e-19 $X=0.0605 $Y=0.135
c13 20 VSS 0.00132257f $X=0.04 $Y=0.135
c14 18 VSS 6.00593e-19 $X=0.081 $Y=0.135
c15 5 VSS 0.00272543f $X=0.081 $Y=0.135
c16 2 VSS 0.0654968f $X=0.081 $Y=0.0675
r17 20 21 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.135 $X2=0.0605 $Y2=0.135
r18 18 21 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.0605 $Y2=0.135
r19 16 24 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r20 16 20 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.04 $Y2=0.135
r21 5 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AND3X2_ASAP7_75T_R%B 2 5 7 16 VSS
c16 16 VSS 0.00419374f $X=0.138 $Y=0.137
c17 5 VSS 9.94886e-19 $X=0.135 $Y=0.135
c18 2 VSS 0.0600755f $X=0.135 $Y=0.0675
r19 5 16 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r20 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r21 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AND3X2_ASAP7_75T_R%C 2 5 7 13 VSS
c13 13 VSS 0.00132189f $X=0.189 $Y=0.137
c14 5 VSS 9.808e-19 $X=0.189 $Y=0.135
c15 2 VSS 0.0583839f $X=0.189 $Y=0.0675
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AND3X2_ASAP7_75T_R%6 2 7 10 13 15 17 22 25 27 28 31 32 35 37 39 40 41
+ 51 53 56 60 61 62 65 66 68 71 74 77 VSS
c46 77 VSS 1.74783e-19 $X=0.225 $Y=0.135
c47 74 VSS 1.31878e-20 $X=0.2655 $Y=0.135
c48 73 VSS 7.16223e-19 $X=0.261 $Y=0.135
c49 71 VSS 1.63496e-19 $X=0.27 $Y=0.135
c50 68 VSS 1.87382e-19 $X=0.225 $Y=0.216
c51 67 VSS 2.19263e-19 $X=0.225 $Y=0.207
c52 66 VSS 3.97206e-19 $X=0.225 $Y=0.2
c53 65 VSS 0.00112931f $X=0.225 $Y=0.184
c54 64 VSS 1.76972e-19 $X=0.225 $Y=0.225
c55 62 VSS 4.69579e-19 $X=0.225 $Y=0.106
c56 61 VSS 3.85466e-19 $X=0.225 $Y=0.086
c57 60 VSS 2.34472e-19 $X=0.225 $Y=0.07
c58 59 VSS 3.64354e-19 $X=0.225 $Y=0.063
c59 58 VSS 7.16147e-19 $X=0.225 $Y=0.126
c60 56 VSS 0.00146362f $X=0.198 $Y=0.234
c61 55 VSS 0.00258369f $X=0.18 $Y=0.234
c62 54 VSS 8.80294e-19 $X=0.153 $Y=0.234
c63 53 VSS 0.00423484f $X=0.144 $Y=0.234
c64 52 VSS 0.00238018f $X=0.107 $Y=0.234
c65 51 VSS 0.00574452f $X=0.095 $Y=0.234
c66 43 VSS 0.00574187f $X=0.216 $Y=0.234
c67 42 VSS 0.00191122f $X=0.207 $Y=0.036
c68 41 VSS 0.00142296f $X=0.198 $Y=0.036
c69 40 VSS 0.00333444f $X=0.18 $Y=0.036
c70 39 VSS 0.00308768f $X=0.144 $Y=0.036
c71 38 VSS 0.0013368f $X=0.107 $Y=0.036
c72 37 VSS 0.00574452f $X=0.095 $Y=0.036
c73 35 VSS 0.00240442f $X=0.054 $Y=0.036
c74 32 VSS 0.00421964f $X=0.216 $Y=0.036
c75 31 VSS 0.0106914f $X=0.162 $Y=0.2025
c76 27 VSS 5.38922e-19 $X=0.179 $Y=0.2025
c77 25 VSS 0.00578446f $X=0.056 $Y=0.2025
c78 22 VSS 3.33606e-19 $X=0.071 $Y=0.2025
c79 17 VSS 3.33606e-19 $X=0.071 $Y=0.0675
c80 13 VSS 0.00462787f $X=0.297 $Y=0.135
c81 10 VSS 0.0639868f $X=0.297 $Y=0.0675
c82 2 VSS 0.0613357f $X=0.243 $Y=0.0675
r83 73 74 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.135 $X2=0.2655 $Y2=0.135
r84 71 74 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.135 $X2=0.2655 $Y2=0.135
r85 71 72 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.27 $Y=0.135 $X2=0.27
+ $Y2=0.135
r86 69 77 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.225 $Y2=0.135
r87 69 73 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.261 $Y2=0.135
r88 67 68 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.207 $X2=0.225 $Y2=0.216
r89 66 67 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.2 $X2=0.225 $Y2=0.207
r90 65 66 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.184 $X2=0.225 $Y2=0.2
r91 64 68 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.225 $X2=0.225 $Y2=0.216
r92 63 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.144 $X2=0.225 $Y2=0.135
r93 63 65 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.144 $X2=0.225 $Y2=0.184
r94 61 62 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.086 $X2=0.225 $Y2=0.106
r95 60 61 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.07 $X2=0.225 $Y2=0.086
r96 59 60 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.063 $X2=0.225 $Y2=0.07
r97 58 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r98 58 62 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.106
r99 57 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.063
r100 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r101 53 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.153 $Y2=0.234
r102 52 53 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.234 $X2=0.144 $Y2=0.234
r103 51 52 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.234 $X2=0.107 $Y2=0.234
r104 49 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r105 49 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.153 $Y2=0.234
r106 45 51 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.095 $Y2=0.234
r107 43 64 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.234 $X2=0.225 $Y2=0.225
r108 43 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.198 $Y2=0.234
r109 41 42 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.207 $Y2=0.036
r110 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r111 39 40 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.18 $Y2=0.036
r112 38 39 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.036 $X2=0.144 $Y2=0.036
r113 37 38 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.036 $X2=0.107 $Y2=0.036
r114 34 37 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.095 $Y2=0.036
r115 34 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r116 32 57 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.036 $X2=0.225 $Y2=0.045
r117 32 42 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.207 $Y2=0.036
r118 31 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r119 28 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r120 27 31 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r121 25 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r122 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r123 20 35 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.054 $Y=0.0675 $X2=0.054 $Y2=0.036
r124 17 20 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r125 13 72 27 $w=2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.297 $Y=0.135
+ $X2=0.27 $Y2=0.135
r126 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.135 $X2=0.297 $Y2=0.2025
r127 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.0675 $X2=0.297 $Y2=0.135
r128 5 72 27 $w=2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.243 $Y=0.135
+ $X2=0.27 $Y2=0.135
r129 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r130 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AND3X2_ASAP7_75T_R%Y 1 2 5 6 7 10 13 18 22 24 26 28 32 34 35 36 VSS
c21 38 VSS 0.00101302f $X=0.351 $Y=0.2045
c22 36 VSS 1.63987e-20 $X=0.351 $Y=0.14575
c23 35 VSS 7.60733e-19 $X=0.351 $Y=0.144
c24 34 VSS 0.00226498f $X=0.351 $Y=0.126
c25 33 VSS 0.00176873f $X=0.351 $Y=0.086
c26 32 VSS 0.00218466f $X=0.352 $Y=0.1475
c27 30 VSS 7.5805e-19 $X=0.351 $Y=0.225
c28 28 VSS 0.00318234f $X=0.313 $Y=0.234
c29 27 VSS 3.63468e-19 $X=0.284 $Y=0.234
c30 26 VSS 0.00201509f $X=0.279 $Y=0.234
c31 25 VSS 0.00755718f $X=0.342 $Y=0.234
c32 24 VSS 0.00318234f $X=0.313 $Y=0.036
c33 23 VSS 3.63468e-19 $X=0.284 $Y=0.036
c34 22 VSS 0.00201509f $X=0.279 $Y=0.036
c35 21 VSS 0.00755718f $X=0.342 $Y=0.036
c36 18 VSS 8.4555e-19 $X=0.27 $Y=0.198
c37 13 VSS 8.4555e-19 $X=0.27 $Y=0.072
c38 10 VSS 0.0110101f $X=0.27 $Y=0.2025
c39 6 VSS 5.81027e-19 $X=0.287 $Y=0.2025
c40 5 VSS 0.0108808f $X=0.27 $Y=0.0675
c41 1 VSS 5.81027e-19 $X=0.287 $Y=0.0675
r42 37 38 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.184 $X2=0.351 $Y2=0.2045
r43 35 36 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.144 $X2=0.351 $Y2=0.14575
r44 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.144
r45 33 34 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.086 $X2=0.351 $Y2=0.126
r46 32 37 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1475 $X2=0.351 $Y2=0.184
r47 32 36 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1475 $X2=0.351 $Y2=0.14575
r48 30 38 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.2045
r49 29 33 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.086
r50 27 28 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.234 $X2=0.313 $Y2=0.234
r51 26 27 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.234 $X2=0.284 $Y2=0.234
r52 25 30 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.234 $X2=0.351 $Y2=0.225
r53 25 28 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.313 $Y2=0.234
r54 23 24 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.036 $X2=0.313 $Y2=0.036
r55 22 23 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.036 $X2=0.284 $Y2=0.036
r56 21 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.036 $X2=0.351 $Y2=0.045
r57 21 24 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.313 $Y2=0.036
r58 16 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.27 $Y=0.225 $X2=0.279 $Y2=0.234
r59 16 18 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.225 $X2=0.27 $Y2=0.198
r60 11 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.27 $Y=0.045 $X2=0.279 $Y2=0.036
r61 11 13 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.045 $X2=0.27 $Y2=0.072
r62 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.198 $X2=0.27
+ $Y2=0.198
r63 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r64 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r65 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.072 $X2=0.27
+ $Y2=0.072
r66 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
r67 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends

.subckt PM_AND3X2_ASAP7_75T_R%8 1 2 VSS
c0 1 VSS 0.00241413f $X=0.125 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends

.subckt PM_AND3X2_ASAP7_75T_R%9 1 2 VSS
c1 1 VSS 0.00183233f $X=0.179 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.145 $Y2=0.0675
.ends


* END of "./AND3x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt AND3x2_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 N_8_M0_d N_A_M0_g N_6_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_9_M1_d N_B_M1_g N_8_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_C_M2_g N_9_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_6_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_6_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 VDD N_A_M5_g N_6_M5_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M6 N_6_M6_d N_B_M6_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M7 VDD N_C_M7_g N_6_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M8 N_Y_M8_d N_6_M8_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M9 N_Y_M9_d N_6_M9_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
*
* 
* .include "AND3x2_ASAP7_75t_R.pex.sp.AND3X2_ASAP7_75T_R.pxi"
* BEGIN of "./AND3x2_ASAP7_75t_R.pex.sp.AND3X2_ASAP7_75T_R.pxi"
* File: AND3x2_ASAP7_75t_R.pex.sp.AND3X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:00:11 2017
* 
x_PM_AND3X2_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M5_g N_A_c_3_p N_A_c_9_p A VSS
+ PM_AND3X2_ASAP7_75T_R%A
x_PM_AND3X2_ASAP7_75T_R%B N_B_M1_g N_B_c_13_n N_B_M6_g B VSS
+ PM_AND3X2_ASAP7_75T_R%B
x_PM_AND3X2_ASAP7_75T_R%C N_C_M2_g N_C_c_30_n N_C_M7_g C VSS
+ PM_AND3X2_ASAP7_75T_R%C
x_PM_AND3X2_ASAP7_75T_R%6 N_6_M3_g N_6_M8_g N_6_M4_g N_6_c_58_n N_6_M9_g
+ N_6_M0_s N_6_M5_s N_6_c_41_n N_6_M7_s N_6_M6_d N_6_c_48_n N_6_c_67_p
+ N_6_c_42_n N_6_c_43_n N_6_c_50_n N_6_c_86_p N_6_c_60_n N_6_c_45_n N_6_c_52_n
+ N_6_c_62_n N_6_c_54_n N_6_c_64_n N_6_c_83_p N_6_c_71_p N_6_c_76_p N_6_c_80_p
+ N_6_c_84_p N_6_c_74_p N_6_c_55_n VSS PM_AND3X2_ASAP7_75T_R%6
x_PM_AND3X2_ASAP7_75T_R%Y N_Y_M4_d N_Y_M3_d N_Y_c_88_n N_Y_M9_d N_Y_M8_d
+ N_Y_c_91_n N_Y_c_94_n N_Y_c_97_n N_Y_c_100_n N_Y_c_101_n N_Y_c_102_n
+ N_Y_c_103_n Y N_Y_c_104_n N_Y_c_106_n N_Y_c_107_n VSS PM_AND3X2_ASAP7_75T_R%Y
x_PM_AND3X2_ASAP7_75T_R%8 N_8_M1_s N_8_M0_d VSS PM_AND3X2_ASAP7_75T_R%8
x_PM_AND3X2_ASAP7_75T_R%9 N_9_M2_s N_9_M1_d VSS PM_AND3X2_ASAP7_75T_R%9
cc_1 N_A_M0_g N_B_M1_g 0.00327995f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_13_n 0.0011545f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A_c_3_p B 8.78098e-19 $X=0.081 $Y=0.135 $X2=0.138 $Y2=0.137
cc_4 A B 0.00129151f $X=0.019 $Y=0.137 $X2=0.138 $Y2=0.137
cc_5 N_A_M0_g N_C_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 A N_6_c_41_n 0.00138243f $X=0.019 $Y=0.137 $X2=0 $Y2=0
cc_7 A N_6_c_42_n 0.00138157f $X=0.019 $Y=0.137 $X2=0 $Y2=0
cc_8 N_A_M0_g N_6_c_43_n 4.30157e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_9 N_A_c_9_p N_6_c_43_n 9.97533e-19 $X=0.0605 $Y=0.135 $X2=0 $Y2=0
cc_10 N_A_M0_g N_6_c_45_n 4.30157e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_11 N_A_c_9_p N_6_c_45_n 9.97533e-19 $X=0.0605 $Y=0.135 $X2=0 $Y2=0
cc_12 N_B_M1_g N_C_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_13 N_B_c_13_n N_C_c_30_n 8.10277e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 B C 0.00567159f $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_15 N_B_M1_g N_6_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 B N_6_c_48_n 0.00137317f $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_17 B N_6_c_42_n 0.00141445f $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_18 N_B_M1_g N_6_c_50_n 3.23062e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 B N_6_c_50_n 0.0039815f $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_20 N_B_M1_g N_6_c_52_n 2.35211e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_21 B N_6_c_52_n 0.00375085f $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_22 B N_6_c_54_n 2.76275e-19 $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_23 B N_6_c_55_n 2.76275e-19 $X=0.138 $Y=0.137 $X2=0 $Y2=0
cc_24 N_C_M2_g N_6_M3_g 0.00284417f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_25 N_C_M2_g N_6_M4_g 2.31381e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 N_C_c_30_n N_6_c_58_n 9.55699e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_27 C N_6_c_48_n 0.00114532f $X=0.189 $Y=0.137 $X2=0 $Y2=0
cc_28 N_C_M2_g N_6_c_60_n 2.57255e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_29 C N_6_c_60_n 0.00123619f $X=0.189 $Y=0.137 $X2=0 $Y2=0
cc_30 N_C_M2_g N_6_c_62_n 2.64606e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_31 C N_6_c_62_n 0.00125368f $X=0.189 $Y=0.137 $X2=0 $Y2=0
cc_32 C N_6_c_64_n 0.010785f $X=0.189 $Y=0.137 $X2=0 $Y2=0
cc_33 N_6_c_58_n N_Y_M4_d 3.67694e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_34 N_6_c_58_n N_Y_c_88_n 5.03898e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_35 N_6_c_67_p N_Y_c_88_n 0.00134941f $X=0.216 $Y=0.036 $X2=0.081 $Y2=0.135
cc_36 N_6_c_58_n N_Y_M9_d 3.67694e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_37 N_6_c_58_n N_Y_c_91_n 5.03898e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_38 N_6_c_48_n N_Y_c_91_n 3.14194e-19 $X=0.162 $Y=0.2025 $X2=0 $Y2=0
cc_39 N_6_c_71_p N_Y_c_91_n 0.00134941f $X=0.225 $Y=0.184 $X2=0 $Y2=0
cc_40 N_6_c_58_n N_Y_c_94_n 2.02739e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_41 N_6_c_54_n N_Y_c_94_n 0.00177067f $X=0.225 $Y=0.07 $X2=0 $Y2=0
cc_42 N_6_c_74_p N_Y_c_94_n 4.88032e-19 $X=0.2655 $Y=0.135 $X2=0 $Y2=0
cc_43 N_6_c_58_n N_Y_c_97_n 2.02739e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_44 N_6_c_76_p N_Y_c_97_n 0.00177067f $X=0.225 $Y=0.2 $X2=0.081 $Y2=0.135
cc_45 N_6_c_74_p N_Y_c_97_n 4.88032e-19 $X=0.2655 $Y=0.135 $X2=0.081 $Y2=0.135
cc_46 N_6_c_67_p N_Y_c_100_n 0.00177067f $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_47 N_6_M4_g N_Y_c_101_n 2.91155e-19 $X=0.297 $Y=0.0675 $X2=0.019 $Y2=0.137
cc_48 N_6_c_80_p N_Y_c_102_n 0.00177067f $X=0.225 $Y=0.216 $X2=0 $Y2=0
cc_49 N_6_M4_g N_Y_c_103_n 2.91155e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_50 N_6_c_58_n N_Y_c_104_n 3.73466e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_51 N_6_c_83_p N_Y_c_104_n 4.12559e-19 $X=0.225 $Y=0.106 $X2=0 $Y2=0
cc_52 N_6_c_84_p N_Y_c_106_n 4.01628e-19 $X=0.27 $Y=0.135 $X2=0 $Y2=0
cc_53 N_6_c_71_p N_Y_c_107_n 4.09799e-19 $X=0.225 $Y=0.184 $X2=0 $Y2=0
cc_54 N_6_c_86_p N_9_M2_s 3.56327e-19 $X=0.18 $Y=0.036 $X2=0.081 $Y2=0.0675

* END of "./AND3x2_ASAP7_75t_R.pex.sp.AND3X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: AND3x4_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:00:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AND3x4_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./AND3x4_ASAP7_75t_R.pex.sp.pex"
* File: AND3x4_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:00:34 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AND3X4_ASAP7_75T_R%C 2 7 10 13 25 VSS
c10 25 VSS 0.0277251f $X=0.08 $Y=0.137
c11 13 VSS 0.00586133f $X=0.135 $Y=0.135
c12 10 VSS 0.0663694f $X=0.135 $Y=0.0675
c13 2 VSS 0.065408f $X=0.081 $Y=0.0675
r14 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r15 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081 $Y=0.135
+ $X2=0.135 $Y2=0.135
r16 5 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AND3X4_ASAP7_75T_R%B 2 7 10 13 23 VSS
c23 23 VSS 0.0103964f $X=0.296 $Y=0.137
c24 13 VSS 0.00667135f $X=0.351 $Y=0.135
c25 10 VSS 0.0640309f $X=0.351 $Y=0.0675
c26 2 VSS 0.0676956f $X=0.297 $Y=0.0675
r27 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r28 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297 $Y=0.135
+ $X2=0.351 $Y2=0.135
r29 5 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r30 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r31 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AND3X4_ASAP7_75T_R%A 2 8 11 13 22 VSS
c24 22 VSS 0.00438186f $X=0.458 $Y=0.137
c25 11 VSS 0.00361229f $X=0.459 $Y=0.135
c26 8 VSS 0.0650347f $X=0.459 $Y=0.0675
c27 2 VSS 0.063631f $X=0.405 $Y=0.0675
r28 11 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r29 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r30 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r31 5 11 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405 $Y=0.135
+ $X2=0.459 $Y2=0.135
r32 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AND3X4_ASAP7_75T_R%6 2 7 10 15 18 23 26 29 31 33 34 38 41 43 46 48 51
+ 53 55 63 64 68 69 70 71 72 74 77 79 82 84 85 86 89 90 96 VSS
c60 96 VSS 3.1582e-19 $X=0.567 $Y=0.135
c61 93 VSS 0.00196352f $X=0.604 $Y=0.135
c62 90 VSS 0.00134722f $X=0.567 $Y=0.207
c63 89 VSS 0.00283959f $X=0.567 $Y=0.189
c64 88 VSS 0.00109324f $X=0.567 $Y=0.225
c65 86 VSS 9.28104e-19 $X=0.567 $Y=0.117
c66 85 VSS 0.00104363f $X=0.567 $Y=0.099
c67 84 VSS 0.00118835f $X=0.567 $Y=0.081
c68 83 VSS 0.00109324f $X=0.567 $Y=0.063
c69 82 VSS 4.21868e-19 $X=0.567 $Y=0.126
c70 80 VSS 0.00376564f $X=0.529 $Y=0.036
c71 79 VSS 0.00689979f $X=0.5 $Y=0.036
c72 77 VSS 0.00331686f $X=0.432 $Y=0.036
c73 74 VSS 0.00676815f $X=0.558 $Y=0.036
c74 73 VSS 0.00376564f $X=0.529 $Y=0.234
c75 72 VSS 0.00298485f $X=0.5 $Y=0.234
c76 71 VSS 0.00429135f $X=0.487 $Y=0.234
c77 70 VSS 0.00705347f $X=0.45 $Y=0.234
c78 69 VSS 0.00861853f $X=0.3715 $Y=0.234
c79 68 VSS 0.0100259f $X=0.311 $Y=0.234
c80 64 VSS 0.00343051f $X=0.198 $Y=0.234
c81 63 VSS 0.00569711f $X=0.161 $Y=0.234
c82 55 VSS 0.00158099f $X=0.108 $Y=0.234
c83 53 VSS 0.00677413f $X=0.558 $Y=0.234
c84 51 VSS 0.00837437f $X=0.434 $Y=0.2025
c85 48 VSS 4.53693e-19 $X=0.449 $Y=0.2025
c86 46 VSS 0.00644867f $X=0.272 $Y=0.2025
c87 43 VSS 3.33606e-19 $X=0.287 $Y=0.2025
c88 41 VSS 0.00657477f $X=0.106 $Y=0.2025
c89 33 VSS 6.4978e-19 $X=0.449 $Y=0.0675
c90 29 VSS 0.017755f $X=0.783 $Y=0.135
c91 26 VSS 0.0645347f $X=0.783 $Y=0.0675
c92 18 VSS 0.0644226f $X=0.729 $Y=0.0675
c93 10 VSS 0.0644226f $X=0.675 $Y=0.0675
c94 2 VSS 0.0652433f $X=0.621 $Y=0.0675
r95 93 94 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.604 $Y=0.135 $X2=0.604
+ $Y2=0.135
r96 91 96 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.135 $X2=0.567 $Y2=0.135
r97 91 93 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.135 $X2=0.604 $Y2=0.135
r98 89 90 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.567 $Y2=0.207
r99 88 90 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.225 $X2=0.567 $Y2=0.207
r100 87 96 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.144 $X2=0.567 $Y2=0.135
r101 87 89 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.144 $X2=0.567 $Y2=0.189
r102 85 86 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.099 $X2=0.567 $Y2=0.117
r103 84 85 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.567 $Y2=0.099
r104 83 84 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.063 $X2=0.567 $Y2=0.081
r105 82 96 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.126 $X2=0.567 $Y2=0.135
r106 82 86 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.126 $X2=0.567 $Y2=0.117
r107 81 83 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.045 $X2=0.567 $Y2=0.063
r108 79 80 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5
+ $Y=0.036 $X2=0.529 $Y2=0.036
r109 76 79 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.5 $Y2=0.036
r110 76 77 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036
+ $X2=0.432 $Y2=0.036
r111 74 81 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.036 $X2=0.567 $Y2=0.045
r112 74 80 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.529 $Y2=0.036
r113 72 73 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.5
+ $Y=0.234 $X2=0.529 $Y2=0.234
r114 71 72 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.487
+ $Y=0.234 $X2=0.5 $Y2=0.234
r115 70 71 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.487 $Y2=0.234
r116 68 69 4.10802 $w=1.8e-08 $l=6.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.234 $X2=0.3715 $Y2=0.234
r117 66 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.45 $Y2=0.234
r118 66 69 4.10802 $w=1.8e-08 $l=6.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.3715 $Y2=0.234
r119 63 64 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.161
+ $Y=0.234 $X2=0.198 $Y2=0.234
r120 61 68 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.311 $Y2=0.234
r121 61 64 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.198 $Y2=0.234
r122 55 63 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.161 $Y2=0.234
r123 53 88 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.234 $X2=0.567 $Y2=0.225
r124 53 73 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.529 $Y2=0.234
r125 51 66 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r126 48 51 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.434 $Y2=0.2025
r127 46 61 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r128 43 46 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.272 $Y2=0.2025
r129 41 55 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r130 38 41 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.106 $Y2=0.2025
r131 37 77 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r132 34 37 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r133 33 37 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r134 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.135 $X2=0.783 $Y2=0.2025
r135 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.135
r136 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.135 $X2=0.783 $Y2=0.135
r137 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.135 $X2=0.729 $Y2=0.2025
r138 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.729 $Y=0.0675 $X2=0.729 $Y2=0.135
r139 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.675
+ $Y=0.135 $X2=0.729 $Y2=0.135
r140 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.135 $X2=0.675 $Y2=0.2025
r141 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.675 $Y=0.0675 $X2=0.675 $Y2=0.135
r142 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621
+ $Y=0.135 $X2=0.675 $Y2=0.135
r143 5 94 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.621
+ $Y=0.135 $X2=0.604 $Y2=0.135
r144 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r145 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
.ends

.subckt PM_AND3X4_ASAP7_75T_R%7 1 2 6 7 12 13 18 19 20 21 22 23 VSS
c21 23 VSS 0.00263599f $X=0.29 $Y=0.036
c22 22 VSS 0.00570028f $X=0.256 $Y=0.036
c23 21 VSS 0.00514322f $X=0.198 $Y=0.036
c24 20 VSS 0.00679243f $X=0.161 $Y=0.036
c25 19 VSS 0.00504846f $X=0.324 $Y=0.036
c26 18 VSS 0.00428455f $X=0.324 $Y=0.036
c27 13 VSS 0.00915316f $X=0.108 $Y=0.036
c28 12 VSS 0.00157935f $X=0.108 $Y=0.036
c29 6 VSS 6.06106e-19 $X=0.341 $Y=0.0675
c30 1 VSS 5.58795e-19 $X=0.125 $Y=0.0675
r31 22 23 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.036 $X2=0.29 $Y2=0.036
r32 21 22 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.256 $Y2=0.036
r33 20 21 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.161
+ $Y=0.036 $X2=0.198 $Y2=0.036
r34 18 23 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.29 $Y2=0.036
r35 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r36 12 20 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.161 $Y2=0.036
r37 12 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r38 10 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r39 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r40 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r41 5 13 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r42 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r43 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends

.subckt PM_AND3X4_ASAP7_75T_R%8 1 4 6 7 10 11 14 23 24 26 28 29 VSS
c31 29 VSS 2.77631e-19 $X=0.45 $Y=0.072
c32 28 VSS 0.00307218f $X=0.418 $Y=0.072
c33 26 VSS 5.9526e-19 $X=0.486 $Y=0.072
c34 24 VSS 1.76677e-19 $X=0.338 $Y=0.072
c35 23 VSS 4.26015e-19 $X=0.311 $Y=0.072
c36 14 VSS 0.00563836f $X=0.484 $Y=0.0675
c37 10 VSS 7.08605e-19 $X=0.378 $Y=0.0675
c38 6 VSS 6.69874e-19 $X=0.395 $Y=0.0675
c39 4 VSS 0.00440126f $X=0.272 $Y=0.0675
c40 1 VSS 3.2378e-19 $X=0.287 $Y=0.0675
r41 28 29 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.072 $X2=0.45 $Y2=0.072
r42 26 29 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.072 $X2=0.45 $Y2=0.072
r43 23 24 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.072 $X2=0.338 $Y2=0.072
r44 21 28 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.418 $Y2=0.072
r45 21 24 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.338 $Y2=0.072
r46 17 23 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.072 $X2=0.311 $Y2=0.072
r47 14 26 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.072 $X2=0.486
+ $Y2=0.072
r48 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.484 $Y2=0.0675
r49 10 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.072 $X2=0.378
+ $Y2=0.072
r50 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.378 $Y2=0.0675
r51 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.0675 $X2=0.378 $Y2=0.0675
r52 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.072 $X2=0.27
+ $Y2=0.072
r53 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.272 $Y2=0.0675
.ends

.subckt PM_AND3X4_ASAP7_75T_R%Y 1 2 6 7 11 12 15 16 17 20 21 24 28 29 40 41 VSS
c19 42 VSS 7.62145e-19 $X=0.837 $Y=0.144
c20 41 VSS 0.00529405f $X=0.837 $Y=0.126
c21 40 VSS 0.00529405f $X=0.8355 $Y=0.1465
c22 29 VSS 0.0265237f $X=0.828 $Y=0.234
c23 28 VSS 0.0092975f $X=0.756 $Y=0.036
c24 24 VSS 0.00913719f $X=0.648 $Y=0.036
c25 21 VSS 0.0265237f $X=0.828 $Y=0.036
c26 20 VSS 0.0092975f $X=0.756 $Y=0.2025
c27 16 VSS 5.38922e-19 $X=0.773 $Y=0.2025
c28 15 VSS 0.00930584f $X=0.648 $Y=0.2025
c29 11 VSS 5.72268e-19 $X=0.665 $Y=0.2025
c30 6 VSS 5.38922e-19 $X=0.773 $Y=0.0675
c31 1 VSS 5.72268e-19 $X=0.665 $Y=0.0675
r32 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.126 $X2=0.837 $Y2=0.144
r33 40 42 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.1465 $X2=0.837 $Y2=0.144
r34 38 40 5.33025 $w=1.8e-08 $l=7.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.1465
r35 37 41 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.045 $X2=0.837 $Y2=0.126
r36 31 35 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.756 $Y2=0.234
r37 29 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r38 29 35 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.756 $Y2=0.234
r39 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r40 23 27 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.756 $Y2=0.036
r41 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036 $X2=0.648
+ $Y2=0.036
r42 21 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.036 $X2=0.837 $Y2=0.045
r43 21 27 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.756 $Y2=0.036
r44 20 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234 $X2=0.756
+ $Y2=0.234
r45 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r46 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r47 15 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234 $X2=0.648
+ $Y2=0.234
r48 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.648 $Y2=0.2025
r49 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.648 $Y2=0.2025
r50 10 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.756
+ $Y=0.0675 $X2=0.756 $Y2=0.036
r51 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.756 $Y2=0.0675
r52 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.756 $Y2=0.0675
r53 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.648
+ $Y=0.0675 $X2=0.648 $Y2=0.036
r54 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.631
+ $Y=0.0675 $X2=0.648 $Y2=0.0675
r55 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.665
+ $Y=0.0675 $X2=0.648 $Y2=0.0675
.ends


* END of "./AND3x4_ASAP7_75t_R.pex.sp.pex"
* 
.subckt AND3x4_ASAP7_75t_R  VSS VDD C B A Y
* 
* Y	Y
* A	A
* B	B
* C	C
M0 N_7_M0_d N_C_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_7_M1_d N_C_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_7_M2_d N_B_M2_g N_8_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_7_M3_d N_B_M3_g N_8_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 N_6_M4_d N_A_M4_g N_8_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 N_6_M5_d N_A_M5_g N_8_M5_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 N_Y_M6_d N_6_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611 $Y=0.027
M7 N_Y_M7_d N_6_M7_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665 $Y=0.027
M8 N_Y_M8_d N_6_M8_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M9 N_Y_M9_d N_6_M9_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773 $Y=0.027
M10 N_6_M10_d N_C_M10_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M11 VDD N_B_M11_g N_6_M11_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M12 VDD N_A_M12_g N_6_M12_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M13 N_Y_M13_d N_6_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M14 N_Y_M14_d N_6_M14_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
M15 N_Y_M15_d N_6_M15_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M16 N_Y_M16_d N_6_M16_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
*
* 
* .include "AND3x4_ASAP7_75t_R.pex.sp.AND3X4_ASAP7_75T_R.pxi"
* BEGIN of "./AND3x4_ASAP7_75t_R.pex.sp.AND3X4_ASAP7_75T_R.pxi"
* File: AND3x4_ASAP7_75t_R.pex.sp.AND3X4_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:00:34 2017
* 
x_PM_AND3X4_ASAP7_75T_R%C N_C_M0_g N_C_M10_g N_C_M1_g N_C_c_2_p C VSS
+ PM_AND3X4_ASAP7_75T_R%C
x_PM_AND3X4_ASAP7_75T_R%B N_B_M2_g N_B_M11_g N_B_M3_g N_B_c_15_p B VSS
+ PM_AND3X4_ASAP7_75T_R%B
x_PM_AND3X4_ASAP7_75T_R%A N_A_M4_g N_A_M5_g N_A_c_37_n N_A_M12_g A VSS
+ PM_AND3X4_ASAP7_75T_R%A
x_PM_AND3X4_ASAP7_75T_R%6 N_6_M6_g N_6_M13_g N_6_M7_g N_6_M14_g N_6_M8_g
+ N_6_M15_g N_6_M9_g N_6_c_69_n N_6_M16_g N_6_M5_d N_6_M4_d N_6_M10_d N_6_c_58_n
+ N_6_M11_s N_6_c_63_n N_6_M12_s N_6_c_71_n N_6_c_116_p N_6_c_59_n N_6_c_61_n
+ N_6_c_64_n N_6_c_65_n N_6_c_68_n N_6_c_73_n N_6_c_75_n N_6_c_96_p N_6_c_109_p
+ N_6_c_77_n N_6_c_78_n N_6_c_79_n N_6_c_94_p N_6_c_91_p N_6_c_80_n N_6_c_81_n
+ N_6_c_82_n N_6_c_83_n VSS PM_AND3X4_ASAP7_75T_R%6
x_PM_AND3X4_ASAP7_75T_R%7 N_7_M1_d N_7_M0_d N_7_M3_d N_7_M2_d N_7_c_119_n
+ N_7_c_121_n N_7_c_124_n N_7_c_125_n N_7_c_122_n N_7_c_126_n N_7_c_127_n
+ N_7_c_128_n VSS PM_AND3X4_ASAP7_75T_R%7
x_PM_AND3X4_ASAP7_75T_R%8 N_8_M2_s N_8_c_139_n N_8_M4_s N_8_M3_s N_8_c_150_n
+ N_8_M5_s N_8_c_144_n N_8_c_140_n N_8_c_156_n N_8_c_145_n N_8_c_143_n
+ N_8_c_159_n VSS PM_AND3X4_ASAP7_75T_R%8
x_PM_AND3X4_ASAP7_75T_R%Y N_Y_M7_d N_Y_M6_d N_Y_M9_d N_Y_M8_d N_Y_M14_d
+ N_Y_M13_d N_Y_c_173_n N_Y_M16_d N_Y_M15_d N_Y_c_175_n N_Y_c_176_n N_Y_c_181_n
+ N_Y_c_182_n N_Y_c_183_n Y N_Y_c_188_n VSS PM_AND3X4_ASAP7_75T_R%Y
cc_1 C B 8.29454e-19 $X=0.08 $Y=0.137 $X2=0.296 $Y2=0.137
cc_2 N_C_c_2_p N_6_c_58_n 7.57503e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_3 N_C_c_2_p N_6_c_59_n 4.82735e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_4 C N_6_c_59_n 5.75458e-19 $X=0.08 $Y=0.137 $X2=0 $Y2=0
cc_5 N_C_M1_g N_6_c_61_n 4.61191e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_6 N_C_c_2_p N_7_M1_d 3.68024e-19 $X=0.135 $Y=0.135 $X2=0.297 $Y2=0.0675
cc_7 N_C_c_2_p N_7_c_119_n 5.15952e-19 $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.135
cc_8 C N_7_c_119_n 5.30913e-19 $X=0.08 $Y=0.137 $X2=0.351 $Y2=0.135
cc_9 N_C_c_2_p N_7_c_121_n 7.57503e-19 $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.135
cc_10 N_C_M1_g N_7_c_122_n 4.61191e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_11 N_B_M2_g N_A_M4_g 2.71887e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_12 N_B_M3_g N_A_M4_g 0.00364308f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_13 N_B_M3_g N_A_M5_g 3.00908e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_14 N_B_c_15_p N_A_c_37_n 0.00147059f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_15 B N_6_c_58_n 8.05623e-19 $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_16 B N_6_c_63_n 7.68375e-19 $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_17 B N_6_c_64_n 0.00373882f $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_18 N_B_M2_g N_6_c_65_n 4.30157e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_19 N_B_c_15_p N_6_c_65_n 8.41375e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_20 B N_6_c_65_n 0.00234629f $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_21 N_B_M3_g N_6_c_68_n 4.65034e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_22 N_B_c_15_p N_7_M3_d 3.67702e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_23 N_B_M2_g N_7_c_124_n 2.2196e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_24 N_B_c_15_p N_7_c_125_n 7.57503e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_25 B N_7_c_126_n 0.00376119f $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_26 B N_7_c_127_n 7.18834e-19 $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_27 B N_7_c_128_n 7.18834e-19 $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_28 B N_8_c_139_n 4.0584e-19 $X=0.296 $Y=0.137 $X2=0.081 $Y2=0.135
cc_29 N_B_M2_g N_8_c_140_n 3.33408e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_30 N_B_c_15_p N_8_c_140_n 0.00100715f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_31 B N_8_c_140_n 0.00255431f $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_32 N_B_M3_g N_8_c_143_n 4.96522e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_33 N_A_c_37_n N_6_c_69_n 2.45398e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_34 N_A_c_37_n N_6_M5_d 3.67193e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_35 N_A_c_37_n N_6_c_71_n 7.57503e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_36 A N_6_c_71_n 8.19478e-19 $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_37 N_A_M4_g N_6_c_73_n 4.65034e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_38 N_A_c_37_n N_6_c_73_n 4.9959e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_39 N_A_M5_g N_6_c_75_n 2.38524e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_40 A N_6_c_75_n 0.00376514f $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_41 N_A_c_37_n N_6_c_77_n 7.57503e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_42 N_A_M5_g N_6_c_78_n 2.38524e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_43 A N_6_c_79_n 3.26956e-19 $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_44 A N_6_c_80_n 4.27572e-19 $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_45 A N_6_c_81_n 3.26956e-19 $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_46 A N_6_c_82_n 3.45331e-19 $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_47 A N_6_c_83_n 3.26956e-19 $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_48 A N_8_c_144_n 9.62431e-19 $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_49 N_A_M5_g N_8_c_145_n 2.53669e-19 $X=0.459 $Y=0.0675 $X2=0.297 $Y2=0.135
cc_50 A N_8_c_145_n 0.00373988f $X=0.458 $Y=0.137 $X2=0.297 $Y2=0.135
cc_51 N_A_M4_g N_8_c_143_n 4.96522e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_52 N_A_c_37_n N_8_c_143_n 8.63627e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_53 N_6_c_58_n N_7_c_121_n 0.00105045f $X=0.106 $Y=0.2025 $X2=0.135 $Y2=0.135
cc_54 N_6_c_78_n N_7_c_124_n 3.04405e-19 $X=0.5 $Y=0.036 $X2=0 $Y2=0
cc_55 N_6_c_63_n N_8_c_139_n 0.00132173f $X=0.272 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_56 N_6_c_77_n N_8_c_150_n 0.0032943f $X=0.432 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_57 N_6_c_78_n N_8_c_150_n 4.51951e-19 $X=0.5 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_58 N_6_c_77_n N_8_c_144_n 0.00364651f $X=0.432 $Y=0.036 $X2=0 $Y2=0
cc_59 N_6_c_78_n N_8_c_144_n 0.00316793f $X=0.5 $Y=0.036 $X2=0 $Y2=0
cc_60 N_6_c_91_p N_8_c_144_n 3.59874e-19 $X=0.567 $Y=0.099 $X2=0 $Y2=0
cc_61 N_6_c_65_n N_8_c_140_n 2.65029e-19 $X=0.311 $Y=0.234 $X2=0 $Y2=0
cc_62 N_6_c_68_n N_8_c_156_n 2.65029e-19 $X=0.3715 $Y=0.234 $X2=0 $Y2=0
cc_63 N_6_c_94_p N_8_c_145_n 6.1248e-19 $X=0.567 $Y=0.081 $X2=0 $Y2=0
cc_64 N_6_c_73_n N_8_c_143_n 2.65029e-19 $X=0.45 $Y=0.234 $X2=0.081 $Y2=0.135
cc_65 N_6_c_96_p N_8_c_159_n 2.65029e-19 $X=0.5 $Y=0.234 $X2=0.081 $Y2=0.135
cc_66 N_6_c_77_n N_8_c_159_n 0.00233206f $X=0.432 $Y=0.036 $X2=0.081 $Y2=0.135
cc_67 N_6_c_78_n N_8_c_159_n 0.00679229f $X=0.5 $Y=0.036 $X2=0.081 $Y2=0.135
cc_68 N_6_c_69_n N_Y_M7_d 3.80663e-19 $X=0.783 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_69 N_6_c_69_n N_Y_M9_d 3.80663e-19 $X=0.783 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_70 N_6_c_69_n N_Y_M14_d 3.80663e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_71 N_6_c_69_n N_Y_c_173_n 8.00061e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_72 N_6_c_69_n N_Y_M16_d 3.80663e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_73 N_6_c_69_n N_Y_c_175_n 8.00061e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_74 N_6_M7_g N_Y_c_176_n 4.59284e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_75 N_6_M8_g N_Y_c_176_n 4.59284e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_76 N_6_M9_g N_Y_c_176_n 4.59284e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_77 N_6_c_69_n N_Y_c_176_n 0.00191346f $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_78 N_6_c_109_p N_Y_c_176_n 4.15041e-19 $X=0.558 $Y=0.036 $X2=0 $Y2=0
cc_79 N_6_c_69_n N_Y_c_181_n 8.00061e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_80 N_6_c_69_n N_Y_c_182_n 8.00061e-19 $X=0.783 $Y=0.135 $X2=0.081 $Y2=0.135
cc_81 N_6_M7_g N_Y_c_183_n 4.59284e-19 $X=0.675 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_82 N_6_M8_g N_Y_c_183_n 4.59284e-19 $X=0.729 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_83 N_6_M9_g N_Y_c_183_n 4.59284e-19 $X=0.783 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_84 N_6_c_69_n N_Y_c_183_n 0.00191346f $X=0.783 $Y=0.135 $X2=0.081 $Y2=0.135
cc_85 N_6_c_116_p N_Y_c_183_n 4.33639e-19 $X=0.558 $Y=0.234 $X2=0.081 $Y2=0.135
cc_86 N_6_c_69_n N_Y_c_188_n 5.76695e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_87 N_7_c_128_n N_8_M2_s 3.13602e-19 $X=0.29 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_88 N_7_c_125_n N_8_c_139_n 0.00350506f $X=0.324 $Y=0.036 $X2=0.081 $Y2=0.135
cc_89 N_7_c_128_n N_8_c_139_n 0.00279986f $X=0.29 $Y=0.036 $X2=0.081 $Y2=0.135
cc_90 N_7_c_124_n N_8_c_150_n 4.49606e-19 $X=0.324 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_91 N_7_c_125_n N_8_c_150_n 0.00318639f $X=0.324 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_92 N_7_c_128_n N_8_c_140_n 0.00352525f $X=0.29 $Y=0.036 $X2=0 $Y2=0
cc_93 N_7_c_124_n N_8_c_156_n 0.00352525f $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_94 N_7_c_125_n N_8_c_156_n 0.00233206f $X=0.324 $Y=0.036 $X2=0 $Y2=0

* END of "./AND3x4_ASAP7_75t_R.pex.sp.AND3X4_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: AND4x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:00:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AND4x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./AND4x1_ASAP7_75t_R.pex.sp.pex"
* File: AND4x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:00:56 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AND4X1_ASAP7_75T_R%A 2 5 7 13 VSS
c11 13 VSS 0.00188896f $X=0.081 $Y=0.138
c12 5 VSS 0.00222734f $X=0.081 $Y=0.135
c13 2 VSS 0.0640699f $X=0.081 $Y=0.0675
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AND4X1_ASAP7_75T_R%B 2 5 7 13 VSS
c10 13 VSS 0.00208027f $X=0.135 $Y=0.138
c11 5 VSS 0.00114876f $X=0.135 $Y=0.135
c12 2 VSS 0.0601793f $X=0.135 $Y=0.0675
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r14 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r15 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_AND4X1_ASAP7_75T_R%C 2 5 7 13 VSS
c12 13 VSS 0.00227424f $X=0.189 $Y=0.138
c13 5 VSS 0.00180716f $X=0.189 $Y=0.135
c14 2 VSS 0.0596433f $X=0.189 $Y=0.0675
r15 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_AND4X1_ASAP7_75T_R%D 2 5 7 15 VSS
c9 15 VSS 0.00169432f $X=0.243 $Y=0.138
c10 5 VSS 0.00112275f $X=0.243 $Y=0.135
c11 2 VSS 0.0600042f $X=0.243 $Y=0.0675
r12 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_AND4X1_ASAP7_75T_R%7 2 5 7 9 14 15 18 19 20 23 27 30 31 34 40 45 47
+ 50 51 54 VSS
c25 58 VSS 6.76599e-19 $X=0.297 $Y=0.1765
c26 54 VSS 5.90801e-19 $X=0.297 $Y=0.135
c27 52 VSS 4.85855e-19 $X=0.297 $Y=0.189
c28 51 VSS 1.80795e-19 $X=0.252 $Y=0.198
c29 50 VSS 0.00403754f $X=0.288 $Y=0.198
c30 49 VSS 8.72341e-19 $X=0.243 $Y=0.225
c31 47 VSS 0.00146362f $X=0.198 $Y=0.234
c32 46 VSS 0.00673385f $X=0.18 $Y=0.234
c33 45 VSS 0.00146362f $X=0.144 $Y=0.234
c34 44 VSS 0.00368081f $X=0.126 $Y=0.234
c35 40 VSS 0.00146362f $X=0.09 $Y=0.234
c36 39 VSS 0.0057813f $X=0.072 $Y=0.234
c37 35 VSS 0.00337635f $X=0.036 $Y=0.234
c38 34 VSS 0.0065785f $X=0.234 $Y=0.234
c39 31 VSS 0.0033144f $X=0.054 $Y=0.036
c40 30 VSS 0.005377f $X=0.054 $Y=0.036
c41 28 VSS 0.00330943f $X=0.036 $Y=0.036
c42 27 VSS 0.00580229f $X=0.027 $Y=0.2
c43 26 VSS 0.00112176f $X=0.027 $Y=0.07
c44 25 VSS 0.00110243f $X=0.027 $Y=0.225
c45 23 VSS 0.0104396f $X=0.216 $Y=0.2025
c46 19 VSS 6.1012e-19 $X=0.233 $Y=0.2025
c47 18 VSS 0.0104576f $X=0.108 $Y=0.2025
c48 14 VSS 6.1012e-19 $X=0.125 $Y=0.2025
c49 9 VSS 3.40659e-19 $X=0.071 $Y=0.0675
c50 5 VSS 0.00229683f $X=0.297 $Y=0.135
c51 2 VSS 0.0652694f $X=0.297 $Y=0.0675
r52 57 58 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.164 $X2=0.297 $Y2=0.1765
r53 54 57 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.164
r54 52 58 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.1765
r55 50 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.198 $X2=0.297 $Y2=0.189
r56 50 51 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.252 $Y2=0.198
r57 48 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.243 $Y=0.207 $X2=0.252 $Y2=0.198
r58 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.207 $X2=0.243 $Y2=0.225
r59 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r60 45 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.18 $Y2=0.234
r61 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r62 42 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.198 $Y2=0.234
r63 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r64 37 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r65 37 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.09 $Y2=0.234
r66 35 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.072 $Y2=0.234
r67 34 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.234 $X2=0.243 $Y2=0.225
r68 34 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.216 $Y2=0.234
r69 30 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r70 28 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.054 $Y2=0.036
r71 26 27 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.2
r72 25 35 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.225 $X2=0.036 $Y2=0.234
r73 25 27 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.2
r74 24 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r75 24 26 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r76 23 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234 $X2=0.216
+ $Y2=0.234
r77 20 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r78 19 23 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r79 18 37 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r80 15 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r81 14 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r82 12 31 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r83 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r84 5 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r85 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r86 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AND4X1_ASAP7_75T_R%Y 1 6 9 13 21 23 25 VSS
c7 31 VSS 0.00447704f $X=0.342 $Y=0.036
c8 30 VSS 0.00278493f $X=0.351 $Y=0.036
c9 28 VSS 0.00641345f $X=0.324 $Y=0.036
c10 25 VSS 0.00374407f $X=0.351 $Y=0.207
c11 23 VSS 9.47326e-19 $X=0.351 $Y=0.09225
c12 22 VSS 0.00126f $X=0.351 $Y=0.07
c13 21 VSS 0.00131406f $X=0.3515 $Y=0.1145
c14 19 VSS 7.23378e-19 $X=0.351 $Y=0.225
c15 13 VSS 0.00194221f $X=0.324 $Y=0.234
c16 11 VSS 0.00648807f $X=0.342 $Y=0.234
c17 9 VSS 0.00694916f $X=0.322 $Y=0.2025
c18 4 VSS 4.09605e-19 $X=0.322 $Y=0.0675
r19 31 32 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.3465 $Y2=0.036
r20 30 32 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.036 $X2=0.3465 $Y2=0.036
r21 27 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r22 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r23 24 25 5.90741 $w=1.8e-08 $l=8.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.12 $X2=0.351 $Y2=0.207
r24 22 23 1.5108 $w=1.8e-08 $l=2.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.07 $X2=0.351 $Y2=0.09225
r25 21 24 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1145 $X2=0.351 $Y2=0.12
r26 21 23 1.5108 $w=1.8e-08 $l=2.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1145 $X2=0.351 $Y2=0.09225
r27 19 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.207
r28 18 30 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.036
r29 18 22 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.07
r30 11 19 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.234 $X2=0.351 $Y2=0.225
r31 11 13 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.324 $Y2=0.234
r32 9 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r33 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2025 $X2=0.322 $Y2=0.2025
r34 4 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r35 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
.ends

.subckt PM_AND4X1_ASAP7_75T_R%9 1 2 VSS
c0 1 VSS 0.00228146f $X=0.125 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends

.subckt PM_AND4X1_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00228146f $X=0.179 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.145 $Y2=0.0675
.ends

.subckt PM_AND4X1_ASAP7_75T_R%11 1 2 VSS
c0 1 VSS 0.00228146f $X=0.233 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.199 $Y2=0.0675
.ends


* END of "./AND4x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt AND4x1_ASAP7_75t_R  VSS VDD A B C D Y
* 
* Y	Y
* D	D
* C	C
* B	B
* A	A
M0 N_9_M0_d N_A_M0_g N_7_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_10_M1_d N_B_M1_g N_9_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_11_M2_d N_C_M2_g N_10_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 VSS N_D_M3_g N_11_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_Y_M4_d N_7_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_7_M5_d N_A_M5_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M6 VDD N_B_M6_g N_7_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M7 N_7_M7_d N_C_M7_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M8 VDD N_D_M8_g N_7_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M9 N_Y_M9_d N_7_M9_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
*
* 
* .include "AND4x1_ASAP7_75t_R.pex.sp.AND4X1_ASAP7_75T_R.pxi"
* BEGIN of "./AND4x1_ASAP7_75t_R.pex.sp.AND4X1_ASAP7_75T_R.pxi"
* File: AND4x1_ASAP7_75t_R.pex.sp.AND4X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:00:56 2017
* 
x_PM_AND4X1_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M5_g A VSS
+ PM_AND4X1_ASAP7_75T_R%A
x_PM_AND4X1_ASAP7_75T_R%B N_B_M1_g N_B_c_13_n N_B_M6_g B VSS
+ PM_AND4X1_ASAP7_75T_R%B
x_PM_AND4X1_ASAP7_75T_R%C N_C_M2_g N_C_c_24_n N_C_M7_g C VSS
+ PM_AND4X1_ASAP7_75T_R%C
x_PM_AND4X1_ASAP7_75T_R%D N_D_M3_g N_D_c_36_n N_D_M8_g D VSS
+ PM_AND4X1_ASAP7_75T_R%D
x_PM_AND4X1_ASAP7_75T_R%7 N_7_M4_g N_7_c_59_n N_7_M9_g N_7_M0_s N_7_M6_s
+ N_7_M5_d N_7_c_43_n N_7_M8_s N_7_M7_d N_7_c_54_n N_7_c_44_n N_7_c_45_n
+ N_7_c_47_n N_7_c_65_p N_7_c_48_n N_7_c_51_n N_7_c_55_n N_7_c_66_p N_7_c_57_n
+ N_7_c_61_n VSS PM_AND4X1_ASAP7_75T_R%7
x_PM_AND4X1_ASAP7_75T_R%Y N_Y_M4_d N_Y_M9_d N_Y_c_69_n N_Y_c_71_n Y N_Y_c_68_n
+ N_Y_c_74_n VSS PM_AND4X1_ASAP7_75T_R%Y
x_PM_AND4X1_ASAP7_75T_R%9 N_9_M1_s N_9_M0_d VSS PM_AND4X1_ASAP7_75T_R%9
x_PM_AND4X1_ASAP7_75T_R%10 N_10_M2_s N_10_M1_d VSS PM_AND4X1_ASAP7_75T_R%10
x_PM_AND4X1_ASAP7_75T_R%11 N_11_M3_s N_11_M2_d VSS PM_AND4X1_ASAP7_75T_R%11
cc_1 N_A_M0_g N_B_M1_g 0.00357042f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_13_n 7.51046e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 A B 0.00588464f $X=0.081 $Y=0.138 $X2=0.135 $Y2=0.138
cc_4 N_A_M0_g N_C_M2_g 2.71887e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 A N_7_c_43_n 0.00114532f $X=0.081 $Y=0.138 $X2=0 $Y2=0
cc_6 A N_7_c_44_n 0.00500621f $X=0.081 $Y=0.138 $X2=0 $Y2=0
cc_7 N_A_M0_g N_7_c_45_n 9.16735e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_8 A N_7_c_45_n 9.05543e-19 $X=0.081 $Y=0.138 $X2=0 $Y2=0
cc_9 A N_7_c_47_n 0.0013295f $X=0.081 $Y=0.138 $X2=0 $Y2=0
cc_10 N_A_M0_g N_7_c_48_n 2.64924e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_11 A N_7_c_48_n 0.00125383f $X=0.081 $Y=0.138 $X2=0 $Y2=0
cc_12 N_B_M1_g N_C_M2_g 0.00327995f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_13 N_B_c_13_n N_C_c_24_n 7.51247e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 B C 0.00592435f $X=0.135 $Y=0.138 $X2=0.081 $Y2=0.138
cc_15 N_B_M1_g N_D_M3_g 2.66145e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 B N_7_c_43_n 0.00114532f $X=0.135 $Y=0.138 $X2=0 $Y2=0
cc_17 N_B_M1_g N_7_c_51_n 2.64606e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_18 B N_7_c_51_n 0.00125368f $X=0.135 $Y=0.138 $X2=0 $Y2=0
cc_19 N_C_M2_g N_D_M3_g 0.00343649f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_20 N_C_c_24_n N_D_c_36_n 7.51247e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 C D 0.0047228f $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_22 N_C_M2_g N_7_M4_g 2.31381e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_23 C N_7_c_54_n 0.00124979f $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_24 N_C_M2_g N_7_c_55_n 2.64924e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_25 C N_7_c_55_n 0.00125383f $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_26 C N_7_c_57_n 4.59663e-19 $X=0.189 $Y=0.138 $X2=0 $Y2=0
cc_27 N_D_M3_g N_7_M4_g 0.00287344f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_28 N_D_c_36_n N_7_c_59_n 7.73819e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_29 D N_7_c_57_n 0.00133641f $X=0.243 $Y=0.138 $X2=0 $Y2=0
cc_30 D N_7_c_61_n 0.00198065f $X=0.243 $Y=0.138 $X2=0 $Y2=0
cc_31 D N_Y_c_68_n 5.24405e-19 $X=0.243 $Y=0.138 $X2=0 $Y2=0
cc_32 N_7_c_54_n N_Y_c_69_n 2.81228e-19 $X=0.216 $Y=0.2025 $X2=0 $Y2=0
cc_33 N_7_c_61_n N_Y_c_69_n 0.00134786f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_34 N_7_M4_g N_Y_c_71_n 2.28931e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.138
cc_35 N_7_c_65_p N_Y_c_71_n 4.69503e-19 $X=0.234 $Y=0.234 $X2=0.081 $Y2=0.138
cc_36 N_7_c_66_p N_Y_c_71_n 6.32542e-19 $X=0.288 $Y=0.198 $X2=0.081 $Y2=0.138
cc_37 N_7_c_61_n N_Y_c_74_n 0.0035324f $X=0.297 $Y=0.135 $X2=0 $Y2=0

* END of "./AND4x1_ASAP7_75t_R.pex.sp.AND4X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: AND4x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:01:19 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AND4x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./AND4x2_ASAP7_75t_R.pex.sp.pex"
* File: AND4x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:01:19 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AND4X2_ASAP7_75T_R%A 2 7 10 13 21 VSS
c23 21 VSS 0.0197815f $X=0.061 $Y=0.1355
c24 13 VSS 0.00758098f $X=0.135 $Y=0.136
c25 10 VSS 0.0645939f $X=0.135 $Y=0.0675
c26 2 VSS 0.06799f $X=0.081 $Y=0.0675
r27 21 25 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.136 $X2=0.064
+ $Y2=0.136
r28 10 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.136
r29 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.136 $X2=0.135 $Y2=0.136
r30 5 25 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.136 $X2=0.064 $Y2=0.136
r31 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.136 $X2=0.081 $Y2=0.2025
r32 2 5 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.136
.ends

.subckt PM_AND4X2_ASAP7_75T_R%B 2 8 11 13 18 20 VSS
c27 20 VSS 0.00218956f $X=0.25 $Y=0.136
c28 18 VSS 0.00237675f $X=0.247 $Y=0.1195
c29 11 VSS 0.00800251f $X=0.243 $Y=0.136
c30 8 VSS 0.0681968f $X=0.243 $Y=0.0675
c31 2 VSS 0.0644017f $X=0.189 $Y=0.0675
r32 18 20 1.12037 $w=1.8e-08 $l=1.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.25
+ $Y=0.1195 $X2=0.25 $Y2=0.136
r33 11 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.25 $Y=0.136 $X2=0.25
+ $Y2=0.136
r34 11 13 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.136 $X2=0.243 $Y2=0.2025
r35 8 11 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.136
r36 5 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.136 $X2=0.243 $Y2=0.136
r37 2 5 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.136
.ends

.subckt PM_AND4X2_ASAP7_75T_R%C 2 7 10 13 20 23 25 VSS
c28 25 VSS 0.001827f $X=0.396 $Y=0.198
c29 20 VSS 0.00283532f $X=0.396 $Y=0.135
c30 13 VSS 0.00532398f $X=0.459 $Y=0.135
c31 10 VSS 0.0633454f $X=0.459 $Y=0.0675
c32 2 VSS 0.0674908f $X=0.405 $Y=0.0675
r33 23 25 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.393
+ $Y=0.198 $X2=0.396 $Y2=0.198
r34 18 25 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.189 $X2=0.396 $Y2=0.198
r35 18 20 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.189 $X2=0.396 $Y2=0.135
r36 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r37 5 13 57.2727 $w=2.2e-08 $l=6.3e-08 $layer=LIG $thickness=5e-08 $X=0.396
+ $Y=0.135 $X2=0.459 $Y2=0.135
r38 5 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.396 $Y=0.135 $X2=0.396
+ $Y2=0.135
r39 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r40 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AND4X2_ASAP7_75T_R%D 2 8 11 13 18 23 VSS
c26 23 VSS 0.00249815f $X=0.573 $Y=0.1525
c27 18 VSS 0.0128783f $X=0.576 $Y=0.134
c28 11 VSS 0.0110457f $X=0.567 $Y=0.134
c29 8 VSS 0.0678644f $X=0.567 $Y=0.0675
c30 2 VSS 0.0644557f $X=0.513 $Y=0.0675
r31 18 23 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.134 $X2=0.576 $Y2=0.1525
r32 11 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.576 $Y=0.134 $X2=0.576
+ $Y2=0.134
r33 11 13 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.134 $X2=0.567 $Y2=0.2025
r34 8 11 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.134
r35 5 11 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.134 $X2=0.567 $Y2=0.134
r36 2 5 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.134
.ends

.subckt PM_AND4X2_ASAP7_75T_R%7 2 7 10 13 15 17 18 21 22 25 27 30 32 35 37 40 44
+ 45 46 47 48 49 50 55 57 63 64 65 69 70 71 75 78 79 83 90 91 99 VSS
c68 99 VSS 0.00362026f $X=0.126 $Y=0.234
c69 91 VSS 2.62765e-19 $X=0.126 $Y=0.072
c70 90 VSS 1.70385e-19 $X=0.135 $Y=0.072
c71 83 VSS 0.00200635f $X=0.719 $Y=0.134
c72 80 VSS 0.00223614f $X=0.697 $Y=0.191
c73 79 VSS 0.00315862f $X=0.684 $Y=0.191
c74 78 VSS 5.38661e-19 $X=0.63 $Y=0.191
c75 77 VSS 0.00235454f $X=0.71 $Y=0.191
c76 76 VSS 2.6744e-19 $X=0.621 $Y=0.216
c77 75 VSS 1.98421e-19 $X=0.621 $Y=0.207
c78 74 VSS 2.52582e-19 $X=0.621 $Y=0.225
c79 72 VSS 4.75743e-19 $X=0.5895 $Y=0.234
c80 71 VSS 0.00465252f $X=0.585 $Y=0.234
c81 70 VSS 0.0108256f $X=0.541 $Y=0.234
c82 69 VSS 0.00151116f $X=0.446 $Y=0.234
c83 65 VSS 3.5855e-19 $X=0.43 $Y=0.234
c84 64 VSS 0.00384272f $X=0.428 $Y=0.234
c85 63 VSS 0.00719489f $X=0.387 $Y=0.234
c86 62 VSS 0.00953627f $X=0.345 $Y=0.234
c87 58 VSS 7.3748e-19 $X=0.2645 $Y=0.234
c88 57 VSS 0.00522587f $X=0.259 $Y=0.234
c89 56 VSS 0.00278169f $X=0.212 $Y=0.234
c90 55 VSS 0.00551485f $X=0.202 $Y=0.234
c91 51 VSS 0.00132597f $X=0.144 $Y=0.234
c92 50 VSS 0.00525392f $X=0.612 $Y=0.234
c93 49 VSS 4.00321e-19 $X=0.135 $Y=0.207
c94 48 VSS 6.09591e-19 $X=0.135 $Y=0.189
c95 46 VSS 3.15512e-19 $X=0.135 $Y=0.127
c96 45 VSS 2.18318e-19 $X=0.135 $Y=0.117
c97 44 VSS 8.2592e-20 $X=0.135 $Y=0.099
c98 43 VSS 9.3434e-19 $X=0.135 $Y=0.225
c99 40 VSS 0.00929132f $X=0.592 $Y=0.2025
c100 35 VSS 0.00887882f $X=0.43 $Y=0.2025
c101 30 VSS 0.00886505f $X=0.268 $Y=0.2025
c102 25 VSS 0.00865038f $X=0.106 $Y=0.2025
c103 21 VSS 0.00276064f $X=0.108 $Y=0.0675
c104 17 VSS 5.66579e-19 $X=0.125 $Y=0.0675
c105 13 VSS 0.00841531f $X=0.783 $Y=0.134
c106 10 VSS 0.0647445f $X=0.783 $Y=0.0675
c107 2 VSS 0.0654861f $X=0.729 $Y=0.0675
r108 99 100 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r109 98 100 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r110 95 99 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r111 91 92 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.1305 $Y2=0.072
r112 90 92 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.072 $X2=0.1305 $Y2=0.072
r113 87 91 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.072 $X2=0.126 $Y2=0.072
r114 83 84 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.719 $Y=0.134 $X2=0.719
+ $Y2=0.134
r115 81 83 3.25926 $w=1.8e-08 $l=4.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.719
+ $Y=0.182 $X2=0.719 $Y2=0.134
r116 79 80 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.684
+ $Y=0.191 $X2=0.697 $Y2=0.191
r117 78 79 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.191 $X2=0.684 $Y2=0.191
r118 77 81 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.71 $Y=0.191 $X2=0.719 $Y2=0.182
r119 77 80 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.71
+ $Y=0.191 $X2=0.697 $Y2=0.191
r120 75 76 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.207 $X2=0.621 $Y2=0.216
r121 74 76 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.216
r122 73 78 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.621 $Y=0.2 $X2=0.63 $Y2=0.191
r123 73 75 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.2 $X2=0.621 $Y2=0.207
r124 71 72 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.585
+ $Y=0.234 $X2=0.5895 $Y2=0.234
r125 70 71 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.541
+ $Y=0.234 $X2=0.585 $Y2=0.234
r126 69 70 6.45062 $w=1.8e-08 $l=9.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.446
+ $Y=0.234 $X2=0.541 $Y2=0.234
r127 67 72 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.5895 $Y2=0.234
r128 64 65 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.428
+ $Y=0.234 $X2=0.43 $Y2=0.234
r129 63 64 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.387
+ $Y=0.234 $X2=0.428 $Y2=0.234
r130 62 63 2.85185 $w=1.8e-08 $l=4.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.345
+ $Y=0.234 $X2=0.387 $Y2=0.234
r131 60 69 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.446 $Y2=0.234
r132 60 65 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.43 $Y2=0.234
r133 57 58 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.259
+ $Y=0.234 $X2=0.2645 $Y2=0.234
r134 56 57 3.19136 $w=1.8e-08 $l=4.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.212
+ $Y=0.234 $X2=0.259 $Y2=0.234
r135 55 56 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.234 $X2=0.212 $Y2=0.234
r136 53 62 5.09259 $w=1.8e-08 $l=7.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.345 $Y2=0.234
r137 53 58 0.373457 $w=1.8e-08 $l=5.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.2645 $Y2=0.234
r138 51 98 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.135 $Y2=0.234
r139 51 55 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.202 $Y2=0.234
r140 50 74 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r141 50 67 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.594 $Y2=0.234
r142 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.135 $Y2=0.207
r143 47 48 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.145 $X2=0.135 $Y2=0.189
r144 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.127 $X2=0.135 $Y2=0.145
r145 45 46 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.117 $X2=0.135 $Y2=0.127
r146 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.099 $X2=0.135 $Y2=0.117
r147 43 98 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.234
r148 43 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.207
r149 42 90 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.081 $X2=0.135 $Y2=0.072
r150 42 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.081 $X2=0.135 $Y2=0.099
r151 40 67 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r152 37 40 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2025 $X2=0.592 $Y2=0.2025
r153 35 60 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r154 32 35 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.43 $Y2=0.2025
r155 30 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r156 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.268 $Y2=0.2025
r157 25 95 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r158 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.106 $Y2=0.2025
r159 21 87 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.072
+ $X2=0.108 $Y2=0.072
r160 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r161 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r162 13 15 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.134 $X2=0.783 $Y2=0.2025
r163 10 13 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.783 $Y=0.0675 $X2=0.783 $Y2=0.134
r164 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.134 $X2=0.783 $Y2=0.134
r165 5 84 9.09091 $w=2.2e-08 $l=1e-08 $layer=LIG $thickness=5e-08 $X=0.729
+ $Y=0.134 $X2=0.719 $Y2=0.134
r166 5 7 256.635 $w=2e-08 $l=6.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.134 $X2=0.729 $Y2=0.2025
r167 2 5 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0675 $X2=0.729 $Y2=0.134
.ends

.subckt PM_AND4X2_ASAP7_75T_R%8 1 6 7 11 14 17 18 24 25 27 30 31 32 33 VSS
c27 33 VSS 0.00264484f $X=0.236 $Y=0.036
c28 32 VSS 0.00469161f $X=0.202 $Y=0.036
c29 31 VSS 0.00283808f $X=0.27 $Y=0.036
c30 30 VSS 0.00476776f $X=0.27 $Y=0.036
c31 28 VSS 9.52863e-19 $X=0.153 $Y=0.036
c32 27 VSS 0.00394048f $X=0.144 $Y=0.036
c33 26 VSS 0.00156718f $X=0.094 $Y=0.036
c34 25 VSS 0.00221358f $X=0.078 $Y=0.036
c35 24 VSS 0.00225071f $X=0.162 $Y=0.036
c36 18 VSS 0.00372502f $X=0.054 $Y=0.036
c37 17 VSS 0.00243247f $X=0.054 $Y=0.036
c38 14 VSS 5.8013e-19 $X=0.268 $Y=0.0675
c39 6 VSS 6.1381e-19 $X=0.179 $Y=0.0675
c40 1 VSS 4.56326e-19 $X=0.071 $Y=0.0675
r41 32 33 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.202
+ $Y=0.036 $X2=0.236 $Y2=0.036
r42 30 33 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.236 $Y2=0.036
r43 30 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r44 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.153 $Y2=0.036
r45 26 27 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.036 $X2=0.144 $Y2=0.036
r46 25 26 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.036 $X2=0.094 $Y2=0.036
r47 23 32 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.202 $Y2=0.036
r48 23 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.153 $Y2=0.036
r49 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r50 17 25 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.078 $Y2=0.036
r51 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r52 14 31 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r53 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.268 $Y2=0.0675
r54 10 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r55 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r56 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r57 4 18 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r58 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends

.subckt PM_AND4X2_ASAP7_75T_R%9 1 2 5 6 7 10 12 18 20 21 22 24 25 26 VSS
c29 27 VSS 2.05513e-19 $X=0.43 $Y=0.072
c30 26 VSS 4.90599e-19 $X=0.428 $Y=0.072
c31 25 VSS 3.72924e-19 $X=0.405 $Y=0.072
c32 24 VSS 0.00107587f $X=0.364 $Y=0.072
c33 23 VSS 0.00421258f $X=0.345 $Y=0.072
c34 22 VSS 4.97474e-19 $X=0.284 $Y=0.072
c35 21 VSS 5.73955e-20 $X=0.259 $Y=0.072
c36 20 VSS 3.15578e-20 $X=0.219 $Y=0.072
c37 18 VSS 2.48882e-19 $X=0.432 $Y=0.072
c38 12 VSS 3.17346e-19 $X=0.216 $Y=0.072
c39 10 VSS 0.0029383f $X=0.432 $Y=0.0675
c40 6 VSS 5.75221e-19 $X=0.449 $Y=0.0675
c41 5 VSS 0.00418138f $X=0.216 $Y=0.0675
c42 1 VSS 6.10138e-19 $X=0.233 $Y=0.0675
r43 26 27 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.428
+ $Y=0.072 $X2=0.43 $Y2=0.072
r44 25 26 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.072 $X2=0.428 $Y2=0.072
r45 24 25 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.364
+ $Y=0.072 $X2=0.405 $Y2=0.072
r46 23 24 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.345
+ $Y=0.072 $X2=0.364 $Y2=0.072
r47 22 23 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.072 $X2=0.345 $Y2=0.072
r48 21 22 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.259
+ $Y=0.072 $X2=0.284 $Y2=0.072
r49 20 21 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.219
+ $Y=0.072 $X2=0.259 $Y2=0.072
r50 18 27 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.072 $X2=0.43 $Y2=0.072
r51 12 20 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.072 $X2=0.219 $Y2=0.072
r52 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.072 $X2=0.432
+ $Y2=0.072
r53 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r54 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r55 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072 $X2=0.216
+ $Y2=0.072
r56 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r57 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends

.subckt PM_AND4X2_ASAP7_75T_R%10 1 6 7 11 14 18 22 23 24 26 27 28 29 VSS
c25 29 VSS 0.00365761f $X=0.567 $Y=0.036
c26 28 VSS 0.00817887f $X=0.541 $Y=0.036
c27 27 VSS 0.00837007f $X=0.594 $Y=0.036
c28 26 VSS 0.00433925f $X=0.594 $Y=0.036
c29 24 VSS 0.00175149f $X=0.466 $Y=0.036
c30 23 VSS 0.00726403f $X=0.446 $Y=0.036
c31 22 VSS 0.00551011f $X=0.486 $Y=0.036
c32 18 VSS 0.00348789f $X=0.378 $Y=0.036
c33 14 VSS 5.33282e-19 $X=0.592 $Y=0.0675
c34 6 VSS 5.38922e-19 $X=0.503 $Y=0.0675
c35 1 VSS 4.30437e-19 $X=0.395 $Y=0.0675
r36 28 29 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.541
+ $Y=0.036 $X2=0.567 $Y2=0.036
r37 26 29 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.567 $Y2=0.036
r38 26 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036 $X2=0.594
+ $Y2=0.036
r39 23 24 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.446
+ $Y=0.036 $X2=0.466 $Y2=0.036
r40 21 28 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.541 $Y2=0.036
r41 21 24 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.466 $Y2=0.036
r42 21 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036 $X2=0.486
+ $Y2=0.036
r43 17 23 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.446 $Y2=0.036
r44 17 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r45 14 27 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.594
+ $Y=0.0675 $X2=0.594 $Y2=0.036
r46 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0675 $X2=0.592 $Y2=0.0675
r47 10 22 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0675 $X2=0.486 $Y2=0.036
r48 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.486 $Y2=0.0675
r49 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.0675 $X2=0.486 $Y2=0.0675
r50 4 18 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r51 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.38 $Y2=0.0675
.ends

.subckt PM_AND4X2_ASAP7_75T_R%Y 1 2 6 7 10 11 14 16 24 27 VSS
c13 28 VSS 6.5344e-19 $X=0.837 $Y=0.2115
c14 27 VSS 0.00467692f $X=0.837 $Y=0.2
c15 26 VSS 0.00223165f $X=0.837 $Y=0.112
c16 25 VSS 0.00198469f $X=0.837 $Y=0.081
c17 24 VSS 6.57878e-19 $X=0.831 $Y=0.223
c18 16 VSS 0.0146565f $X=0.828 $Y=0.234
c19 14 VSS 0.00905362f $X=0.756 $Y=0.036
c20 11 VSS 0.0147042f $X=0.828 $Y=0.036
c21 10 VSS 0.00943367f $X=0.756 $Y=0.2025
c22 6 VSS 5.72268e-19 $X=0.773 $Y=0.2025
c23 1 VSS 5.72268e-19 $X=0.773 $Y=0.0675
r24 27 28 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.2 $X2=0.837 $Y2=0.2115
r25 26 27 5.97531 $w=1.8e-08 $l=8.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.112 $X2=0.837 $Y2=0.2
r26 25 26 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.081 $X2=0.837 $Y2=0.112
r27 24 28 0.780864 $w=1.8e-08 $l=1.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.223 $X2=0.837 $Y2=0.2115
r28 22 24 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.225 $X2=0.837 $Y2=0.223
r29 21 25 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.837
+ $Y=0.045 $X2=0.837 $Y2=0.081
r30 16 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.234 $X2=0.837 $Y2=0.225
r31 16 18 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.234 $X2=0.756 $Y2=0.234
r32 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036 $X2=0.756
+ $Y2=0.036
r33 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.828 $Y=0.036 $X2=0.837 $Y2=0.045
r34 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.828
+ $Y=0.036 $X2=0.756 $Y2=0.036
r35 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234 $X2=0.756
+ $Y2=0.234
r36 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.2025 $X2=0.756 $Y2=0.2025
r37 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.756 $Y2=0.2025
r38 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.756
+ $Y=0.0675 $X2=0.756 $Y2=0.036
r39 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.739
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
r40 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.773
+ $Y=0.0675 $X2=0.756 $Y2=0.0675
.ends


* END of "./AND4x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt AND4x2_ASAP7_75t_R  VSS VDD A B C D Y
* 
* Y	Y
* D	D
* C	C
* B	B
* A	A
M0 N_7_M0_d N_A_M0_g N_8_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_7_M1_d N_A_M1_g N_8_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_9_M2_d N_B_M2_g N_8_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_9_M3_d N_B_M3_g N_8_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_9_M4_d N_C_M4_g N_10_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 N_9_M5_d N_C_M5_g N_10_M5_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 VSS N_D_M6_g N_10_M6_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M7 VSS N_D_M7_g N_10_M7_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M8 N_Y_M8_d N_7_M8_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719 $Y=0.027
M9 N_Y_M9_d N_7_M9_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773 $Y=0.027
M10 N_7_M10_d N_A_M10_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M11 N_7_M11_d N_B_M11_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M12 N_7_M12_d N_C_M12_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M13 N_7_M13_d N_D_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M14 N_Y_M14_d N_7_M14_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.162
M15 N_Y_M15_d N_7_M15_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
*
* 
* .include "AND4x2_ASAP7_75t_R.pex.sp.AND4X2_ASAP7_75T_R.pxi"
* BEGIN of "./AND4x2_ASAP7_75t_R.pex.sp.AND4X2_ASAP7_75T_R.pxi"
* File: AND4x2_ASAP7_75t_R.pex.sp.AND4X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:01:19 2017
* 
x_PM_AND4X2_ASAP7_75T_R%A N_A_M0_g N_A_M10_g N_A_M1_g N_A_c_4_p A VSS
+ PM_AND4X2_ASAP7_75T_R%A
x_PM_AND4X2_ASAP7_75T_R%B N_B_M2_g N_B_M3_g N_B_c_27_n N_B_M11_g B N_B_c_30_p
+ VSS PM_AND4X2_ASAP7_75T_R%B
x_PM_AND4X2_ASAP7_75T_R%C N_C_M4_g N_C_M12_g N_C_M5_g N_C_c_51_n N_C_c_52_n C
+ N_C_c_53_n VSS PM_AND4X2_ASAP7_75T_R%C
x_PM_AND4X2_ASAP7_75T_R%D N_D_M6_g N_D_M7_g N_D_c_82_n N_D_M13_g N_D_c_83_n D
+ VSS PM_AND4X2_ASAP7_75T_R%D
x_PM_AND4X2_ASAP7_75T_R%7 N_7_M8_g N_7_M14_g N_7_M9_g N_7_c_137_n N_7_M15_g
+ N_7_M1_d N_7_M0_d N_7_c_106_n N_7_M10_d N_7_c_107_n N_7_M11_d N_7_c_119_n
+ N_7_M12_d N_7_c_129_n N_7_M13_d N_7_c_138_n N_7_c_108_n N_7_c_122_n
+ N_7_c_109_n N_7_c_110_n N_7_c_112_n N_7_c_124_n N_7_c_170_p N_7_c_125_n
+ N_7_c_127_n N_7_c_132_n N_7_c_133_n N_7_c_135_n N_7_c_158_p N_7_c_136_n
+ N_7_c_142_n N_7_c_144_n N_7_c_145_n N_7_c_147_n N_7_c_148_n N_7_c_152_p
+ N_7_c_115_n N_7_c_117_n VSS PM_AND4X2_ASAP7_75T_R%7
x_PM_AND4X2_ASAP7_75T_R%8 N_8_M0_s N_8_M2_s N_8_M1_s N_8_M3_s N_8_c_196_p
+ N_8_c_174_n N_8_c_175_n N_8_c_184_n N_8_c_176_n N_8_c_177_n N_8_c_178_n
+ N_8_c_179_n N_8_c_180_n N_8_c_191_p VSS PM_AND4X2_ASAP7_75T_R%8
x_PM_AND4X2_ASAP7_75T_R%9 N_9_M3_d N_9_M2_d N_9_c_201_n N_9_M5_d N_9_M4_d
+ N_9_c_207_n N_9_c_203_n N_9_c_226_p N_9_c_218_n N_9_c_204_n N_9_c_220_n
+ N_9_c_209_n N_9_c_222_p N_9_c_210_n VSS PM_AND4X2_ASAP7_75T_R%9
x_PM_AND4X2_ASAP7_75T_R%10 N_10_M4_s N_10_M6_s N_10_M5_s N_10_M7_s N_10_c_235_n
+ N_10_c_230_n N_10_c_250_n N_10_c_232_n N_10_c_233_n N_10_c_236_n N_10_c_237_n
+ N_10_c_239_n N_10_c_241_n VSS PM_AND4X2_ASAP7_75T_R%10
x_PM_AND4X2_ASAP7_75T_R%Y N_Y_M9_d N_Y_M8_d N_Y_M15_d N_Y_M14_d N_Y_c_257_n
+ N_Y_c_254_n N_Y_c_261_n N_Y_c_262_n Y N_Y_c_265_n VSS PM_AND4X2_ASAP7_75T_R%Y
cc_1 N_A_M0_g N_B_M2_g 3.03912e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_A_M1_g N_B_M2_g 0.0036697f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A_M1_g N_B_M3_g 2.74891e-19 $X=0.135 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_4 N_A_c_4_p N_B_c_27_n 0.00138172f $X=0.135 $Y=0.136 $X2=0.243 $Y2=0.136
cc_5 N_A_c_4_p N_7_M1_d 3.74131e-19 $X=0.135 $Y=0.136 $X2=0.25 $Y2=0.1195
cc_6 N_A_c_4_p N_7_c_106_n 7.60428e-19 $X=0.135 $Y=0.136 $X2=0.25 $Y2=0.136
cc_7 N_A_c_4_p N_7_c_107_n 8.43851e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_8 A N_7_c_108_n 4.8654e-19 $X=0.061 $Y=0.1355 $X2=0 $Y2=0
cc_9 N_A_c_4_p N_7_c_109_n 4.8859e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_10 N_A_c_4_p N_7_c_110_n 0.00136752f $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_11 A N_7_c_110_n 5.23274e-19 $X=0.061 $Y=0.1355 $X2=0 $Y2=0
cc_12 N_A_M1_g N_7_c_112_n 4.86515e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_13 N_A_c_4_p N_7_c_112_n 4.97174e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_14 A N_7_c_112_n 6.74927e-19 $X=0.061 $Y=0.1355 $X2=0 $Y2=0
cc_15 N_A_c_4_p N_7_c_115_n 4.99795e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_16 A N_7_c_115_n 6.07916e-19 $X=0.061 $Y=0.1355 $X2=0 $Y2=0
cc_17 N_A_c_4_p N_7_c_117_n 2.85448e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_18 A N_7_c_117_n 7.22154e-19 $X=0.061 $Y=0.1355 $X2=0 $Y2=0
cc_19 A N_8_M0_s 2.23359e-19 $X=0.061 $Y=0.1355 $X2=0.189 $Y2=0.0675
cc_20 A N_8_c_174_n 0.00147537f $X=0.061 $Y=0.1355 $X2=0.25 $Y2=0.1195
cc_21 A N_8_c_175_n 0.00233258f $X=0.061 $Y=0.1355 $X2=0.247 $Y2=0.1195
cc_22 N_A_c_4_p N_8_c_176_n 3.35575e-19 $X=0.135 $Y=0.136 $X2=0 $Y2=0
cc_23 N_A_M1_g N_8_c_177_n 2.35211e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_24 N_B_c_27_n N_C_c_51_n 4.40768e-19 $X=0.243 $Y=0.136 $X2=0.135 $Y2=0.136
cc_25 B N_C_c_52_n 8.37738e-19 $X=0.247 $Y=0.1195 $X2=0 $Y2=0
cc_26 N_B_c_30_p N_C_c_53_n 4.08302e-19 $X=0.25 $Y=0.136 $X2=0.064 $Y2=0.136
cc_27 N_B_c_27_n N_7_c_119_n 2.10963e-19 $X=0.243 $Y=0.136 $X2=0 $Y2=0
cc_28 B N_7_c_119_n 4.18098e-19 $X=0.247 $Y=0.1195 $X2=0 $Y2=0
cc_29 N_B_c_30_p N_7_c_119_n 8.95126e-19 $X=0.25 $Y=0.136 $X2=0 $Y2=0
cc_30 B N_7_c_122_n 3.38877e-19 $X=0.247 $Y=0.1195 $X2=0 $Y2=0
cc_31 B N_7_c_109_n 8.78989e-19 $X=0.247 $Y=0.1195 $X2=0 $Y2=0
cc_32 N_B_c_30_p N_7_c_124_n 3.68337e-19 $X=0.25 $Y=0.136 $X2=0 $Y2=0
cc_33 N_B_M2_g N_7_c_125_n 4.56095e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_34 N_B_c_27_n N_7_c_125_n 4.01894e-19 $X=0.243 $Y=0.136 $X2=0 $Y2=0
cc_35 N_B_M3_g N_7_c_127_n 2.64526e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B_c_30_p N_7_c_127_n 0.00452342f $X=0.25 $Y=0.136 $X2=0 $Y2=0
cc_37 N_B_M3_g N_8_c_178_n 2.2196e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_38 B N_8_c_179_n 4.21932e-19 $X=0.247 $Y=0.1195 $X2=0 $Y2=0
cc_39 N_B_M2_g N_8_c_180_n 4.61191e-19 $X=0.189 $Y=0.0675 $X2=0.064 $Y2=0.136
cc_40 N_B_c_27_n N_8_c_180_n 2.65146e-19 $X=0.243 $Y=0.136 $X2=0.064 $Y2=0.136
cc_41 N_B_c_27_n N_9_M3_d 3.70805e-19 $X=0.243 $Y=0.136 $X2=0.081 $Y2=0.0675
cc_42 N_B_c_27_n N_9_c_201_n 7.60428e-19 $X=0.243 $Y=0.136 $X2=0.081 $Y2=0.136
cc_43 B N_9_c_201_n 8.87973e-19 $X=0.247 $Y=0.1195 $X2=0.081 $Y2=0.136
cc_44 N_B_c_27_n N_9_c_203_n 2.30331e-19 $X=0.243 $Y=0.136 $X2=0.135 $Y2=0.136
cc_45 N_B_M3_g N_9_c_204_n 2.85825e-19 $X=0.243 $Y=0.0675 $X2=0.061 $Y2=0.1355
cc_46 B N_9_c_204_n 0.00398489f $X=0.247 $Y=0.1195 $X2=0.061 $Y2=0.1355
cc_47 N_C_M4_g N_D_M6_g 2.98169e-19 $X=0.405 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_48 N_C_M5_g N_D_M6_g 0.00354623f $X=0.459 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_49 N_C_M5_g N_D_M7_g 2.34385e-19 $X=0.459 $Y=0.0675 $X2=0.243 $Y2=0.0675
cc_50 N_C_c_51_n N_D_c_82_n 0.00161002f $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.136
cc_51 N_C_c_52_n N_D_c_83_n 2.49014e-19 $X=0.396 $Y=0.135 $X2=0.247 $Y2=0.1195
cc_52 N_C_c_52_n D 2.49014e-19 $X=0.396 $Y=0.135 $X2=0 $Y2=0
cc_53 N_C_c_51_n N_7_c_129_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_54 N_C_c_52_n N_7_c_129_n 8.41502e-19 $X=0.396 $Y=0.135 $X2=0 $Y2=0
cc_55 N_C_c_53_n N_7_c_129_n 0.00135469f $X=0.396 $Y=0.198 $X2=0 $Y2=0
cc_56 N_C_c_52_n N_7_c_132_n 6.38598e-19 $X=0.396 $Y=0.135 $X2=0 $Y2=0
cc_57 N_C_M4_g N_7_c_133_n 2.64781e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_C_c_53_n N_7_c_133_n 0.00403472f $X=0.396 $Y=0.198 $X2=0 $Y2=0
cc_59 N_C_c_51_n N_7_c_135_n 3.80706e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_60 N_C_M5_g N_7_c_136_n 4.58656e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_61 N_C_c_51_n N_9_M5_d 3.80371e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_62 N_C_c_51_n N_9_c_207_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.243 $Y2=0.136
cc_63 N_C_c_52_n N_9_c_207_n 2.91667e-19 $X=0.396 $Y=0.135 $X2=0.243 $Y2=0.136
cc_64 N_C_c_52_n N_9_c_209_n 0.00557875f $X=0.396 $Y=0.135 $X2=0 $Y2=0
cc_65 N_C_c_51_n N_9_c_210_n 5.89092e-19 $X=0.459 $Y=0.135 $X2=0.189 $Y2=0.136
cc_66 N_C_c_52_n N_10_M4_s 2.04552e-19 $X=0.396 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_67 N_C_c_51_n N_10_c_230_n 2.00015e-19 $X=0.459 $Y=0.135 $X2=0.247 $Y2=0.1195
cc_68 N_C_c_52_n N_10_c_230_n 0.00135993f $X=0.396 $Y=0.135 $X2=0.247 $Y2=0.1195
cc_69 N_C_M4_g N_10_c_232_n 2.64781e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_70 N_C_M5_g N_10_c_233_n 3.89858e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_71 N_C_c_51_n N_10_c_233_n 2.53248e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_72 N_D_c_82_n N_7_c_137_n 4.64422e-19 $X=0.567 $Y=0.134 $X2=0.459 $Y2=0.135
cc_73 N_D_c_83_n N_7_c_138_n 4.53921e-19 $X=0.576 $Y=0.134 $X2=0 $Y2=0
cc_74 D N_7_c_138_n 8.44726e-19 $X=0.573 $Y=0.1525 $X2=0 $Y2=0
cc_75 N_D_M6_g N_7_c_136_n 4.61191e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_76 N_D_c_82_n N_7_c_136_n 4.89004e-19 $X=0.567 $Y=0.134 $X2=0 $Y2=0
cc_77 N_D_M7_g N_7_c_142_n 2.65027e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_78 D N_7_c_142_n 0.00428211f $X=0.573 $Y=0.1525 $X2=0 $Y2=0
cc_79 D N_7_c_144_n 6.41437e-19 $X=0.573 $Y=0.1525 $X2=0 $Y2=0
cc_80 N_D_c_83_n N_7_c_145_n 6.86517e-19 $X=0.576 $Y=0.134 $X2=0 $Y2=0
cc_81 D N_7_c_145_n 6.41437e-19 $X=0.573 $Y=0.1525 $X2=0 $Y2=0
cc_82 N_D_c_83_n N_7_c_147_n 6.86517e-19 $X=0.576 $Y=0.134 $X2=0 $Y2=0
cc_83 N_D_c_83_n N_7_c_148_n 7.38337e-19 $X=0.576 $Y=0.134 $X2=0 $Y2=0
cc_84 N_D_c_83_n N_10_c_235_n 2.87556e-19 $X=0.576 $Y=0.134 $X2=0 $Y2=0
cc_85 N_D_c_83_n N_10_c_236_n 0.00398859f $X=0.576 $Y=0.134 $X2=0 $Y2=0
cc_86 N_D_c_82_n N_10_c_237_n 2.10963e-19 $X=0.567 $Y=0.134 $X2=0 $Y2=0
cc_87 N_D_c_83_n N_10_c_237_n 0.00342538f $X=0.576 $Y=0.134 $X2=0 $Y2=0
cc_88 N_D_M6_g N_10_c_239_n 4.56095e-19 $X=0.513 $Y=0.0675 $X2=0.396 $Y2=0.135
cc_89 N_D_c_82_n N_10_c_239_n 8.90257e-19 $X=0.567 $Y=0.134 $X2=0.396 $Y2=0.135
cc_90 N_D_M7_g N_10_c_241_n 2.30186e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_91 N_D_c_83_n N_Y_c_254_n 2.66253e-19 $X=0.576 $Y=0.134 $X2=0 $Y2=0
cc_92 N_7_c_106_n N_8_c_175_n 0.0037765f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_93 N_7_c_115_n N_8_c_175_n 3.32544e-19 $X=0.126 $Y=0.072 $X2=0 $Y2=0
cc_94 N_7_c_106_n N_8_c_184_n 0.00311019f $X=0.108 $Y=0.0675 $X2=0.064 $Y2=0.136
cc_95 N_7_c_152_p N_8_c_184_n 0.00125338f $X=0.135 $Y=0.072 $X2=0.064 $Y2=0.136
cc_96 N_7_c_106_n N_8_c_177_n 0.00250914f $X=0.108 $Y=0.0675 $X2=0 $Y2=0
cc_97 N_7_c_115_n N_8_c_177_n 0.00470294f $X=0.126 $Y=0.072 $X2=0 $Y2=0
cc_98 N_7_c_119_n N_8_c_179_n 0.00136032f $X=0.268 $Y=0.2025 $X2=0 $Y2=0
cc_99 N_7_c_129_n N_9_c_207_n 0.00148182f $X=0.43 $Y=0.2025 $X2=0.135 $Y2=0.0675
cc_100 N_7_c_152_p N_9_c_203_n 3.80515e-19 $X=0.135 $Y=0.072 $X2=0.135 $Y2=0.136
cc_101 N_7_c_158_p N_10_c_233_n 3.04329e-19 $X=0.446 $Y=0.234 $X2=0.064
+ $Y2=0.136
cc_102 N_7_c_138_n N_10_c_237_n 0.00132309f $X=0.592 $Y=0.2025 $X2=0 $Y2=0
cc_103 N_7_c_136_n N_10_c_239_n 3.04329e-19 $X=0.541 $Y=0.234 $X2=0 $Y2=0
cc_104 N_7_c_137_n N_Y_M9_d 3.87022e-19 $X=0.783 $Y=0.134 $X2=0.081 $Y2=0.0675
cc_105 N_7_c_137_n N_Y_M15_d 3.7444e-19 $X=0.783 $Y=0.134 $X2=0.081 $Y2=0.2025
cc_106 N_7_c_137_n N_Y_c_257_n 7.60428e-19 $X=0.783 $Y=0.134 $X2=0.135
+ $Y2=0.0675
cc_107 N_7_c_148_n N_Y_c_257_n 0.00115663f $X=0.719 $Y=0.134 $X2=0.135
+ $Y2=0.0675
cc_108 N_7_M9_g N_Y_c_254_n 4.56718e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_109 N_7_c_137_n N_Y_c_254_n 6.56931e-19 $X=0.783 $Y=0.134 $X2=0 $Y2=0
cc_110 N_7_c_137_n N_Y_c_261_n 8.43851e-19 $X=0.783 $Y=0.134 $X2=0 $Y2=0
cc_111 N_7_M9_g N_Y_c_262_n 4.61823e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_112 N_7_c_137_n N_Y_c_262_n 6.44171e-19 $X=0.783 $Y=0.134 $X2=0 $Y2=0
cc_113 N_7_c_170_p N_Y_c_262_n 2.06604e-19 $X=0.612 $Y=0.234 $X2=0 $Y2=0
cc_114 N_7_c_137_n N_Y_c_265_n 4.78361e-19 $X=0.783 $Y=0.134 $X2=0 $Y2=0
cc_115 N_7_c_148_n N_Y_c_265_n 0.00101786f $X=0.719 $Y=0.134 $X2=0 $Y2=0
cc_116 N_8_c_184_n N_9_c_201_n 0.00378484f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.136
cc_117 N_8_c_179_n N_9_c_201_n 0.00391031f $X=0.27 $Y=0.036 $X2=0.081 $Y2=0.136
cc_118 N_8_c_191_p N_9_c_201_n 0.00258679f $X=0.236 $Y=0.036 $X2=0.081 $Y2=0.136
cc_119 N_8_c_184_n N_9_c_203_n 3.9589e-19 $X=0.162 $Y=0.036 $X2=0.135 $Y2=0.136
cc_120 N_8_c_191_p N_9_c_203_n 0.003517f $X=0.236 $Y=0.036 $X2=0.135 $Y2=0.136
cc_121 N_8_c_178_n N_9_c_218_n 0.003517f $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_122 N_8_c_179_n N_9_c_204_n 4.19603e-19 $X=0.27 $Y=0.036 $X2=0.061 $Y2=0.1355
cc_123 N_8_c_196_p N_9_c_220_n 2.87556e-19 $X=0.268 $Y=0.0675 $X2=0 $Y2=0
cc_124 N_8_c_179_n N_9_c_220_n 0.00215527f $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_125 N_8_c_179_n N_10_c_230_n 0.00136914f $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_126 N_8_c_178_n N_10_c_232_n 6.78329e-19 $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_127 N_9_c_222_p N_10_M4_s 3.3673e-19 $X=0.405 $Y=0.072 $X2=0.189 $Y2=0.0675
cc_128 N_9_c_207_n N_10_c_230_n 0.00372805f $X=0.432 $Y=0.0675 $X2=0.247
+ $Y2=0.1195
cc_129 N_9_c_222_p N_10_c_230_n 0.00268579f $X=0.405 $Y=0.072 $X2=0.247
+ $Y2=0.1195
cc_130 N_9_c_207_n N_10_c_250_n 0.0032866f $X=0.432 $Y=0.0675 $X2=0 $Y2=0
cc_131 N_9_c_226_p N_10_c_250_n 5.01471e-19 $X=0.432 $Y=0.072 $X2=0 $Y2=0
cc_132 N_9_c_207_n N_10_c_232_n 0.00254576f $X=0.432 $Y=0.0675 $X2=0 $Y2=0
cc_133 N_9_c_222_p N_10_c_232_n 0.00705753f $X=0.405 $Y=0.072 $X2=0 $Y2=0

* END of "./AND4x2_ASAP7_75t_R.pex.sp.AND4X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: AND5x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:01:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AND5x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./AND5x1_ASAP7_75t_R.pex.sp.pex"
* File: AND5x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:01:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AND5X1_ASAP7_75T_R%A 2 5 7 13 VSS
c10 13 VSS 0.00172694f $X=0.081 $Y=0.135
c11 5 VSS 0.00325747f $X=0.081 $Y=0.134
c12 2 VSS 0.0653596f $X=0.081 $Y=0.0675
r13 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.134 $X2=0.081
+ $Y2=0.134
r14 5 7 307.213 $w=2e-08 $l=8.2e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.134 $X2=0.081 $Y2=0.216
r15 2 5 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.134
.ends

.subckt PM_AND5X1_ASAP7_75T_R%B 2 5 7 15 VSS
c12 15 VSS 0.0024522f $X=0.135 $Y=0.135
c13 5 VSS 0.0017107f $X=0.135 $Y=0.1345
c14 2 VSS 0.0604599f $X=0.135 $Y=0.0675
r15 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.134 $X2=0.135
+ $Y2=0.134
r16 5 7 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1345 $X2=0.135 $Y2=0.216
r17 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1345
.ends

.subckt PM_AND5X1_ASAP7_75T_R%C 2 5 7 13 VSS
c11 13 VSS 0.00209947f $X=0.189 $Y=0.135
c12 5 VSS 0.00160244f $X=0.189 $Y=0.1345
c13 2 VSS 0.0597904f $X=0.189 $Y=0.0675
r14 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.134 $X2=0.189
+ $Y2=0.134
r15 5 7 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1345 $X2=0.189 $Y2=0.216
r16 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.1345
.ends

.subckt PM_AND5X1_ASAP7_75T_R%D 2 5 7 13 VSS
c13 13 VSS 0.0024709f $X=0.243 $Y=0.135
c14 5 VSS 0.00160623f $X=0.243 $Y=0.1345
c15 2 VSS 0.059515f $X=0.243 $Y=0.0675
r16 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.134 $X2=0.243
+ $Y2=0.134
r17 5 7 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1345 $X2=0.243 $Y2=0.216
r18 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.1345
.ends

.subckt PM_AND5X1_ASAP7_75T_R%E 2 5 7 15 VSS
c10 15 VSS 0.00305094f $X=0.297 $Y=0.135
c11 5 VSS 0.00162408f $X=0.297 $Y=0.1345
c12 2 VSS 0.0594813f $X=0.297 $Y=0.0675
r13 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.134 $X2=0.297
+ $Y2=0.134
r14 5 7 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.1345 $X2=0.297 $Y2=0.216
r15 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.1345
.ends

.subckt PM_AND5X1_ASAP7_75T_R%8 2 5 7 9 14 17 19 20 23 24 25 28 32 35 36 38 48
+ 50 56 58 61 62 63 65 69 VSS
c32 69 VSS 5.06098e-19 $X=0.351 $Y=0.1765
c33 65 VSS 4.53772e-19 $X=0.351 $Y=0.134
c34 63 VSS 4.85855e-19 $X=0.351 $Y=0.189
c35 62 VSS 1.69932e-19 $X=0.306 $Y=0.198
c36 61 VSS 0.00394258f $X=0.342 $Y=0.198
c37 60 VSS 8.65169e-19 $X=0.297 $Y=0.225
c38 58 VSS 0.00146362f $X=0.252 $Y=0.234
c39 57 VSS 0.00631462f $X=0.234 $Y=0.234
c40 56 VSS 0.00146362f $X=0.198 $Y=0.234
c41 55 VSS 0.00284382f $X=0.18 $Y=0.234
c42 51 VSS 9.64186e-19 $X=0.153 $Y=0.234
c43 50 VSS 0.00142296f $X=0.144 $Y=0.234
c44 49 VSS 0.00636214f $X=0.126 $Y=0.234
c45 48 VSS 0.00142296f $X=0.09 $Y=0.234
c46 47 VSS 1.68773e-19 $X=0.072 $Y=0.234
c47 46 VSS 0.00470185f $X=0.07 $Y=0.234
c48 39 VSS 0.0032477f $X=0.027 $Y=0.234
c49 38 VSS 0.0066498f $X=0.288 $Y=0.234
c50 36 VSS 0.00244555f $X=0.054 $Y=0.036
c51 35 VSS 0.00545273f $X=0.054 $Y=0.036
c52 33 VSS 0.00317163f $X=0.027 $Y=0.036
c53 32 VSS 0.00607891f $X=0.018 $Y=0.2
c54 31 VSS 0.00117262f $X=0.018 $Y=0.07
c55 30 VSS 9.13166e-19 $X=0.018 $Y=0.225
c56 28 VSS 0.00838562f $X=0.27 $Y=0.216
c57 24 VSS 5.3314e-19 $X=0.287 $Y=0.216
c58 23 VSS 0.00791982f $X=0.162 $Y=0.216
c59 19 VSS 5.3314e-19 $X=0.179 $Y=0.216
c60 17 VSS 0.00523518f $X=0.056 $Y=0.216
c61 14 VSS 2.53241e-19 $X=0.071 $Y=0.216
c62 9 VSS 4.49354e-19 $X=0.071 $Y=0.0675
c63 5 VSS 0.00201427f $X=0.351 $Y=0.1345
c64 2 VSS 0.064696f $X=0.351 $Y=0.0675
r65 68 69 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.164 $X2=0.351 $Y2=0.1765
r66 65 68 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.134 $X2=0.351 $Y2=0.164
r67 63 69 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.1765
r68 61 63 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.198 $X2=0.351 $Y2=0.189
r69 61 62 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.306 $Y2=0.198
r70 59 62 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.297 $Y=0.207 $X2=0.306 $Y2=0.198
r71 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.207 $X2=0.297 $Y2=0.225
r72 57 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r73 56 57 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.234 $Y2=0.234
r74 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r75 53 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.252 $Y2=0.234
r76 50 51 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.153 $Y2=0.234
r77 49 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r78 48 49 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.126 $Y2=0.234
r79 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r80 46 47 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.07
+ $Y=0.234 $X2=0.072 $Y2=0.234
r81 44 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r82 44 51 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.153 $Y2=0.234
r83 41 46 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.07 $Y2=0.234
r84 39 41 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.054 $Y2=0.234
r85 38 60 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.234 $X2=0.297 $Y2=0.225
r86 38 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.27 $Y2=0.234
r87 35 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r88 33 35 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.054 $Y2=0.036
r89 31 32 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.2
r90 30 39 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r91 30 32 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2
r92 29 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r93 29 31 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r94 28 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r95 25 28 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.216 $X2=0.27 $Y2=0.216
r96 24 28 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.216 $X2=0.27 $Y2=0.216
r97 23 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234 $X2=0.162
+ $Y2=0.234
r98 20 23 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.216 $X2=0.162 $Y2=0.216
r99 19 23 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.216 $X2=0.162 $Y2=0.216
r100 17 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r101 14 17 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.216 $X2=0.056 $Y2=0.216
r102 12 36 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.054 $Y=0.0675 $X2=0.054 $Y2=0.036
r103 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r104 5 65 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.134 $X2=0.351
+ $Y2=0.134
r105 5 7 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.1345 $X2=0.351 $Y2=0.2025
r106 2 5 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.1345
.ends

.subckt PM_AND5X1_ASAP7_75T_R%Y 1 6 9 13 20 28 29 30 VSS
c10 32 VSS 4.55454e-19 $X=0.405 $Y=0.216
c11 30 VSS 3.02858e-19 $X=0.405 $Y=0.1225
c12 29 VSS 0.00319587f $X=0.405 $Y=0.116
c13 28 VSS 0.00360426f $X=0.409 $Y=0.129
c14 26 VSS 4.30151e-19 $X=0.405 $Y=0.225
c15 21 VSS 0.00612739f $X=0.378 $Y=0.036
c16 20 VSS 0.00269153f $X=0.378 $Y=0.036
c17 18 VSS 0.00601235f $X=0.396 $Y=0.036
c18 13 VSS 0.00275846f $X=0.378 $Y=0.234
c19 11 VSS 0.00601314f $X=0.396 $Y=0.234
c20 9 VSS 0.00665728f $X=0.376 $Y=0.2025
c21 4 VSS 2.69461e-19 $X=0.376 $Y=0.0675
r22 31 32 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.207 $X2=0.405 $Y2=0.216
r23 29 30 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.116 $X2=0.405 $Y2=0.1225
r24 28 31 5.2963 $w=1.8e-08 $l=7.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.129 $X2=0.405 $Y2=0.207
r25 28 30 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.129 $X2=0.405 $Y2=0.1225
r26 26 32 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.216
r27 25 29 4.82099 $w=1.8e-08 $l=7.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.116
r28 20 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r29 18 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r30 18 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.378 $Y2=0.036
r31 11 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r32 11 13 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.378 $Y2=0.234
r33 9 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r34 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.2025 $X2=0.376 $Y2=0.2025
r35 4 21 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r36 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.0675 $X2=0.376 $Y2=0.0675
.ends

.subckt PM_AND5X1_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00228332f $X=0.125 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends

.subckt PM_AND5X1_ASAP7_75T_R%11 1 2 VSS
c0 1 VSS 0.00228332f $X=0.179 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.145 $Y2=0.0675
.ends

.subckt PM_AND5X1_ASAP7_75T_R%12 1 2 VSS
c0 1 VSS 0.00228332f $X=0.233 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.199 $Y2=0.0675
.ends

.subckt PM_AND5X1_ASAP7_75T_R%13 1 2 VSS
c0 1 VSS 0.00228332f $X=0.287 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.253 $Y2=0.0675
.ends


* END of "./AND5x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt AND5x1_ASAP7_75t_R  VSS VDD A B C D E Y
* 
* Y	Y
* E	E
* D	D
* C	C
* B	B
* A	A
M0 N_10_M0_d N_A_M0_g N_8_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_11_M1_d N_B_M1_g N_10_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_12_M2_d N_C_M2_g N_11_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_13_M3_d N_D_M3_g N_12_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 VSS N_E_M4_g N_13_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 N_Y_M5_d N_8_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 VDD N_A_M6_g N_8_M6_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M7 N_8_M7_d N_B_M7_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
M8 VDD N_C_M8_g N_8_M8_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.189
M9 N_8_M9_d N_D_M9_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.189
M10 VDD N_E_M10_g N_8_M10_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287
+ $Y=0.189
M11 N_Y_M11_d N_8_M11_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "AND5x1_ASAP7_75t_R.pex.sp.AND5X1_ASAP7_75T_R.pxi"
* BEGIN of "./AND5x1_ASAP7_75t_R.pex.sp.AND5X1_ASAP7_75T_R.pxi"
* File: AND5x1_ASAP7_75t_R.pex.sp.AND5X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:01:41 2017
* 
x_PM_AND5X1_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M6_g A VSS
+ PM_AND5X1_ASAP7_75T_R%A
x_PM_AND5X1_ASAP7_75T_R%B N_B_M1_g N_B_c_12_n N_B_M7_g B VSS
+ PM_AND5X1_ASAP7_75T_R%B
x_PM_AND5X1_ASAP7_75T_R%C N_C_M2_g N_C_c_25_n N_C_M8_g C VSS
+ PM_AND5X1_ASAP7_75T_R%C
x_PM_AND5X1_ASAP7_75T_R%D N_D_M3_g N_D_c_36_n N_D_M9_g D VSS
+ PM_AND5X1_ASAP7_75T_R%D
x_PM_AND5X1_ASAP7_75T_R%E N_E_M4_g N_E_c_49_n N_E_M10_g E VSS
+ PM_AND5X1_ASAP7_75T_R%E
x_PM_AND5X1_ASAP7_75T_R%8 N_8_M5_g N_8_c_78_n N_8_M11_g N_8_M0_s N_8_M6_s
+ N_8_c_57_n N_8_M8_s N_8_M7_d N_8_c_63_n N_8_M10_s N_8_M9_d N_8_c_72_n
+ N_8_c_58_n N_8_c_64_n N_8_c_59_n N_8_c_83_p N_8_c_61_n N_8_c_66_n N_8_c_69_n
+ N_8_c_73_n N_8_c_84_p N_8_c_75_n N_8_c_87_p N_8_c_80_n N_8_c_76_n VSS
+ PM_AND5X1_ASAP7_75T_R%8
x_PM_AND5X1_ASAP7_75T_R%Y N_Y_M5_d N_Y_M11_d N_Y_c_91_n N_Y_c_92_n N_Y_c_89_n Y
+ N_Y_c_90_n N_Y_c_98_n VSS PM_AND5X1_ASAP7_75T_R%Y
x_PM_AND5X1_ASAP7_75T_R%10 N_10_M1_s N_10_M0_d VSS PM_AND5X1_ASAP7_75T_R%10
x_PM_AND5X1_ASAP7_75T_R%11 N_11_M2_s N_11_M1_d VSS PM_AND5X1_ASAP7_75T_R%11
x_PM_AND5X1_ASAP7_75T_R%12 N_12_M3_s N_12_M2_d VSS PM_AND5X1_ASAP7_75T_R%12
x_PM_AND5X1_ASAP7_75T_R%13 N_13_M4_s N_13_M3_d VSS PM_AND5X1_ASAP7_75T_R%13
cc_1 N_A_M0_g N_B_M1_g 0.00333077f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_12_n 7.98811e-19 $X=0.081 $Y=0.134 $X2=0.135 $Y2=0.1345
cc_3 A B 0.00621434f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A_M0_g N_C_M2_g 2.71887e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 A N_8_c_57_n 3.52002e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_6 A N_8_c_58_n 0.00436697f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_7 N_A_c_2_p N_8_c_59_n 3.06446e-19 $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_8 A N_8_c_59_n 0.00134508f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_A_M0_g N_8_c_61_n 2.57864e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_10 A N_8_c_61_n 0.00123648f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 N_B_M1_g N_C_M2_g 0.00357042f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_12 N_B_c_12_n N_C_c_25_n 7.92653e-19 $X=0.135 $Y=0.1345 $X2=0.081 $Y2=0.134
cc_13 B C 0.00817592f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 N_B_M1_g N_D_M3_g 2.71887e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_15 B N_8_c_63_n 3.31541e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_16 B N_8_c_64_n 4.64233e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_17 B N_8_c_59_n 5.56013e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_18 N_B_M1_g N_8_c_66_n 2.57565e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 B N_8_c_66_n 0.00123952f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_20 N_C_M2_g N_D_M3_g 0.00327995f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_21 N_C_c_25_n N_D_c_36_n 7.90494e-19 $X=0.189 $Y=0.1345 $X2=0.081 $Y2=0.134
cc_22 C D 0.00817682f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 N_C_M2_g N_E_M4_g 2.66145e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_24 C N_8_c_63_n 3.31541e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_25 N_C_M2_g N_8_c_69_n 2.64924e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 C N_8_c_69_n 0.00125705f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_27 N_D_M3_g N_E_M4_g 0.00344695f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_28 N_D_c_36_n N_E_c_49_n 7.90494e-19 $X=0.243 $Y=0.1345 $X2=0.135 $Y2=0.1345
cc_29 D E 0.00646431f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_30 N_D_M3_g N_8_M5_g 2.31381e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_31 D N_8_c_72_n 3.24828e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_32 N_D_M3_g N_8_c_73_n 2.64924e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_33 D N_8_c_73_n 0.00125705f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_34 D N_8_c_75_n 4.59663e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_35 D N_8_c_76_n 2.69033e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_36 N_E_M4_g N_8_M5_g 0.00284417f $X=0.297 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_37 N_E_c_49_n N_8_c_78_n 8.31912e-19 $X=0.297 $Y=0.1345 $X2=0.189 $Y2=0.1345
cc_38 E N_8_c_75_n 0.00135016f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_39 E N_8_c_80_n 0.00215568f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_40 E N_Y_c_89_n 3.55123e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_41 E N_Y_c_90_n 4.71495e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_42 N_8_c_80_n N_Y_c_91_n 0.00135034f $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_43 N_8_M5_g N_Y_c_92_n 2.56972e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_44 N_8_c_83_p N_Y_c_92_n 5.2369e-19 $X=0.288 $Y=0.234 $X2=0.081 $Y2=0.135
cc_45 N_8_c_84_p N_Y_c_92_n 0.00100131f $X=0.342 $Y=0.198 $X2=0.081 $Y2=0.135
cc_46 N_8_M5_g N_Y_c_89_n 3.02028e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_8_c_80_n N_Y_c_89_n 2.49025e-19 $X=0.351 $Y=0.134 $X2=0 $Y2=0
cc_48 N_8_c_87_p Y 0.0018612f $X=0.351 $Y=0.189 $X2=0 $Y2=0
cc_49 N_8_c_80_n N_Y_c_98_n 0.0018612f $X=0.351 $Y=0.134 $X2=0 $Y2=0

* END of "./AND5x1_ASAP7_75t_R.pex.sp.AND5X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: AND5x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:02:04 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "AND5x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./AND5x2_ASAP7_75t_R.pex.sp.pex"
* File: AND5x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:02:04 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_AND5X2_ASAP7_75T_R%E 2 8 11 13 30 VSS
c4 30 VSS 0.0203548f $X=0.08 $Y=0.137
c5 11 VSS 0.00958217f $X=0.135 $Y=0.135
c6 8 VSS 0.0668902f $X=0.135 $Y=0.0675
c7 2 VSS 0.0670595f $X=0.081 $Y=0.0675
r8 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r9 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
r10 5 11 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081 $Y=0.135
+ $X2=0.135 $Y2=0.135
r11 5 30 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r12 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_AND5X2_ASAP7_75T_R%D 2 7 10 13 22 VSS
c19 22 VSS 0.00420967f $X=0.296 $Y=0.137
c20 13 VSS 0.0069115f $X=0.351 $Y=0.135
c21 10 VSS 0.0640309f $X=0.351 $Y=0.0675
c22 2 VSS 0.0673211f $X=0.297 $Y=0.0675
r23 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r24 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297 $Y=0.135
+ $X2=0.351 $Y2=0.135
r25 5 22 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r26 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r27 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_AND5X2_ASAP7_75T_R%C 2 8 11 13 20 VSS
c21 20 VSS 0.00395043f $X=0.458 $Y=0.137
c22 11 VSS 0.00422108f $X=0.459 $Y=0.135
c23 8 VSS 0.0661608f $X=0.459 $Y=0.0675
c24 2 VSS 0.063631f $X=0.405 $Y=0.0675
r25 11 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r26 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r27 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r28 5 11 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405 $Y=0.135
+ $X2=0.459 $Y2=0.135
r29 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_AND5X2_ASAP7_75T_R%B 2 7 10 13 20 VSS
c20 20 VSS 0.00332483f $X=0.62 $Y=0.137
c21 13 VSS 0.0069009f $X=0.675 $Y=0.135
c22 10 VSS 0.0640309f $X=0.675 $Y=0.0675
c23 2 VSS 0.0672745f $X=0.621 $Y=0.0675
r24 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0675 $X2=0.675 $Y2=0.135
r25 5 13 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.621 $Y=0.135
+ $X2=0.675 $Y2=0.135
r26 5 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r27 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.2025
r28 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.621
+ $Y=0.0675 $X2=0.621 $Y2=0.135
.ends

.subckt PM_AND5X2_ASAP7_75T_R%A 2 8 11 13 20 VSS
c23 20 VSS 0.00247178f $X=0.728 $Y=0.137
c24 11 VSS 0.00356163f $X=0.783 $Y=0.135
c25 8 VSS 0.0655947f $X=0.783 $Y=0.0675
c26 2 VSS 0.0632415f $X=0.729 $Y=0.0675
r27 11 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.135 $X2=0.783 $Y2=0.2025
r28 8 11 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.783
+ $Y=0.0675 $X2=0.783 $Y2=0.135
r29 5 11 54 $w=2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.729 $Y=0.135
+ $X2=0.783 $Y2=0.135
r30 5 20 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.729 $Y=0.135 $X2=0.729
+ $Y2=0.135
r31 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.729
+ $Y=0.0675 $X2=0.729 $Y2=0.135
.ends

.subckt PM_AND5X2_ASAP7_75T_R%8 2 7 10 13 15 17 18 22 27 30 32 35 37 40 42 45 47
+ 55 56 60 61 65 66 67 69 74 75 76 77 78 81 83 86 88 89 93 VSS
c67 100 VSS 3.92668e-19 $X=0.891 $Y=0.135
c68 97 VSS 0.00210915f $X=0.928 $Y=0.135
c69 94 VSS 0.00155658f $X=0.891 $Y=0.207
c70 93 VSS 0.00278763f $X=0.891 $Y=0.189
c71 92 VSS 0.00109324f $X=0.891 $Y=0.225
c72 90 VSS 0.00104577f $X=0.891 $Y=0.117
c73 89 VSS 0.00101345f $X=0.891 $Y=0.099
c74 88 VSS 0.0011573f $X=0.891 $Y=0.081
c75 87 VSS 0.00109324f $X=0.891 $Y=0.063
c76 86 VSS 3.85713e-19 $X=0.891 $Y=0.126
c77 84 VSS 0.00376564f $X=0.853 $Y=0.036
c78 83 VSS 0.00690555f $X=0.824 $Y=0.036
c79 81 VSS 0.00317566f $X=0.756 $Y=0.036
c80 78 VSS 0.00676815f $X=0.882 $Y=0.036
c81 77 VSS 0.0091941f $X=0.824 $Y=0.234
c82 76 VSS 0.00294577f $X=0.757 $Y=0.234
c83 75 VSS 0.0115403f $X=0.72 $Y=0.234
c84 74 VSS 0.00286286f $X=0.63 $Y=0.234
c85 69 VSS 0.00127724f $X=0.593 $Y=0.234
c86 68 VSS 0.0101873f $X=0.58 $Y=0.234
c87 67 VSS 0.00297135f $X=0.5 $Y=0.234
c88 66 VSS 0.00429135f $X=0.487 $Y=0.234
c89 65 VSS 0.00729429f $X=0.45 $Y=0.234
c90 61 VSS 0.00886827f $X=0.369 $Y=0.234
c91 60 VSS 0.00290097f $X=0.306 $Y=0.234
c92 56 VSS 0.00133102f $X=0.269 $Y=0.234
c93 55 VSS 0.014063f $X=0.256 $Y=0.234
c94 47 VSS 0.0105409f $X=0.882 $Y=0.234
c95 45 VSS 0.00874174f $X=0.758 $Y=0.2025
c96 42 VSS 4.53693e-19 $X=0.773 $Y=0.2025
c97 40 VSS 0.00833579f $X=0.596 $Y=0.2025
c98 37 VSS 3.00769e-19 $X=0.611 $Y=0.2025
c99 35 VSS 0.00804325f $X=0.434 $Y=0.2025
c100 32 VSS 4.53693e-19 $X=0.449 $Y=0.2025
c101 30 VSS 0.00719038f $X=0.272 $Y=0.2025
c102 27 VSS 3.00769e-19 $X=0.287 $Y=0.2025
c103 25 VSS 0.00698584f $X=0.16 $Y=0.2025
c104 17 VSS 6.7506e-19 $X=0.773 $Y=0.0675
c105 13 VSS 0.00765919f $X=0.999 $Y=0.135
c106 10 VSS 0.0641916f $X=0.999 $Y=0.0675
c107 2 VSS 0.065064f $X=0.945 $Y=0.0675
r108 97 98 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.928 $Y=0.135 $X2=0.928
+ $Y2=0.135
r109 95 100 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.135 $X2=0.891 $Y2=0.135
r110 95 97 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.9
+ $Y=0.135 $X2=0.928 $Y2=0.135
r111 93 94 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.189 $X2=0.891 $Y2=0.207
r112 92 94 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.225 $X2=0.891 $Y2=0.207
r113 91 100 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.144 $X2=0.891 $Y2=0.135
r114 91 93 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.144 $X2=0.891 $Y2=0.189
r115 89 90 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.099 $X2=0.891 $Y2=0.117
r116 88 89 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.081 $X2=0.891 $Y2=0.099
r117 87 88 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.063 $X2=0.891 $Y2=0.081
r118 86 100 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.126 $X2=0.891 $Y2=0.135
r119 86 90 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.126 $X2=0.891 $Y2=0.117
r120 85 87 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.891
+ $Y=0.045 $X2=0.891 $Y2=0.063
r121 83 84 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.824
+ $Y=0.036 $X2=0.853 $Y2=0.036
r122 80 83 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.036 $X2=0.824 $Y2=0.036
r123 80 81 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.036
+ $X2=0.756 $Y2=0.036
r124 78 85 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.036 $X2=0.891 $Y2=0.045
r125 78 84 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.036 $X2=0.853 $Y2=0.036
r126 76 77 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.757
+ $Y=0.234 $X2=0.824 $Y2=0.234
r127 74 75 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.234 $X2=0.72 $Y2=0.234
r128 72 76 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.757 $Y2=0.234
r129 72 75 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.756
+ $Y=0.234 $X2=0.72 $Y2=0.234
r130 69 70 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.593
+ $Y=0.234 $X2=0.5935 $Y2=0.234
r131 68 69 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.58
+ $Y=0.234 $X2=0.593 $Y2=0.234
r132 67 68 5.4321 $w=1.8e-08 $l=8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5
+ $Y=0.234 $X2=0.58 $Y2=0.234
r133 66 67 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.487
+ $Y=0.234 $X2=0.5 $Y2=0.234
r134 65 66 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.487 $Y2=0.234
r135 63 74 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.63 $Y2=0.234
r136 63 70 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.5935 $Y2=0.234
r137 60 61 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.234 $X2=0.369 $Y2=0.234
r138 58 65 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.45 $Y2=0.234
r139 58 61 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.369 $Y2=0.234
r140 55 56 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.234 $X2=0.269 $Y2=0.234
r141 53 60 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.306 $Y2=0.234
r142 53 56 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.269 $Y2=0.234
r143 49 55 6.38272 $w=1.8e-08 $l=9.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.256 $Y2=0.234
r144 47 92 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.882 $Y=0.234 $X2=0.891 $Y2=0.225
r145 47 77 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.882
+ $Y=0.234 $X2=0.824 $Y2=0.234
r146 45 72 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.756 $Y=0.234
+ $X2=0.756 $Y2=0.234
r147 42 45 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.2025 $X2=0.758 $Y2=0.2025
r148 40 63 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234
+ $X2=0.594 $Y2=0.234
r149 37 40 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.611 $Y=0.2025 $X2=0.596 $Y2=0.2025
r150 35 58 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234
+ $X2=0.432 $Y2=0.234
r151 32 35 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.434 $Y2=0.2025
r152 30 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r153 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.272 $Y2=0.2025
r154 25 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.234
+ $X2=0.162 $Y2=0.234
r155 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.16 $Y2=0.2025
r156 21 81 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.756 $Y=0.0675 $X2=0.756 $Y2=0.036
r157 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.739 $Y=0.0675 $X2=0.756 $Y2=0.0675
r158 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.773 $Y=0.0675 $X2=0.756 $Y2=0.0675
r159 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.135 $X2=0.999 $Y2=0.2025
r160 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.999 $Y=0.0675 $X2=0.999 $Y2=0.135
r161 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.945
+ $Y=0.135 $X2=0.999 $Y2=0.135
r162 5 98 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.945
+ $Y=0.135 $X2=0.928 $Y2=0.135
r163 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.945
+ $Y=0.135 $X2=0.945 $Y2=0.2025
r164 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.945
+ $Y=0.0675 $X2=0.945 $Y2=0.135
.ends

.subckt PM_AND5X2_ASAP7_75T_R%9 1 2 6 7 12 13 18 19 20 21 VSS
c18 21 VSS 0.0159468f $X=0.256 $Y=0.036
c19 20 VSS 0.0043517f $X=0.148 $Y=0.036
c20 19 VSS 0.00510681f $X=0.324 $Y=0.036
c21 18 VSS 0.0068994f $X=0.324 $Y=0.036
c22 13 VSS 0.0102758f $X=0.108 $Y=0.036
c23 12 VSS 0.00174603f $X=0.108 $Y=0.036
c24 6 VSS 6.4978e-19 $X=0.341 $Y=0.0675
c25 1 VSS 5.58795e-19 $X=0.125 $Y=0.0675
r26 20 21 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.148
+ $Y=0.036 $X2=0.256 $Y2=0.036
r27 18 21 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.256 $Y2=0.036
r28 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r29 12 20 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.148 $Y2=0.036
r30 12 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r31 10 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r32 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r33 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r34 5 13 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r35 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r36 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends

.subckt PM_AND5X2_ASAP7_75T_R%10 1 4 6 7 10 11 14 17 25 26 28 30 31 VSS
c30 31 VSS 2.77631e-19 $X=0.45 $Y=0.072
c31 30 VSS 0.00323868f $X=0.418 $Y=0.072
c32 28 VSS 6.81795e-19 $X=0.486 $Y=0.072
c33 26 VSS 2.77631e-19 $X=0.338 $Y=0.072
c34 25 VSS 8.46035e-21 $X=0.306 $Y=0.072
c35 17 VSS 7.71579e-19 $X=0.27 $Y=0.072
c36 14 VSS 0.0041846f $X=0.484 $Y=0.0675
c37 10 VSS 7.08605e-19 $X=0.378 $Y=0.0675
c38 6 VSS 6.69874e-19 $X=0.395 $Y=0.0675
c39 4 VSS 0.00440468f $X=0.272 $Y=0.0675
c40 1 VSS 3.32862e-19 $X=0.287 $Y=0.0675
r41 30 31 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.418
+ $Y=0.072 $X2=0.45 $Y2=0.072
r42 28 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.072 $X2=0.45 $Y2=0.072
r43 25 26 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.072 $X2=0.338 $Y2=0.072
r44 23 30 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.418 $Y2=0.072
r45 23 26 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.338 $Y2=0.072
r46 17 25 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.072 $X2=0.306 $Y2=0.072
r47 14 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.072 $X2=0.486
+ $Y2=0.072
r48 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.484 $Y2=0.0675
r49 10 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.072 $X2=0.378
+ $Y2=0.072
r50 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.378 $Y2=0.0675
r51 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.0675 $X2=0.378 $Y2=0.0675
r52 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.072 $X2=0.27
+ $Y2=0.072
r53 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.272 $Y2=0.0675
.ends

.subckt PM_AND5X2_ASAP7_75T_R%11 1 2 6 7 13 16 17 18 19 VSS
c27 19 VSS 0.0101873f $X=0.58 $Y=0.036
c28 18 VSS 0.00686773f $X=0.5 $Y=0.036
c29 17 VSS 0.00488896f $X=0.648 $Y=0.036
c30 16 VSS 0.0068994f $X=0.648 $Y=0.036
c31 13 VSS 0.00296838f $X=0.432 $Y=0.036
c32 6 VSS 6.4978e-19 $X=0.665 $Y=0.0675
c33 1 VSS 6.4978e-19 $X=0.449 $Y=0.0675
r34 18 19 5.4321 $w=1.8e-08 $l=8e-08 $layer=M1 $thickness=3.6e-08 $X=0.5
+ $Y=0.036 $X2=0.58 $Y2=0.036
r35 16 19 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.58 $Y2=0.036
r36 16 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036 $X2=0.648
+ $Y2=0.036
r37 12 18 4.61728 $w=1.8e-08 $l=6.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.5 $Y2=0.036
r38 12 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r39 10 17 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.648
+ $Y=0.0675 $X2=0.648 $Y2=0.036
r40 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.648 $Y2=0.0675
r41 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0675 $X2=0.648 $Y2=0.0675
r42 5 13 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r43 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.432 $Y2=0.0675
r44 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.449
+ $Y=0.0675 $X2=0.432 $Y2=0.0675
.ends

.subckt PM_AND5X2_ASAP7_75T_R%12 1 4 6 7 10 11 14 17 25 26 28 30 31 32 33 VSS
c32 33 VSS 1.88159e-19 $X=0.7835 $Y=0.072
c33 32 VSS 1.37234e-20 $X=0.757 $Y=0.072
c34 31 VSS 6.62855e-19 $X=0.742 $Y=0.072
c35 30 VSS 0.00249766f $X=0.72 $Y=0.072
c36 28 VSS 0.0011408f $X=0.81 $Y=0.072
c37 26 VSS 2.77631e-19 $X=0.662 $Y=0.072
c38 25 VSS 8.46035e-21 $X=0.63 $Y=0.072
c39 17 VSS 6.19631e-19 $X=0.594 $Y=0.072
c40 14 VSS 0.00610772f $X=0.808 $Y=0.0675
c41 10 VSS 7.09451e-19 $X=0.702 $Y=0.0675
c42 6 VSS 6.69874e-19 $X=0.719 $Y=0.0675
c43 4 VSS 0.00297328f $X=0.596 $Y=0.0675
c44 1 VSS 3.32862e-19 $X=0.611 $Y=0.0675
r45 32 33 1.79938 $w=1.8e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.757
+ $Y=0.072 $X2=0.7835 $Y2=0.072
r46 31 32 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.742
+ $Y=0.072 $X2=0.757 $Y2=0.072
r47 30 31 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.72
+ $Y=0.072 $X2=0.742 $Y2=0.072
r48 28 33 1.79938 $w=1.8e-08 $l=2.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.81
+ $Y=0.072 $X2=0.7835 $Y2=0.072
r49 25 26 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.63
+ $Y=0.072 $X2=0.662 $Y2=0.072
r50 23 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.072 $X2=0.72 $Y2=0.072
r51 23 26 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.702
+ $Y=0.072 $X2=0.662 $Y2=0.072
r52 17 25 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.072 $X2=0.63 $Y2=0.072
r53 14 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.81 $Y=0.072 $X2=0.81
+ $Y2=0.072
r54 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.793 $Y=0.0675 $X2=0.808 $Y2=0.0675
r55 10 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.702 $Y=0.072 $X2=0.702
+ $Y2=0.072
r56 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.685 $Y=0.0675 $X2=0.702 $Y2=0.0675
r57 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.719 $Y=0.0675 $X2=0.702 $Y2=0.0675
r58 4 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.072 $X2=0.594
+ $Y2=0.072
r59 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.611
+ $Y=0.0675 $X2=0.596 $Y2=0.0675
.ends

.subckt PM_AND5X2_ASAP7_75T_R%Y 1 2 6 7 10 11 14 16 24 25 VSS
c13 26 VSS 9.7518e-19 $X=1.053 $Y=0.144
c14 25 VSS 0.0046845f $X=1.053 $Y=0.126
c15 24 VSS 0.0046845f $X=1.053 $Y=0.1475
c16 16 VSS 0.0145473f $X=1.044 $Y=0.234
c17 14 VSS 0.00914518f $X=0.972 $Y=0.036
c18 11 VSS 0.0145473f $X=1.044 $Y=0.036
c19 10 VSS 0.00931384f $X=0.972 $Y=0.2025
c20 6 VSS 5.72268e-19 $X=0.989 $Y=0.2025
c21 1 VSS 5.72268e-19 $X=0.989 $Y=0.0675
r22 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.126 $X2=1.053 $Y2=0.144
r23 24 26 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.1475 $X2=1.053 $Y2=0.144
r24 22 24 5.26235 $w=1.8e-08 $l=7.75e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.225 $X2=1.053 $Y2=0.1475
r25 21 25 5.5 $w=1.8e-08 $l=8.1e-08 $layer=M1 $thickness=3.6e-08 $X=1.053
+ $Y=0.045 $X2=1.053 $Y2=0.126
r26 16 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.234 $X2=1.053 $Y2=0.225
r27 16 18 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.234 $X2=0.972 $Y2=0.234
r28 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.036 $X2=0.972
+ $Y2=0.036
r29 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=1.044 $Y=0.036 $X2=1.053 $Y2=0.045
r30 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=1.044
+ $Y=0.036 $X2=0.972 $Y2=0.036
r31 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.972 $Y=0.234 $X2=0.972
+ $Y2=0.234
r32 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.955 $Y=0.2025 $X2=0.972 $Y2=0.2025
r33 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.989 $Y=0.2025 $X2=0.972 $Y2=0.2025
r34 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.972
+ $Y=0.0675 $X2=0.972 $Y2=0.036
r35 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.955
+ $Y=0.0675 $X2=0.972 $Y2=0.0675
r36 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.989
+ $Y=0.0675 $X2=0.972 $Y2=0.0675
.ends


* END of "./AND5x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt AND5x2_ASAP7_75t_R  VSS VDD E D C B A Y
* 
* Y	Y
* A	A
* B	B
* C	C
* D	D
* E	E
M0 N_9_M0_d N_E_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_9_M1_d N_E_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_9_M2_d N_D_M2_g N_10_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 N_9_M3_d N_D_M3_g N_10_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 N_11_M4_d N_C_M4_g N_10_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 N_11_M5_d N_C_M5_g N_10_M5_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 N_11_M6_d N_B_M6_g N_12_M6_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M7 N_11_M7_d N_B_M7_g N_12_M7_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M8 N_8_M8_d N_A_M8_g N_12_M8_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.719
+ $Y=0.027
M9 N_8_M9_d N_A_M9_g N_12_M9_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.027
M10 N_Y_M10_d N_8_M10_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.027
M11 N_Y_M11_d N_8_M11_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.027
M12 N_8_M12_d N_E_M12_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M13 VDD N_D_M13_g N_8_M13_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M14 VDD N_C_M14_g N_8_M14_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M15 VDD N_B_M15_g N_8_M15_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M16 VDD N_A_M16_g N_8_M16_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.773
+ $Y=0.162
M17 N_Y_M17_d N_8_M17_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.935
+ $Y=0.162
M18 N_Y_M18_d N_8_M18_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.989
+ $Y=0.162
*
* 
* .include "AND5x2_ASAP7_75t_R.pex.sp.AND5X2_ASAP7_75T_R.pxi"
* BEGIN of "./AND5x2_ASAP7_75t_R.pex.sp.AND5X2_ASAP7_75T_R.pxi"
* File: AND5x2_ASAP7_75t_R.pex.sp.AND5X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:02:04 2017
* 
x_PM_AND5X2_ASAP7_75T_R%E N_E_M0_g N_E_M1_g N_E_c_1_p N_E_M12_g E VSS
+ PM_AND5X2_ASAP7_75T_R%E
x_PM_AND5X2_ASAP7_75T_R%D N_D_M2_g N_D_M13_g N_D_M3_g N_D_c_8_p D VSS
+ PM_AND5X2_ASAP7_75T_R%D
x_PM_AND5X2_ASAP7_75T_R%C N_C_M4_g N_C_M5_g N_C_c_27_n N_C_M14_g C VSS
+ PM_AND5X2_ASAP7_75T_R%C
x_PM_AND5X2_ASAP7_75T_R%B N_B_M6_g N_B_M15_g N_B_M7_g N_B_c_49_p B VSS
+ PM_AND5X2_ASAP7_75T_R%B
x_PM_AND5X2_ASAP7_75T_R%A N_A_M8_g N_A_M9_g N_A_c_68_n N_A_M16_g A VSS
+ PM_AND5X2_ASAP7_75T_R%A
x_PM_AND5X2_ASAP7_75T_R%8 N_8_M10_g N_8_M17_g N_8_M11_g N_8_c_104_n N_8_M18_g
+ N_8_M9_d N_8_M8_d N_8_M12_d N_8_M13_s N_8_c_88_n N_8_M14_s N_8_c_93_n
+ N_8_M15_s N_8_c_99_n N_8_M16_s N_8_c_107_n N_8_c_151_p N_8_c_118_p N_8_c_117_p
+ N_8_c_89_n N_8_c_91_n N_8_c_95_n N_8_c_97_n N_8_c_123_p N_8_c_125_p
+ N_8_c_100_n N_8_c_102_n N_8_c_109_n N_8_c_111_n N_8_c_147_p N_8_c_113_n
+ N_8_c_115_n N_8_c_116_n N_8_c_137_p N_8_c_134_p N_8_c_152_p VSS
+ PM_AND5X2_ASAP7_75T_R%8
x_PM_AND5X2_ASAP7_75T_R%9 N_9_M1_d N_9_M0_d N_9_M3_d N_9_M2_d N_9_c_156_n
+ N_9_c_157_n N_9_c_160_n N_9_c_161_n N_9_c_158_n N_9_c_164_n VSS
+ PM_AND5X2_ASAP7_75T_R%9
x_PM_AND5X2_ASAP7_75T_R%10 N_10_M2_s N_10_c_173_n N_10_M4_s N_10_M3_s
+ N_10_c_191_n N_10_M5_s N_10_c_178_n N_10_c_184_n N_10_c_174_n N_10_c_176_n
+ N_10_c_179_n N_10_c_177_n N_10_c_187_n VSS PM_AND5X2_ASAP7_75T_R%10
x_PM_AND5X2_ASAP7_75T_R%11 N_11_M5_d N_11_M4_d N_11_M7_d N_11_M6_d N_11_c_204_n
+ N_11_c_208_n N_11_c_209_n N_11_c_206_n N_11_c_215_n VSS
+ PM_AND5X2_ASAP7_75T_R%11
x_PM_AND5X2_ASAP7_75T_R%12 N_12_M6_s N_12_c_230_n N_12_M8_s N_12_M7_s
+ N_12_c_235_n N_12_M9_s N_12_c_243_n N_12_c_246_n N_12_c_231_n N_12_c_233_n
+ N_12_c_248_n N_12_c_234_n N_12_c_236_n N_12_c_249_n N_12_c_238_n VSS
+ PM_AND5X2_ASAP7_75T_R%12
x_PM_AND5X2_ASAP7_75T_R%Y N_Y_M11_d N_Y_M10_d N_Y_M18_d N_Y_M17_d N_Y_c_264_n
+ N_Y_c_265_n N_Y_c_268_n N_Y_c_269_n Y N_Y_c_273_n VSS PM_AND5X2_ASAP7_75T_R%Y
cc_1 N_E_c_1_p N_9_M1_d 3.68024e-19 $X=0.135 $Y=0.135 $X2=0.297 $Y2=0.0675
cc_2 N_E_c_1_p N_9_c_156_n 8.1394e-19 $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.135
cc_3 N_E_c_1_p N_9_c_157_n 7.57503e-19 $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.135
cc_4 N_E_M1_g N_9_c_158_n 2.6792e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_5 N_D_M2_g N_C_M4_g 2.71887e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_6 N_D_M3_g N_C_M4_g 0.00364308f $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_7 N_D_M3_g N_C_M5_g 3.00908e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_8 N_D_c_8_p N_C_c_27_n 0.00146676f $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_9 D C 7.05261e-19 $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_10 D N_8_c_88_n 0.00157973f $X=0.296 $Y=0.137 $X2=0.08 $Y2=0.137
cc_11 N_D_M2_g N_8_c_89_n 2.35211e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_12 D N_8_c_89_n 0.00374076f $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_13 N_D_M3_g N_8_c_91_n 4.65034e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_14 N_D_c_8_p N_8_c_91_n 7.23712e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_15 N_D_c_8_p N_9_M3_d 3.67193e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_16 N_D_M2_g N_9_c_160_n 2.38524e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_17 N_D_c_8_p N_9_c_161_n 7.57503e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_18 D N_9_c_161_n 3.21662e-19 $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_19 D N_10_c_173_n 8.82271e-19 $X=0.296 $Y=0.137 $X2=0.081 $Y2=0.135
cc_20 N_D_M2_g N_10_c_174_n 2.53669e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_21 D N_10_c_174_n 0.00372053f $X=0.296 $Y=0.137 $X2=0 $Y2=0
cc_22 N_D_c_8_p N_10_c_176_n 8.63627e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_23 N_D_M3_g N_10_c_177_n 4.96522e-19 $X=0.351 $Y=0.0675 $X2=0.08 $Y2=0.137
cc_24 C B 6.44218e-19 $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_25 N_C_c_27_n N_8_c_93_n 7.57503e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_26 C N_8_c_93_n 0.00157927f $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_27 N_C_M4_g N_8_c_95_n 4.65034e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_28 N_C_c_27_n N_8_c_95_n 4.9959e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_29 N_C_M5_g N_8_c_97_n 2.38524e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_30 C N_8_c_97_n 0.00376514f $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_31 C N_10_c_178_n 9.78138e-19 $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_32 N_C_M5_g N_10_c_179_n 2.53669e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_33 C N_10_c_179_n 0.00373988f $X=0.458 $Y=0.137 $X2=0 $Y2=0
cc_34 N_C_M4_g N_10_c_177_n 4.96522e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_C_c_27_n N_10_c_177_n 8.63627e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_36 N_C_c_27_n N_11_M5_d 3.67193e-19 $X=0.459 $Y=0.135 $X2=0.297 $Y2=0.0675
cc_37 N_C_c_27_n N_11_c_204_n 7.57503e-19 $X=0.459 $Y=0.135 $X2=0.351 $Y2=0.135
cc_38 C N_11_c_204_n 3.21662e-19 $X=0.458 $Y=0.137 $X2=0.351 $Y2=0.135
cc_39 N_C_M5_g N_11_c_206_n 2.38524e-19 $X=0.459 $Y=0.0675 $X2=0.297 $Y2=0.135
cc_40 N_B_M6_g N_A_M8_g 2.71887e-19 $X=0.621 $Y=0.0675 $X2=0.405 $Y2=0.0675
cc_41 N_B_M7_g N_A_M8_g 0.00364308f $X=0.675 $Y=0.0675 $X2=0.405 $Y2=0.0675
cc_42 N_B_M7_g N_A_M9_g 3.00908e-19 $X=0.675 $Y=0.0675 $X2=0.459 $Y2=0.0675
cc_43 N_B_c_49_p N_A_c_68_n 0.00121307f $X=0.675 $Y=0.135 $X2=0.459 $Y2=0.135
cc_44 B A 0.00162725f $X=0.62 $Y=0.137 $X2=0.458 $Y2=0.137
cc_45 B N_8_c_99_n 0.00219806f $X=0.62 $Y=0.137 $X2=0 $Y2=0
cc_46 N_B_M6_g N_8_c_100_n 2.35211e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_47 B N_8_c_100_n 0.00372141f $X=0.62 $Y=0.137 $X2=0 $Y2=0
cc_48 N_B_M7_g N_8_c_102_n 4.65034e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_49 N_B_c_49_p N_8_c_102_n 7.23712e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_50 N_B_c_49_p N_11_M7_d 3.67193e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_51 N_B_M6_g N_11_c_208_n 2.38524e-19 $X=0.621 $Y=0.0675 $X2=0 $Y2=0
cc_52 N_B_c_49_p N_11_c_209_n 7.57503e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_53 B N_11_c_209_n 3.18961e-19 $X=0.62 $Y=0.137 $X2=0 $Y2=0
cc_54 B N_12_c_230_n 9.69496e-19 $X=0.62 $Y=0.137 $X2=0.405 $Y2=0.135
cc_55 N_B_M6_g N_12_c_231_n 2.53669e-19 $X=0.621 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_56 B N_12_c_231_n 0.00372053f $X=0.62 $Y=0.137 $X2=0.405 $Y2=0.135
cc_57 N_B_c_49_p N_12_c_233_n 8.63627e-19 $X=0.675 $Y=0.135 $X2=0 $Y2=0
cc_58 N_B_M7_g N_12_c_234_n 4.96522e-19 $X=0.675 $Y=0.0675 $X2=0 $Y2=0
cc_59 N_A_c_68_n N_8_c_104_n 2.44309e-19 $X=0.783 $Y=0.135 $X2=0.675 $Y2=0.135
cc_60 N_A_c_68_n N_8_M9_d 3.65696e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_61 A N_8_M16_s 2.0764e-19 $X=0.728 $Y=0.137 $X2=0 $Y2=0
cc_62 N_A_c_68_n N_8_c_107_n 7.57503e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_63 A N_8_c_107_n 0.00231513f $X=0.728 $Y=0.137 $X2=0 $Y2=0
cc_64 N_A_M8_g N_8_c_109_n 2.35211e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_65 A N_8_c_109_n 0.00371855f $X=0.728 $Y=0.137 $X2=0 $Y2=0
cc_66 N_A_M9_g N_8_c_111_n 4.65034e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_67 N_A_c_68_n N_8_c_111_n 3.46051e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_68 N_A_c_68_n N_8_c_113_n 7.57503e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_69 A N_8_c_113_n 8.71019e-19 $X=0.728 $Y=0.137 $X2=0 $Y2=0
cc_70 N_A_M9_g N_8_c_115_n 2.65027e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_71 A N_8_c_116_n 4.64816e-19 $X=0.728 $Y=0.137 $X2=0 $Y2=0
cc_72 A N_12_c_235_n 3.18961e-19 $X=0.728 $Y=0.137 $X2=0.675 $Y2=0.0675
cc_73 N_A_M8_g N_12_c_236_n 3.43086e-19 $X=0.729 $Y=0.0675 $X2=0 $Y2=0
cc_74 A N_12_c_236_n 0.00373368f $X=0.728 $Y=0.137 $X2=0 $Y2=0
cc_75 N_A_M9_g N_12_c_238_n 2.10599e-19 $X=0.783 $Y=0.0675 $X2=0 $Y2=0
cc_76 N_A_c_68_n N_12_c_238_n 5.60103e-19 $X=0.783 $Y=0.135 $X2=0 $Y2=0
cc_77 N_8_c_117_p N_9_c_160_n 5.01308e-19 $X=0.269 $Y=0.234 $X2=0 $Y2=0
cc_78 N_8_c_118_p N_9_c_164_n 5.01308e-19 $X=0.256 $Y=0.234 $X2=0 $Y2=0
cc_79 N_8_c_88_n N_10_c_173_n 0.00134615f $X=0.272 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_80 N_8_c_117_p N_10_c_184_n 3.02179e-19 $X=0.269 $Y=0.234 $X2=0 $Y2=0
cc_81 N_8_c_91_n N_10_c_176_n 3.02179e-19 $X=0.369 $Y=0.234 $X2=0 $Y2=0
cc_82 N_8_c_95_n N_10_c_177_n 3.02179e-19 $X=0.45 $Y=0.234 $X2=0.08 $Y2=0.137
cc_83 N_8_c_123_p N_10_c_187_n 3.02179e-19 $X=0.5 $Y=0.234 $X2=0.081 $Y2=0.135
cc_84 N_8_c_93_n N_11_c_204_n 0.00137189f $X=0.434 $Y=0.2025 $X2=0.135
+ $Y2=0.2025
cc_85 N_8_c_125_p N_11_c_208_n 2.9865e-19 $X=0.593 $Y=0.234 $X2=0 $Y2=0
cc_86 N_8_c_115_n N_11_c_208_n 3.04405e-19 $X=0.824 $Y=0.036 $X2=0 $Y2=0
cc_87 N_8_c_95_n N_11_c_206_n 2.9865e-19 $X=0.45 $Y=0.234 $X2=0 $Y2=0
cc_88 N_8_c_123_p N_11_c_215_n 2.9865e-19 $X=0.5 $Y=0.234 $X2=0 $Y2=0
cc_89 N_8_c_99_n N_12_c_230_n 0.00134615f $X=0.596 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_90 N_8_c_113_n N_12_c_235_n 0.00332784f $X=0.756 $Y=0.036 $X2=0.135 $Y2=0.135
cc_91 N_8_c_115_n N_12_c_235_n 4.51951e-19 $X=0.824 $Y=0.036 $X2=0.135 $Y2=0.135
cc_92 N_8_c_113_n N_12_c_243_n 0.00360833f $X=0.756 $Y=0.036 $X2=0 $Y2=0
cc_93 N_8_c_115_n N_12_c_243_n 0.00312695f $X=0.824 $Y=0.036 $X2=0 $Y2=0
cc_94 N_8_c_134_p N_12_c_243_n 4.23807e-19 $X=0.891 $Y=0.099 $X2=0 $Y2=0
cc_95 N_8_c_125_p N_12_c_246_n 4.09962e-19 $X=0.593 $Y=0.234 $X2=0 $Y2=0
cc_96 N_8_c_102_n N_12_c_233_n 4.09962e-19 $X=0.72 $Y=0.234 $X2=0 $Y2=0
cc_97 N_8_c_137_p N_12_c_248_n 6.1248e-19 $X=0.891 $Y=0.081 $X2=0 $Y2=0
cc_98 N_8_c_113_n N_12_c_249_n 0.00126662f $X=0.756 $Y=0.036 $X2=0.081 $Y2=0.135
cc_99 N_8_c_115_n N_12_c_249_n 0.00678122f $X=0.824 $Y=0.036 $X2=0.081 $Y2=0.135
cc_100 N_8_c_111_n N_12_c_238_n 4.09962e-19 $X=0.824 $Y=0.234 $X2=0 $Y2=0
cc_101 N_8_c_113_n N_12_c_238_n 0.00112576f $X=0.756 $Y=0.036 $X2=0 $Y2=0
cc_102 N_8_c_104_n N_Y_M11_d 3.80663e-19 $X=0.999 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_103 N_8_c_104_n N_Y_M18_d 3.80663e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_104 N_8_c_104_n N_Y_c_264_n 8.00061e-19 $X=0.999 $Y=0.135 $X2=0.135 $Y2=0.135
cc_105 N_8_M11_g N_Y_c_265_n 4.59284e-19 $X=0.999 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_106 N_8_c_104_n N_Y_c_265_n 5.51214e-19 $X=0.999 $Y=0.135 $X2=0.135 $Y2=0.135
cc_107 N_8_c_147_p N_Y_c_265_n 3.9751e-19 $X=0.882 $Y=0.036 $X2=0.135 $Y2=0.135
cc_108 N_8_c_104_n N_Y_c_268_n 8.00061e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_109 N_8_M11_g N_Y_c_269_n 4.59284e-19 $X=0.999 $Y=0.0675 $X2=0 $Y2=0
cc_110 N_8_c_104_n N_Y_c_269_n 5.51214e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_111 N_8_c_151_p N_Y_c_269_n 4.03429e-19 $X=0.882 $Y=0.234 $X2=0 $Y2=0
cc_112 N_8_c_152_p Y 3.18599e-19 $X=0.891 $Y=0.189 $X2=0 $Y2=0
cc_113 N_8_c_104_n N_Y_c_273_n 5.13752e-19 $X=0.999 $Y=0.135 $X2=0 $Y2=0
cc_114 N_8_c_137_p N_Y_c_273_n 3.16757e-19 $X=0.891 $Y=0.081 $X2=0 $Y2=0
cc_115 N_9_c_160_n N_10_M2_s 3.13602e-19 $X=0.324 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_116 N_9_c_160_n N_10_c_173_n 0.00282786f $X=0.324 $Y=0.036 $X2=0.081
+ $Y2=0.135
cc_117 N_9_c_161_n N_10_c_173_n 0.0036466f $X=0.324 $Y=0.036 $X2=0.081 $Y2=0.135
cc_118 N_9_c_160_n N_10_c_191_n 4.49606e-19 $X=0.324 $Y=0.036 $X2=0.135
+ $Y2=0.135
cc_119 N_9_c_161_n N_10_c_191_n 0.0032943f $X=0.324 $Y=0.036 $X2=0.135 $Y2=0.135
cc_120 N_9_c_160_n N_10_c_184_n 0.00703507f $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_121 N_9_c_161_n N_10_c_176_n 0.00233206f $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_122 N_9_c_160_n N_11_c_206_n 3.11218e-19 $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_123 N_10_c_191_n N_11_c_204_n 0.0032943f $X=0.378 $Y=0.0675 $X2=0.351
+ $Y2=0.135
cc_124 N_10_c_178_n N_11_c_204_n 0.0036466f $X=0.484 $Y=0.0675 $X2=0.351
+ $Y2=0.135
cc_125 N_10_c_187_n N_11_c_204_n 0.00233206f $X=0.45 $Y=0.072 $X2=0.351
+ $Y2=0.135
cc_126 N_10_c_191_n N_11_c_206_n 4.49606e-19 $X=0.378 $Y=0.0675 $X2=0.297
+ $Y2=0.135
cc_127 N_10_c_178_n N_11_c_206_n 0.00315444f $X=0.484 $Y=0.0675 $X2=0.297
+ $Y2=0.135
cc_128 N_10_c_187_n N_11_c_206_n 0.00706398f $X=0.45 $Y=0.072 $X2=0.297
+ $Y2=0.135
cc_129 N_10_c_178_n N_12_c_230_n 0.00132424f $X=0.484 $Y=0.0675 $X2=0.297
+ $Y2=0.135
cc_130 N_10_c_179_n N_12_c_246_n 6.78329e-19 $X=0.486 $Y=0.072 $X2=0 $Y2=0
cc_131 N_11_c_208_n N_12_M6_s 3.13602e-19 $X=0.648 $Y=0.036 $X2=0.405 $Y2=0.0675
cc_132 N_11_c_208_n N_12_c_230_n 0.00282786f $X=0.648 $Y=0.036 $X2=0.405
+ $Y2=0.135
cc_133 N_11_c_209_n N_12_c_230_n 0.0036466f $X=0.648 $Y=0.036 $X2=0.405
+ $Y2=0.135
cc_134 N_11_c_208_n N_12_c_235_n 4.49606e-19 $X=0.648 $Y=0.036 $X2=0.459
+ $Y2=0.135
cc_135 N_11_c_209_n N_12_c_235_n 0.00340637f $X=0.648 $Y=0.036 $X2=0.459
+ $Y2=0.135
cc_136 N_11_c_208_n N_12_c_246_n 0.00703507f $X=0.648 $Y=0.036 $X2=0 $Y2=0
cc_137 N_11_c_209_n N_12_c_233_n 0.00233206f $X=0.648 $Y=0.036 $X2=0 $Y2=0

* END of "./AND5x2_ASAP7_75t_R.pex.sp.AND5X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: OR2x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:59:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OR2x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./OR2x2_ASAP7_75t_R.pex.sp.pex"
* File: OR2x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:59:18 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OR2X2_ASAP7_75T_R%B 2 5 7 18 21 26 VSS
c9 26 VSS 0.0159636f $X=0.019 $Y=0.134
c10 21 VSS 2.10262e-19 $X=0.046 $Y=0.135
c11 20 VSS 0.00102817f $X=0.04 $Y=0.135
c12 18 VSS 5.96772e-19 $X=0.063 $Y=0.135
c13 5 VSS 0.00501581f $X=0.081 $Y=0.1355
c14 2 VSS 0.0648497f $X=0.081 $Y=0.054
r15 20 21 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.135 $X2=0.046 $Y2=0.135
r16 18 21 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.135 $X2=0.046 $Y2=0.135
r17 18 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.063 $Y=0.135 $X2=0.063
+ $Y2=0.135
r18 16 26 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r19 16 20 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.04 $Y2=0.135
r20 5 19 15.6522 $w=2.3e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1355 $X2=0.063 $Y2=0.1355
r21 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1355 $X2=0.081 $Y2=0.2025
r22 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.1355
.ends

.subckt PM_OR2X2_ASAP7_75T_R%A 2 5 7 12 VSS
c19 12 VSS 0.0026637f $X=0.137 $Y=0.134
c20 5 VSS 0.00111013f $X=0.135 $Y=0.1355
c21 2 VSS 0.0589852f $X=0.135 $Y=0.054
r22 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r23 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.2025
r24 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.1355
.ends

.subckt PM_OR2X2_ASAP7_75T_R%5 2 7 10 13 15 17 18 21 22 25 32 35 36 38 43 46 47
+ 48 50 51 52 55 58 61 VSS
c36 61 VSS 2.27295e-19 $X=0.171 $Y=0.135
c37 58 VSS 1.31878e-20 $X=0.21 $Y=0.135
c38 57 VSS 7.16223e-19 $X=0.207 $Y=0.135
c39 55 VSS 9.02817e-20 $X=0.213 $Y=0.135
c40 52 VSS 5.02861e-19 $X=0.171 $Y=0.2045
c41 51 VSS 0.00112536f $X=0.171 $Y=0.184
c42 50 VSS 4.22387e-19 $X=0.171 $Y=0.225
c43 48 VSS 5.61558e-19 $X=0.171 $Y=0.086
c44 47 VSS 3.64354e-19 $X=0.171 $Y=0.063
c45 46 VSS 0.00117391f $X=0.171 $Y=0.126
c46 44 VSS 0.00147742f $X=0.153 $Y=0.036
c47 43 VSS 0.00283359f $X=0.144 $Y=0.036
c48 38 VSS 0.00216909f $X=0.108 $Y=0.036
c49 36 VSS 0.00421964f $X=0.162 $Y=0.036
c50 35 VSS 0.00314023f $X=0.144 $Y=0.234
c51 34 VSS 0.00134454f $X=0.107 $Y=0.234
c52 33 VSS 0.00172465f $X=0.094 $Y=0.234
c53 32 VSS 0.0042162f $X=0.077 $Y=0.234
c54 27 VSS 0.00603283f $X=0.162 $Y=0.234
c55 25 VSS 0.00469785f $X=0.056 $Y=0.2025
c56 22 VSS 4.64427e-19 $X=0.071 $Y=0.2025
c57 21 VSS 0.00817362f $X=0.108 $Y=0.054
c58 17 VSS 6.05457e-19 $X=0.125 $Y=0.054
c59 13 VSS 0.00499257f $X=0.243 $Y=0.135
c60 10 VSS 0.0639847f $X=0.243 $Y=0.0675
c61 2 VSS 0.0613335f $X=0.189 $Y=0.0675
r62 57 58 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.135 $X2=0.21 $Y2=0.135
r63 55 58 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.213
+ $Y=0.135 $X2=0.21 $Y2=0.135
r64 55 56 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.213 $Y=0.135 $X2=0.213
+ $Y2=0.135
r65 53 61 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.171 $Y2=0.135
r66 53 57 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.207 $Y2=0.135
r67 51 52 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.184 $X2=0.171 $Y2=0.2045
r68 50 52 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.225 $X2=0.171 $Y2=0.2045
r69 49 61 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.144 $X2=0.171 $Y2=0.135
r70 49 51 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.144 $X2=0.171 $Y2=0.184
r71 47 48 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.063 $X2=0.171 $Y2=0.086
r72 46 61 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.126 $X2=0.171 $Y2=0.135
r73 46 48 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.126 $X2=0.171 $Y2=0.086
r74 45 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.045 $X2=0.171 $Y2=0.063
r75 43 44 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.153 $Y2=0.036
r76 38 43 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.144 $Y2=0.036
r77 36 45 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.036 $X2=0.171 $Y2=0.045
r78 36 44 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.153 $Y2=0.036
r79 34 35 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.234 $X2=0.144 $Y2=0.234
r80 33 34 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.234 $X2=0.107 $Y2=0.234
r81 32 33 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.077
+ $Y=0.234 $X2=0.094 $Y2=0.234
r82 29 32 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.077 $Y2=0.234
r83 27 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.234 $X2=0.171 $Y2=0.225
r84 27 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.144 $Y2=0.234
r85 25 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r86 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r87 21 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r88 18 21 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.054 $X2=0.108 $Y2=0.054
r89 17 21 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.054 $X2=0.108 $Y2=0.054
r90 13 56 27.2727 $w=2.2e-08 $l=3e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.213 $Y2=0.135
r91 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r92 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r93 5 56 21.8182 $w=2.2e-08 $l=2.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.213 $Y2=0.135
r94 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r95 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OR2X2_ASAP7_75T_R%Y 1 2 5 6 7 10 13 18 22 24 26 28 32 34 35 36 VSS
c16 38 VSS 0.00101302f $X=0.297 $Y=0.2045
c17 36 VSS 7.93583e-20 $X=0.297 $Y=0.14575
c18 35 VSS 7.62744e-19 $X=0.297 $Y=0.144
c19 34 VSS 0.00229014f $X=0.297 $Y=0.126
c20 33 VSS 0.00176873f $X=0.297 $Y=0.086
c21 32 VSS 0.00218466f $X=0.297 $Y=0.1475
c22 30 VSS 7.5805e-19 $X=0.297 $Y=0.225
c23 28 VSS 0.00288612f $X=0.2575 $Y=0.234
c24 27 VSS 1.17723e-19 $X=0.227 $Y=0.234
c25 26 VSS 0.00201509f $X=0.225 $Y=0.234
c26 25 VSS 0.00815468f $X=0.288 $Y=0.234
c27 24 VSS 0.00288612f $X=0.2575 $Y=0.036
c28 23 VSS 1.17723e-19 $X=0.227 $Y=0.036
c29 22 VSS 0.00201509f $X=0.225 $Y=0.036
c30 21 VSS 0.00815468f $X=0.288 $Y=0.036
c31 18 VSS 9.20467e-19 $X=0.216 $Y=0.198
c32 13 VSS 9.20467e-19 $X=0.216 $Y=0.072
c33 10 VSS 0.0108958f $X=0.216 $Y=0.2025
c34 6 VSS 5.945e-19 $X=0.233 $Y=0.2025
c35 5 VSS 0.0111568f $X=0.216 $Y=0.0675
c36 1 VSS 5.945e-19 $X=0.233 $Y=0.0675
r37 37 38 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.184 $X2=0.297 $Y2=0.2045
r38 35 36 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.144 $X2=0.297 $Y2=0.14575
r39 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.144
r40 33 34 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.086 $X2=0.297 $Y2=0.126
r41 32 37 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1475 $X2=0.297 $Y2=0.184
r42 32 36 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1475 $X2=0.297 $Y2=0.14575
r43 30 38 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.225 $X2=0.297 $Y2=0.2045
r44 29 33 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.086
r45 27 28 2.07099 $w=1.8e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.227
+ $Y=0.234 $X2=0.2575 $Y2=0.234
r46 26 27 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.234 $X2=0.227 $Y2=0.234
r47 25 30 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.234 $X2=0.297 $Y2=0.225
r48 25 28 2.07099 $w=1.8e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.234 $X2=0.2575 $Y2=0.234
r49 23 24 2.07099 $w=1.8e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.227
+ $Y=0.036 $X2=0.2575 $Y2=0.036
r50 22 23 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.036 $X2=0.227 $Y2=0.036
r51 21 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r52 21 24 2.07099 $w=1.8e-08 $l=3.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.2575 $Y2=0.036
r53 16 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.225 $X2=0.225 $Y2=0.234
r54 16 18 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.225 $X2=0.216 $Y2=0.198
r55 11 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.045 $X2=0.225 $Y2=0.036
r56 11 13 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.045 $X2=0.216 $Y2=0.072
r57 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r58 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r59 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r60 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072 $X2=0.216
+ $Y2=0.072
r61 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r62 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends

.subckt PM_OR2X2_ASAP7_75T_R%7 1 2 VSS
c0 1 VSS 0.00242246f $X=0.125 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends


* END of "./OR2x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt OR2x2_ASAP7_75t_R  VSS VDD B A Y
* 
* Y	Y
* A	A
* B	B
M0 N_5_M0_d N_B_M0_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 VSS N_A_M1_g N_5_M1_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_5_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_5_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_7_M4_d N_B_M4_g N_5_M4_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 VDD N_A_M5_g N_7_M5_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M6 N_Y_M6_d N_5_M6_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M7 N_Y_M7_d N_5_M7_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
*
* 
* .include "OR2x2_ASAP7_75t_R.pex.sp.OR2X2_ASAP7_75T_R.pxi"
* BEGIN of "./OR2x2_ASAP7_75t_R.pex.sp.OR2X2_ASAP7_75T_R.pxi"
* File: OR2x2_ASAP7_75t_R.pex.sp.OR2X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:59:18 2017
* 
x_PM_OR2X2_ASAP7_75T_R%B N_B_M0_g N_B_c_2_p N_B_M4_g N_B_c_3_p N_B_c_8_p B VSS
+ PM_OR2X2_ASAP7_75T_R%B
x_PM_OR2X2_ASAP7_75T_R%A N_A_M1_g N_A_c_11_n N_A_M5_g A VSS
+ PM_OR2X2_ASAP7_75T_R%A
x_PM_OR2X2_ASAP7_75T_R%5 N_5_M2_g N_5_M6_g N_5_M3_g N_5_c_36_n N_5_M7_g N_5_M1_s
+ N_5_M0_d N_5_c_37_n N_5_M4_s N_5_c_30_n N_5_c_31_n N_5_c_39_n N_5_c_50_p
+ N_5_c_33_n N_5_c_41_n N_5_c_43_n N_5_c_53_p N_5_c_44_n N_5_c_45_n N_5_c_46_n
+ N_5_c_47_n N_5_c_63_p N_5_c_54_p N_5_c_48_n VSS PM_OR2X2_ASAP7_75T_R%5
x_PM_OR2X2_ASAP7_75T_R%Y N_Y_M3_d N_Y_M2_d N_Y_c_66_n N_Y_M7_d N_Y_M6_d
+ N_Y_c_68_n N_Y_c_69_n N_Y_c_71_n N_Y_c_73_n N_Y_c_74_n N_Y_c_75_n N_Y_c_76_n Y
+ N_Y_c_77_n N_Y_c_79_n N_Y_c_80_n VSS PM_OR2X2_ASAP7_75T_R%Y
x_PM_OR2X2_ASAP7_75T_R%7 N_7_M5_s N_7_M4_d VSS PM_OR2X2_ASAP7_75T_R%7
cc_1 N_B_M0_g N_A_M1_g 0.00344695f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_B_c_2_p N_A_c_11_n 0.00176726f $X=0.081 $Y=0.1355 $X2=0.135 $Y2=0.1355
cc_3 N_B_c_3_p A 4.06677e-19 $X=0.063 $Y=0.135 $X2=0.137 $Y2=0.134
cc_4 B A 0.00132855f $X=0.019 $Y=0.134 $X2=0.137 $Y2=0.134
cc_5 N_B_M0_g N_5_M2_g 2.31381e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_6 B N_5_c_30_n 0.00117106f $X=0.019 $Y=0.134 $X2=0 $Y2=0
cc_7 N_B_c_2_p N_5_c_31_n 3.23506e-19 $X=0.081 $Y=0.1355 $X2=0 $Y2=0
cc_8 N_B_c_8_p N_5_c_31_n 5.57559e-19 $X=0.046 $Y=0.135 $X2=0 $Y2=0
cc_9 B N_5_c_33_n 5.21568e-19 $X=0.019 $Y=0.134 $X2=0 $Y2=0
cc_10 N_A_M1_g N_5_M2_g 0.00284417f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_11 N_A_M1_g N_5_M3_g 2.31381e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_12 N_A_c_11_n N_5_c_36_n 0.00126003f $X=0.135 $Y=0.1355 $X2=0 $Y2=0
cc_13 A N_5_c_37_n 0.00183722f $X=0.137 $Y=0.134 $X2=0.046 $Y2=0.135
cc_14 A N_5_c_30_n 7.93203e-19 $X=0.137 $Y=0.134 $X2=0.018 $Y2=0.135
cc_15 N_A_M1_g N_5_c_39_n 2.38073e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_16 A N_5_c_39_n 0.00400414f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_17 N_A_M1_g N_5_c_41_n 2.34993e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_18 A N_5_c_41_n 0.00372832f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_19 A N_5_c_43_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_20 A N_5_c_44_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_21 A N_5_c_45_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_22 A N_5_c_46_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_23 A N_5_c_47_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_24 A N_5_c_48_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_25 N_5_c_36_n N_Y_M3_d 3.8044e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.054
cc_26 N_5_c_50_p N_Y_c_66_n 0.00135341f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.1355
cc_27 N_5_c_36_n N_Y_M7_d 3.8044e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_28 N_5_c_46_n N_Y_c_68_n 0.00135523f $X=0.171 $Y=0.184 $X2=0 $Y2=0
cc_29 N_5_c_53_p N_Y_c_69_n 0.00175807f $X=0.171 $Y=0.063 $X2=0 $Y2=0
cc_30 N_5_c_54_p N_Y_c_69_n 4.86094e-19 $X=0.21 $Y=0.135 $X2=0 $Y2=0
cc_31 N_5_c_47_n N_Y_c_71_n 0.00177145f $X=0.171 $Y=0.2045 $X2=0.063 $Y2=0.135
cc_32 N_5_c_54_p N_Y_c_71_n 4.86094e-19 $X=0.21 $Y=0.135 $X2=0.063 $Y2=0.135
cc_33 N_5_c_50_p N_Y_c_73_n 0.00175807f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_34 N_5_M3_g N_Y_c_74_n 2.89885e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_5_c_45_n N_Y_c_75_n 0.00177145f $X=0.171 $Y=0.225 $X2=0.019 $Y2=0.134
cc_36 N_5_M3_g N_Y_c_76_n 2.89885e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_37 N_5_c_36_n N_Y_c_77_n 4.56156e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_38 N_5_c_43_n N_Y_c_77_n 4.04965e-19 $X=0.171 $Y=0.126 $X2=0 $Y2=0
cc_39 N_5_c_63_p N_Y_c_79_n 3.74579e-19 $X=0.213 $Y=0.135 $X2=0 $Y2=0
cc_40 N_5_c_46_n N_Y_c_80_n 4.03366e-19 $X=0.171 $Y=0.184 $X2=0 $Y2=0

* END of "./OR2x2_ASAP7_75t_R.pex.sp.OR2X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: OR2x4_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:59:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OR2x4_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./OR2x4_ASAP7_75t_R.pex.sp.pex"
* File: OR2x4_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:59:41 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OR2X4_ASAP7_75T_R%B 2 5 7 18 21 26 VSS
c9 26 VSS 0.0159636f $X=0.019 $Y=0.134
c10 21 VSS 2.10262e-19 $X=0.046 $Y=0.135
c11 20 VSS 0.00102817f $X=0.04 $Y=0.135
c12 18 VSS 5.96772e-19 $X=0.063 $Y=0.135
c13 5 VSS 0.00501581f $X=0.081 $Y=0.1355
c14 2 VSS 0.0648497f $X=0.081 $Y=0.054
r15 20 21 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.135 $X2=0.046 $Y2=0.135
r16 18 21 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.135 $X2=0.046 $Y2=0.135
r17 18 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.063 $Y=0.135 $X2=0.063
+ $Y2=0.135
r18 16 26 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r19 16 20 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.04 $Y2=0.135
r20 5 19 15.6522 $w=2.3e-08 $l=1.8e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.1355 $X2=0.063 $Y2=0.1355
r21 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1355 $X2=0.081 $Y2=0.2025
r22 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.1355
.ends

.subckt PM_OR2X4_ASAP7_75T_R%A 2 5 7 12 VSS
c19 12 VSS 0.00266013f $X=0.137 $Y=0.134
c20 5 VSS 0.00111013f $X=0.135 $Y=0.1355
c21 2 VSS 0.0589852f $X=0.135 $Y=0.054
r22 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r23 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.2025
r24 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.1355
.ends

.subckt PM_OR2X4_ASAP7_75T_R%5 2 7 10 15 18 23 26 29 31 33 34 37 38 41 48 51 52
+ 54 59 62 63 64 66 67 68 74 77 VSS
c45 77 VSS 2.27295e-19 $X=0.171 $Y=0.135
c46 74 VSS 1.31878e-20 $X=0.21 $Y=0.135
c47 73 VSS 7.16223e-19 $X=0.207 $Y=0.135
c48 71 VSS 1.52796e-19 $X=0.213 $Y=0.135
c49 68 VSS 5.02861e-19 $X=0.171 $Y=0.2045
c50 67 VSS 0.00114186f $X=0.171 $Y=0.184
c51 66 VSS 4.22387e-19 $X=0.171 $Y=0.225
c52 64 VSS 5.61558e-19 $X=0.171 $Y=0.086
c53 63 VSS 3.64354e-19 $X=0.171 $Y=0.063
c54 62 VSS 0.00119042f $X=0.171 $Y=0.126
c55 60 VSS 0.00147742f $X=0.153 $Y=0.036
c56 59 VSS 0.00283359f $X=0.144 $Y=0.036
c57 54 VSS 0.00216909f $X=0.108 $Y=0.036
c58 52 VSS 0.00421964f $X=0.162 $Y=0.036
c59 51 VSS 0.00314023f $X=0.144 $Y=0.234
c60 50 VSS 0.00134454f $X=0.107 $Y=0.234
c61 49 VSS 0.00172465f $X=0.094 $Y=0.234
c62 48 VSS 0.0042162f $X=0.077 $Y=0.234
c63 43 VSS 0.00603283f $X=0.162 $Y=0.234
c64 41 VSS 0.00469785f $X=0.056 $Y=0.2025
c65 38 VSS 4.64427e-19 $X=0.071 $Y=0.2025
c66 37 VSS 0.00817362f $X=0.108 $Y=0.054
c67 33 VSS 6.05457e-19 $X=0.125 $Y=0.054
c68 29 VSS 0.0158073f $X=0.351 $Y=0.135
c69 26 VSS 0.0639847f $X=0.351 $Y=0.0675
c70 18 VSS 0.0638949f $X=0.297 $Y=0.0675
c71 10 VSS 0.0636879f $X=0.243 $Y=0.0675
c72 2 VSS 0.0611266f $X=0.189 $Y=0.0675
r73 73 74 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.135 $X2=0.21 $Y2=0.135
r74 71 74 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.213
+ $Y=0.135 $X2=0.21 $Y2=0.135
r75 71 72 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.213 $Y=0.135 $X2=0.213
+ $Y2=0.135
r76 69 77 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.171 $Y2=0.135
r77 69 73 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.207 $Y2=0.135
r78 67 68 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.184 $X2=0.171 $Y2=0.2045
r79 66 68 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.225 $X2=0.171 $Y2=0.2045
r80 65 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.144 $X2=0.171 $Y2=0.135
r81 65 67 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.144 $X2=0.171 $Y2=0.184
r82 63 64 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.063 $X2=0.171 $Y2=0.086
r83 62 77 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.126 $X2=0.171 $Y2=0.135
r84 62 64 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.126 $X2=0.171 $Y2=0.086
r85 61 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.045 $X2=0.171 $Y2=0.063
r86 59 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.153 $Y2=0.036
r87 54 59 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.144 $Y2=0.036
r88 52 61 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.036 $X2=0.171 $Y2=0.045
r89 52 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.153 $Y2=0.036
r90 50 51 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.234 $X2=0.144 $Y2=0.234
r91 49 50 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.234 $X2=0.107 $Y2=0.234
r92 48 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.077
+ $Y=0.234 $X2=0.094 $Y2=0.234
r93 45 48 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.077 $Y2=0.234
r94 43 66 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.234 $X2=0.171 $Y2=0.225
r95 43 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.144 $Y2=0.234
r96 41 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r97 38 41 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r98 37 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r99 34 37 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.054 $X2=0.108 $Y2=0.054
r100 33 37 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.054 $X2=0.108 $Y2=0.054
r101 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r102 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r103 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r104 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.135 $X2=0.297 $Y2=0.2025
r105 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.0675 $X2=0.297 $Y2=0.135
r106 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.297 $Y2=0.135
r107 13 72 27.2727 $w=2.2e-08 $l=3e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.213 $Y2=0.135
r108 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.135 $X2=0.243 $Y2=0.2025
r109 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.243 $Y=0.0675 $X2=0.243 $Y2=0.135
r110 5 72 21.8182 $w=2.2e-08 $l=2.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.213 $Y2=0.135
r111 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r112 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OR2X4_ASAP7_75T_R%Y 1 2 5 6 7 10 11 12 15 16 17 20 23 28 31 32 34 35
+ 36 38 41 46 49 51 56 58 VSS
c25 64 VSS 0.00150149f $X=0.324 $Y=0.234
c26 63 VSS 0.00150149f $X=0.324 $Y=0.036
c27 62 VSS 0.00101302f $X=0.405 $Y=0.2045
c28 60 VSS 7.51787e-20 $X=0.405 $Y=0.14575
c29 59 VSS 8.65162e-19 $X=0.405 $Y=0.144
c30 58 VSS 0.00285296f $X=0.405 $Y=0.126
c31 57 VSS 0.00176873f $X=0.405 $Y=0.086
c32 56 VSS 0.00274913f $X=0.407 $Y=0.1475
c33 54 VSS 7.5805e-19 $X=0.405 $Y=0.225
c34 51 VSS 0.0112873f $X=0.396 $Y=0.234
c35 49 VSS 0.0112873f $X=0.396 $Y=0.036
c36 46 VSS 0.00117559f $X=0.324 $Y=0.198
c37 41 VSS 0.00117559f $X=0.324 $Y=0.072
c38 38 VSS 0.00528351f $X=0.271 $Y=0.234
c39 37 VSS 1.17723e-19 $X=0.227 $Y=0.234
c40 36 VSS 0.0020097f $X=0.225 $Y=0.234
c41 35 VSS 0.00508372f $X=0.315 $Y=0.234
c42 34 VSS 0.00528351f $X=0.271 $Y=0.036
c43 33 VSS 1.17723e-19 $X=0.227 $Y=0.036
c44 32 VSS 0.0020097f $X=0.225 $Y=0.036
c45 31 VSS 0.00508372f $X=0.315 $Y=0.036
c46 28 VSS 5.20536e-19 $X=0.216 $Y=0.198
c47 23 VSS 5.20536e-19 $X=0.216 $Y=0.072
c48 20 VSS 0.0105054f $X=0.324 $Y=0.2025
c49 16 VSS 5.38922e-19 $X=0.341 $Y=0.2025
c50 15 VSS 0.0108809f $X=0.216 $Y=0.2025
c51 11 VSS 5.945e-19 $X=0.233 $Y=0.2025
c52 10 VSS 0.0105054f $X=0.324 $Y=0.0675
c53 6 VSS 5.38922e-19 $X=0.341 $Y=0.0675
c54 5 VSS 0.0111419f $X=0.216 $Y=0.0675
c55 1 VSS 5.945e-19 $X=0.233 $Y=0.0675
r56 61 62 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.184 $X2=0.405 $Y2=0.2045
r57 59 60 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.144 $X2=0.405 $Y2=0.14575
r58 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.126 $X2=0.405 $Y2=0.144
r59 57 58 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.086 $X2=0.405 $Y2=0.126
r60 56 61 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.1475 $X2=0.405 $Y2=0.184
r61 56 60 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.1475 $X2=0.405 $Y2=0.14575
r62 54 62 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.2045
r63 53 57 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.086
r64 52 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.234 $X2=0.324 $Y2=0.234
r65 51 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r66 51 52 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.333 $Y2=0.234
r67 50 63 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.036 $X2=0.324 $Y2=0.036
r68 49 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r69 49 50 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.333 $Y2=0.036
r70 44 64 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.225 $X2=0.324 $Y2=0.234
r71 44 46 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.225 $X2=0.324 $Y2=0.198
r72 39 63 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.045 $X2=0.324 $Y2=0.036
r73 39 41 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.045 $X2=0.324 $Y2=0.072
r74 37 38 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.227
+ $Y=0.234 $X2=0.271 $Y2=0.234
r75 36 37 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.234 $X2=0.227 $Y2=0.234
r76 35 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.315
+ $Y=0.234 $X2=0.324 $Y2=0.234
r77 35 38 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.315
+ $Y=0.234 $X2=0.271 $Y2=0.234
r78 33 34 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.227
+ $Y=0.036 $X2=0.271 $Y2=0.036
r79 32 33 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.036 $X2=0.227 $Y2=0.036
r80 31 63 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.315
+ $Y=0.036 $X2=0.324 $Y2=0.036
r81 31 34 2.98765 $w=1.8e-08 $l=4.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.315
+ $Y=0.036 $X2=0.271 $Y2=0.036
r82 26 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.225 $X2=0.225 $Y2=0.234
r83 26 28 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.225 $X2=0.216 $Y2=0.198
r84 21 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.045 $X2=0.225 $Y2=0.036
r85 21 23 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.045 $X2=0.216 $Y2=0.072
r86 20 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.198 $X2=0.324
+ $Y2=0.198
r87 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r88 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r89 15 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198 $X2=0.216
+ $Y2=0.198
r90 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r91 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r92 10 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.072 $X2=0.324
+ $Y2=0.072
r93 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r94 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r95 5 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.072 $X2=0.216
+ $Y2=0.072
r96 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.199
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
r97 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.216 $Y2=0.0675
.ends

.subckt PM_OR2X4_ASAP7_75T_R%7 1 2 VSS
c0 1 VSS 0.00242246f $X=0.125 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends


* END of "./OR2x4_ASAP7_75t_R.pex.sp.pex"
* 
.subckt OR2x4_ASAP7_75t_R  VSS VDD B A Y
* 
* Y	Y
* A	A
* B	B
M0 N_5_M0_d N_B_M0_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 VSS N_A_M1_g N_5_M1_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_5_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_5_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_5_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_5_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_7_M6_d N_B_M6_g N_5_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 VDD N_A_M7_g N_7_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M8 N_Y_M8_d N_5_M8_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M9 N_Y_M9_d N_5_M9_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M10 N_Y_M10_d N_5_M10_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_Y_M11_d N_5_M11_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "OR2x4_ASAP7_75t_R.pex.sp.OR2X4_ASAP7_75T_R.pxi"
* BEGIN of "./OR2x4_ASAP7_75t_R.pex.sp.OR2X4_ASAP7_75T_R.pxi"
* File: OR2x4_ASAP7_75t_R.pex.sp.OR2X4_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:59:41 2017
* 
x_PM_OR2X4_ASAP7_75T_R%B N_B_M0_g N_B_c_2_p N_B_M6_g N_B_c_3_p N_B_c_8_p B VSS
+ PM_OR2X4_ASAP7_75T_R%B
x_PM_OR2X4_ASAP7_75T_R%A N_A_M1_g N_A_c_11_n N_A_M7_g A VSS
+ PM_OR2X4_ASAP7_75T_R%A
x_PM_OR2X4_ASAP7_75T_R%5 N_5_M2_g N_5_M8_g N_5_M3_g N_5_M9_g N_5_M4_g N_5_M10_g
+ N_5_M5_g N_5_c_36_n N_5_M11_g N_5_M1_s N_5_M0_d N_5_c_37_n N_5_M6_s N_5_c_30_n
+ N_5_c_31_n N_5_c_39_n N_5_c_50_p N_5_c_33_n N_5_c_41_n N_5_c_43_n N_5_c_57_p
+ N_5_c_44_n N_5_c_45_n N_5_c_46_n N_5_c_47_n N_5_c_58_p N_5_c_48_n VSS
+ PM_OR2X4_ASAP7_75T_R%5
x_PM_OR2X4_ASAP7_75T_R%Y N_Y_M3_d N_Y_M2_d N_Y_c_75_n N_Y_M5_d N_Y_M4_d
+ N_Y_c_77_n N_Y_M9_d N_Y_M8_d N_Y_c_79_n N_Y_M11_d N_Y_M10_d N_Y_c_81_n
+ N_Y_c_82_n N_Y_c_84_n N_Y_c_86_n N_Y_c_87_n N_Y_c_88_n N_Y_c_90_n N_Y_c_91_n
+ N_Y_c_92_n N_Y_c_94_n N_Y_c_95_n N_Y_c_96_n N_Y_c_97_n Y N_Y_c_98_n VSS
+ PM_OR2X4_ASAP7_75T_R%Y
x_PM_OR2X4_ASAP7_75T_R%7 N_7_M7_s N_7_M6_d VSS PM_OR2X4_ASAP7_75T_R%7
cc_1 N_B_M0_g N_A_M1_g 0.00344695f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_B_c_2_p N_A_c_11_n 0.00176726f $X=0.081 $Y=0.1355 $X2=0.135 $Y2=0.1355
cc_3 N_B_c_3_p A 4.06677e-19 $X=0.063 $Y=0.135 $X2=0.137 $Y2=0.134
cc_4 B A 0.00132855f $X=0.019 $Y=0.134 $X2=0.137 $Y2=0.134
cc_5 N_B_M0_g N_5_M2_g 2.31381e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_6 B N_5_c_30_n 0.00117106f $X=0.019 $Y=0.134 $X2=0 $Y2=0
cc_7 N_B_c_2_p N_5_c_31_n 3.23506e-19 $X=0.081 $Y=0.1355 $X2=0 $Y2=0
cc_8 N_B_c_8_p N_5_c_31_n 5.57559e-19 $X=0.046 $Y=0.135 $X2=0 $Y2=0
cc_9 B N_5_c_33_n 5.21568e-19 $X=0.019 $Y=0.134 $X2=0 $Y2=0
cc_10 N_A_M1_g N_5_M2_g 0.00284417f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_11 N_A_M1_g N_5_M3_g 2.31381e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_12 N_A_c_11_n N_5_c_36_n 0.00125168f $X=0.135 $Y=0.1355 $X2=0.081 $Y2=0.1355
cc_13 A N_5_c_37_n 0.00183722f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_14 A N_5_c_30_n 7.93203e-19 $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_15 N_A_M1_g N_5_c_39_n 2.38073e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_16 A N_5_c_39_n 0.00400414f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_17 N_A_M1_g N_5_c_41_n 2.34993e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_18 A N_5_c_41_n 0.00372832f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_19 A N_5_c_43_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_20 A N_5_c_44_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_21 A N_5_c_45_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_22 A N_5_c_46_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_23 A N_5_c_47_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_24 A N_5_c_48_n 0.00197581f $X=0.137 $Y=0.134 $X2=0 $Y2=0
cc_25 N_5_c_36_n N_Y_M3_d 3.8044e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.054
cc_26 N_5_c_50_p N_Y_c_75_n 0.00112671f $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.1355
cc_27 N_5_c_36_n N_Y_M5_d 3.80663e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_28 N_5_c_36_n N_Y_c_77_n 8.00061e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_29 N_5_c_36_n N_Y_M9_d 3.8044e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_30 N_5_c_46_n N_Y_c_79_n 0.00112854f $X=0.171 $Y=0.184 $X2=0 $Y2=0
cc_31 N_5_c_36_n N_Y_M11_d 3.80663e-19 $X=0.351 $Y=0.135 $X2=0.027 $Y2=0.135
cc_32 N_5_c_36_n N_Y_c_81_n 8.00061e-19 $X=0.351 $Y=0.135 $X2=0.04 $Y2=0.135
cc_33 N_5_c_57_p N_Y_c_82_n 0.00177252f $X=0.171 $Y=0.063 $X2=0 $Y2=0
cc_34 N_5_c_58_p N_Y_c_82_n 4.86094e-19 $X=0.21 $Y=0.135 $X2=0 $Y2=0
cc_35 N_5_c_47_n N_Y_c_84_n 0.00179083f $X=0.171 $Y=0.2045 $X2=0 $Y2=0
cc_36 N_5_c_58_p N_Y_c_84_n 4.86094e-19 $X=0.21 $Y=0.135 $X2=0 $Y2=0
cc_37 N_5_M4_g N_Y_c_86_n 2.89885e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_38 N_5_c_50_p N_Y_c_87_n 0.00177252f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_39 N_5_M3_g N_Y_c_88_n 2.89885e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_40 N_5_c_36_n N_Y_c_88_n 7.93486e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_41 N_5_M4_g N_Y_c_90_n 2.89885e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_42 N_5_c_45_n N_Y_c_91_n 0.00179083f $X=0.171 $Y=0.225 $X2=0 $Y2=0
cc_43 N_5_M3_g N_Y_c_92_n 2.89885e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_5_c_36_n N_Y_c_92_n 7.93486e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_45 N_5_c_36_n N_Y_c_94_n 2.47493e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_46 N_5_c_36_n N_Y_c_95_n 2.47493e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_47 N_5_M5_g N_Y_c_96_n 2.89885e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_48 N_5_M5_g N_Y_c_97_n 2.89885e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_49 N_5_c_36_n N_Y_c_98_n 9.13063e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0

* END of "./OR2x4_ASAP7_75t_R.pex.sp.OR2X4_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: OR2x6_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:00:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OR2x6_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./OR2x6_ASAP7_75t_R.pex.sp.pex"
* File: OR2x6_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:00:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OR2X6_ASAP7_75T_R%B 2 5 7 10 13 15 24 25 26 27 28 30 35 42 49 VSS
c32 49 VSS 0.00148483f $X=0.243 $Y=0.1575
c33 47 VSS 3.08436e-19 $X=0.243 $Y=0.162
c34 42 VSS 3.41081e-19 $X=0.243 $Y=0.135
c35 35 VSS 0.00726985f $X=0.081 $Y=0.162
c36 30 VSS 3.05217e-19 $X=0.081 $Y=0.135
c37 28 VSS 1.5262e-19 $X=0.148 $Y=0.162
c38 27 VSS 3.20044e-19 $X=0.144 $Y=0.162
c39 26 VSS 6.79482e-19 $X=0.126 $Y=0.162
c40 25 VSS 1.33656e-19 $X=0.109 $Y=0.162
c41 13 VSS 0.00149016f $X=0.243 $Y=0.135
c42 10 VSS 0.059021f $X=0.243 $Y=0.054
c43 5 VSS 0.00213343f $X=0.081 $Y=0.135
c44 2 VSS 0.0630726f $X=0.081 $Y=0.054
r45 48 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.153 $X2=0.243 $Y2=0.1575
r46 47 49 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.162 $X2=0.243 $Y2=0.1575
r47 42 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.153
r48 36 37 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.153 $X2=0.081 $Y2=0.1575
r49 35 37 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.162 $X2=0.081 $Y2=0.1575
r50 30 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.153
r51 27 28 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.162 $X2=0.148 $Y2=0.162
r52 26 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.162 $X2=0.144 $Y2=0.162
r53 25 26 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.162 $X2=0.126 $Y2=0.162
r54 24 28 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.172
+ $Y=0.162 $X2=0.148 $Y2=0.162
r55 22 35 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.162 $X2=0.081 $Y2=0.162
r56 22 25 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.162 $X2=0.109 $Y2=0.162
r57 21 47 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.162 $X2=0.243 $Y2=0.162
r58 21 24 4.20988 $w=1.8e-08 $l=6.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.162 $X2=0.172 $Y2=0.162
r59 13 42 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r60 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r61 10 13 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.135
r62 5 30 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r63 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r64 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OR2X6_ASAP7_75T_R%A 2 7 10 13 15 17 19 20 23 24 25 28 VSS
c22 31 VSS 1.91948e-19 $X=0.135 $Y=0.098
c23 30 VSS 1.95531e-19 $X=0.135 $Y=0.088
c24 28 VSS 3.70061e-19 $X=0.135 $Y=0.108
c25 25 VSS 2.70577e-20 $X=0.11 $Y=0.072
c26 24 VSS 1.62967e-19 $X=0.094 $Y=0.072
c27 23 VSS 5.31938e-19 $X=0.09 $Y=0.072
c28 22 VSS 0.00592527f $X=0.072 $Y=0.072
c29 21 VSS 0.0017909f $X=0.027 $Y=0.072
c30 20 VSS 0.00101993f $X=0.126 $Y=0.072
c31 17 VSS 0.00896867f $X=0.018 $Y=0.081
c32 13 VSS 0.00723545f $X=0.189 $Y=0.108
c33 10 VSS 0.0621765f $X=0.189 $Y=0.054
c34 2 VSS 0.0622716f $X=0.135 $Y=0.054
r35 30 31 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.088 $X2=0.135 $Y2=0.098
r36 28 31 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.108 $X2=0.135 $Y2=0.098
r37 26 30 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.081 $X2=0.135 $Y2=0.088
r38 24 25 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.072 $X2=0.11 $Y2=0.072
r39 23 24 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.094 $Y2=0.072
r40 22 23 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.072 $X2=0.09 $Y2=0.072
r41 21 22 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.072 $X2=0.072 $Y2=0.072
r42 20 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.126 $Y=0.072 $X2=0.135 $Y2=0.081
r43 20 25 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.11 $Y2=0.072
r44 17 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.081 $X2=0.027 $Y2=0.072
r45 17 19 3.59877 $w=1.8e-08 $l=5.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.081 $X2=0.018 $Y2=0.134
r46 13 15 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.108 $X2=0.189 $Y2=0.2025
r47 10 13 202.311 $w=2e-08 $l=5.4e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.108
r48 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.108 $X2=0.189 $Y2=0.108
r49 5 28 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.108 $X2=0.135
+ $Y2=0.108
r50 5 7 354.044 $w=2e-08 $l=9.45e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.108 $X2=0.135 $Y2=0.2025
r51 2 5 202.311 $w=2e-08 $l=5.4e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.108
.ends

.subckt PM_OR2X6_ASAP7_75T_R%5 2 7 10 15 18 23 26 31 34 39 42 45 47 49 50 53 54
+ 55 59 60 63 64 72 73 74 79 85 86 90 93 VSS
c55 93 VSS 2.02535e-19 $X=0.297 $Y=0.128
c56 92 VSS 6.23903e-19 $X=0.297 $Y=0.121
c57 90 VSS 7.13603e-19 $X=0.297 $Y=0.135
c58 86 VSS 5.57048e-20 $X=0.252 $Y=0.079
c59 85 VSS 0.00391688f $X=0.288 $Y=0.079
c60 84 VSS 3.30458e-19 $X=0.243 $Y=0.0665
c61 83 VSS 8.65169e-19 $X=0.243 $Y=0.063
c62 82 VSS 3.0506e-19 $X=0.243 $Y=0.07
c63 80 VSS 0.00229019f $X=0.27 $Y=0.198
c64 79 VSS 0.00352732f $X=0.252 $Y=0.198
c65 74 VSS 0.00158614f $X=0.288 $Y=0.198
c66 73 VSS 0.00532351f $X=0.18 $Y=0.036
c67 72 VSS 0.00511986f $X=0.144 $Y=0.036
c68 64 VSS 0.00792543f $X=0.234 $Y=0.036
c69 63 VSS 0.00440707f $X=0.162 $Y=0.2025
c70 59 VSS 7.89519e-19 $X=0.179 $Y=0.2025
c71 58 VSS 0.00873399f $X=0.216 $Y=0.054
c72 54 VSS 5.3314e-19 $X=0.233 $Y=0.054
c73 53 VSS 0.00873066f $X=0.108 $Y=0.054
c74 49 VSS 6.87793e-19 $X=0.125 $Y=0.054
c75 45 VSS 0.0246939f $X=0.567 $Y=0.135
c76 42 VSS 0.0645347f $X=0.567 $Y=0.0675
c77 34 VSS 0.0644226f $X=0.513 $Y=0.0675
c78 26 VSS 0.0642127f $X=0.459 $Y=0.0675
c79 18 VSS 0.0640423f $X=0.405 $Y=0.0675
c80 10 VSS 0.0640423f $X=0.351 $Y=0.0675
c81 2 VSS 0.0601423f $X=0.297 $Y=0.0675
r82 94 95 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.171 $X2=0.297 $Y2=0.18
r83 92 93 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.121 $X2=0.297 $Y2=0.128
r84 90 94 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.171
r85 90 93 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.128
r86 88 95 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.189 $X2=0.297 $Y2=0.18
r87 87 92 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.088 $X2=0.297 $Y2=0.121
r88 85 87 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.079 $X2=0.297 $Y2=0.088
r89 85 86 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.079 $X2=0.252 $Y2=0.079
r90 83 84 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.063 $X2=0.243 $Y2=0.0665
r91 82 86 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.243 $Y=0.07 $X2=0.252 $Y2=0.079
r92 82 84 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.07 $X2=0.243 $Y2=0.0665
r93 81 83 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.045 $X2=0.243 $Y2=0.063
r94 79 80 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.27 $Y2=0.198
r95 76 79 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.198 $X2=0.252 $Y2=0.198
r96 74 88 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.198 $X2=0.297 $Y2=0.189
r97 74 80 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.27 $Y2=0.198
r98 72 73 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.18 $Y2=0.036
r99 70 73 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.18 $Y2=0.036
r100 66 72 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.144 $Y2=0.036
r101 64 81 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.234 $Y=0.036 $X2=0.243 $Y2=0.045
r102 64 70 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.216 $Y2=0.036
r103 63 76 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.198
+ $X2=0.162 $Y2=0.198
r104 60 63 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.162 $Y2=0.2025
r105 59 63 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.2025 $X2=0.162 $Y2=0.2025
r106 58 70 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r107 55 58 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.054 $X2=0.216 $Y2=0.054
r108 54 58 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.054 $X2=0.216 $Y2=0.054
r109 53 66 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r110 50 53 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.054 $X2=0.108 $Y2=0.054
r111 49 53 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.054 $X2=0.108 $Y2=0.054
r112 45 47 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.135 $X2=0.567 $Y2=0.2025
r113 42 45 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.567 $Y=0.0675 $X2=0.567 $Y2=0.135
r114 37 45 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.567 $Y2=0.135
r115 37 39 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r116 34 37 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r117 29 37 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.513 $Y2=0.135
r118 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r119 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r120 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r121 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r122 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r123 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r124 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r125 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r126 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r127 5 90 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r128 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r129 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OR2X6_ASAP7_75T_R%Y 1 2 6 7 11 12 16 17 20 21 22 25 26 27 30 31 33 44
+ 47 51 54 58 VSS
c30 62 VSS 4.55454e-19 $X=0.621 $Y=0.216
c31 60 VSS 0.00270058f $X=0.621 $Y=0.10875
c32 59 VSS 0.00131846f $X=0.621 $Y=0.07
c33 58 VSS 0.00635587f $X=0.6215 $Y=0.1475
c34 56 VSS 4.30151e-19 $X=0.621 $Y=0.225
c35 54 VSS 0.00929752f $X=0.54 $Y=0.036
c36 51 VSS 0.00928909f $X=0.432 $Y=0.036
c37 47 VSS 0.0101927f $X=0.324 $Y=0.036
c38 44 VSS 0.0384823f $X=0.612 $Y=0.036
c39 33 VSS 0.00332891f $X=0.324 $Y=0.234
c40 31 VSS 0.0376498f $X=0.612 $Y=0.234
c41 30 VSS 0.00929752f $X=0.54 $Y=0.2025
c42 26 VSS 5.38922e-19 $X=0.557 $Y=0.2025
c43 25 VSS 0.00928903f $X=0.432 $Y=0.2025
c44 21 VSS 5.38922e-19 $X=0.449 $Y=0.2025
c45 20 VSS 0.0104341f $X=0.324 $Y=0.2025
c46 16 VSS 5.25448e-19 $X=0.341 $Y=0.2025
c47 11 VSS 5.38922e-19 $X=0.557 $Y=0.0675
c48 6 VSS 5.38922e-19 $X=0.449 $Y=0.0675
c49 1 VSS 5.72268e-19 $X=0.341 $Y=0.0675
r50 61 62 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.207 $X2=0.621 $Y2=0.216
r51 59 60 2.63117 $w=1.8e-08 $l=3.875e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.07 $X2=0.621 $Y2=0.10875
r52 58 61 4.04012 $w=1.8e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.1475 $X2=0.621 $Y2=0.207
r53 58 60 2.63117 $w=1.8e-08 $l=3.875e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.1475 $X2=0.621 $Y2=0.10875
r54 56 62 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.225 $X2=0.621 $Y2=0.216
r55 55 59 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.045 $X2=0.621 $Y2=0.07
r56 53 54 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r57 50 53 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.54 $Y2=0.036
r58 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r59 46 50 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.432 $Y2=0.036
r60 46 47 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r61 44 55 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.036 $X2=0.621 $Y2=0.045
r62 44 53 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.54 $Y2=0.036
r63 39 42 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.54 $Y2=0.234
r64 33 39 7.33333 $w=1.8e-08 $l=1.08e-07 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.432 $Y2=0.234
r65 31 56 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.612 $Y=0.234 $X2=0.621 $Y2=0.225
r66 31 42 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.234 $X2=0.54 $Y2=0.234
r67 30 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r68 27 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.2025 $X2=0.54 $Y2=0.2025
r69 26 30 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.2025 $X2=0.54 $Y2=0.2025
r70 25 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r71 22 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r72 21 25 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r73 20 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r74 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.324 $Y2=0.2025
r75 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.324 $Y2=0.2025
r76 15 54 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r77 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.523 $Y=0.0675 $X2=0.54 $Y2=0.0675
r78 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.557 $Y=0.0675 $X2=0.54 $Y2=0.0675
r79 10 51 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r80 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r81 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r82 5 47 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r83 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.324 $Y2=0.0675
r84 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.0675 $X2=0.324 $Y2=0.0675
.ends

.subckt PM_OR2X6_ASAP7_75T_R%7 1 2 VSS
c3 1 VSS 0.00207522f $X=0.125 $Y=0.2025
r4 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends

.subckt PM_OR2X6_ASAP7_75T_R%8 1 2 VSS
c2 1 VSS 0.00227757f $X=0.233 $Y=0.2025
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.199 $Y2=0.2025
.ends


* END of "./OR2x6_ASAP7_75t_R.pex.sp.pex"
* 
.subckt OR2x6_ASAP7_75t_R  VSS VDD B A Y
* 
* Y	Y
* A	A
* B	B
M0 N_5_M0_d N_B_M0_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 VSS N_A_M1_g N_5_M1_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_A_M2_g N_5_M2_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 N_5_M3_d N_B_M3_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_5_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_5_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_5_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_5_M7_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_Y_M8_d N_5_M8_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M9 N_Y_M9_d N_5_M9_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M10 VDD N_B_M10_g N_7_M10_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M11 N_7_M11_d N_A_M11_g N_5_M11_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M12 N_8_M12_d N_A_M12_g N_5_M12_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M13 VDD N_B_M13_g N_8_M13_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M14 N_Y_M14_d N_5_M14_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M15 N_Y_M15_d N_5_M15_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M16 N_Y_M16_d N_5_M16_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M17 N_Y_M17_d N_5_M17_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M18 N_Y_M18_d N_5_M18_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M19 N_Y_M19_d N_5_M19_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
*
* 
* .include "OR2x6_ASAP7_75t_R.pex.sp.OR2X6_ASAP7_75T_R.pxi"
* BEGIN of "./OR2x6_ASAP7_75t_R.pex.sp.OR2X6_ASAP7_75T_R.pxi"
* File: OR2x6_ASAP7_75t_R.pex.sp.OR2X6_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:00:03 2017
* 
x_PM_OR2X6_ASAP7_75T_R%B N_B_M0_g N_B_c_8_p N_B_M10_g N_B_M3_g N_B_c_16_p
+ N_B_M13_g B N_B_c_12_p N_B_c_30_p N_B_c_3_p N_B_c_7_p N_B_c_9_p N_B_c_18_p
+ N_B_c_26_p N_B_c_6_p VSS PM_OR2X6_ASAP7_75T_R%B
x_PM_OR2X6_ASAP7_75T_R%A N_A_M1_g N_A_M11_g N_A_M2_g N_A_c_39_n N_A_M12_g
+ N_A_c_40_n A N_A_c_47_p N_A_c_42_n N_A_c_44_n N_A_c_48_p N_A_c_45_n VSS
+ PM_OR2X6_ASAP7_75T_R%A
x_PM_OR2X6_ASAP7_75T_R%5 N_5_M4_g N_5_M14_g N_5_M5_g N_5_M15_g N_5_M6_g
+ N_5_M16_g N_5_M7_g N_5_M17_g N_5_M8_g N_5_M18_g N_5_M9_g N_5_c_57_n N_5_M19_g
+ N_5_M1_s N_5_M0_d N_5_c_58_n N_5_M3_d N_5_M2_s N_5_M12_s N_5_M11_s N_5_c_59_n
+ N_5_c_61_n N_5_c_75_n N_5_c_62_n N_5_c_96_p N_5_c_63_n N_5_c_105_p N_5_c_66_n
+ N_5_c_68_n N_5_c_69_n VSS PM_OR2X6_ASAP7_75T_R%5
x_PM_OR2X6_ASAP7_75T_R%Y N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M6_d N_Y_M9_d N_Y_M8_d
+ N_Y_M15_d N_Y_M14_d N_Y_c_114_n N_Y_M17_d N_Y_M16_d N_Y_c_117_n N_Y_M19_d
+ N_Y_M18_d N_Y_c_119_n N_Y_c_120_n N_Y_c_125_n N_Y_c_128_n N_Y_c_135_n
+ N_Y_c_137_n N_Y_c_138_n Y VSS PM_OR2X6_ASAP7_75T_R%Y
x_PM_OR2X6_ASAP7_75T_R%7 N_7_M11_d N_7_M10_s VSS PM_OR2X6_ASAP7_75T_R%7
x_PM_OR2X6_ASAP7_75T_R%8 N_8_M13_s N_8_M12_d VSS PM_OR2X6_ASAP7_75T_R%8
cc_1 N_B_M0_g N_A_M1_g 0.00344695f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_B_M3_g N_A_M1_g 2.66145e-19 $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_3 N_B_c_3_p N_A_M1_g 4.46756e-19 $X=0.144 $Y=0.162 $X2=0.135 $Y2=0.054
cc_4 N_B_M0_g N_A_M2_g 2.66145e-19 $X=0.081 $Y=0.054 $X2=0.189 $Y2=0.054
cc_5 N_B_M3_g N_A_M2_g 0.00344695f $X=0.243 $Y=0.054 $X2=0.189 $Y2=0.054
cc_6 N_B_c_6_p N_A_M2_g 3.81735e-19 $X=0.243 $Y=0.1575 $X2=0.189 $Y2=0.054
cc_7 N_B_c_7_p N_A_c_39_n 8.53719e-19 $X=0.148 $Y=0.162 $X2=0.189 $Y2=0.108
cc_8 N_B_c_8_p N_A_c_40_n 2.70475e-19 $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.081
cc_9 N_B_c_9_p N_A_c_40_n 0.00331833f $X=0.081 $Y=0.135 $X2=0.018 $Y2=0.081
cc_10 N_B_M0_g N_A_c_42_n 3.94529e-19 $X=0.081 $Y=0.054 $X2=0.09 $Y2=0.072
cc_11 N_B_c_9_p N_A_c_42_n 7.91413e-19 $X=0.081 $Y=0.135 $X2=0.09 $Y2=0.072
cc_12 N_B_c_12_p N_A_c_44_n 3.98522e-19 $X=0.109 $Y=0.162 $X2=0.094 $Y2=0.072
cc_13 N_B_c_3_p N_A_c_45_n 9.68728e-19 $X=0.144 $Y=0.162 $X2=0.135 $Y2=0.108
cc_14 N_B_M3_g N_5_M4_g 0.00284417f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_15 N_B_M3_g N_5_M5_g 2.31381e-19 $X=0.243 $Y=0.054 $X2=0.189 $Y2=0.054
cc_16 N_B_c_16_p N_5_c_57_n 9.68814e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_17 N_B_c_12_p N_5_c_58_n 2.36853e-19 $X=0.109 $Y=0.162 $X2=0 $Y2=0
cc_18 N_B_c_18_p N_5_c_59_n 0.00101747f $X=0.081 $Y=0.162 $X2=0 $Y2=0
cc_19 N_B_c_6_p N_5_c_59_n 0.002123f $X=0.243 $Y=0.1575 $X2=0 $Y2=0
cc_20 N_B_c_7_p N_5_c_61_n 6.58693e-19 $X=0.148 $Y=0.162 $X2=0 $Y2=0
cc_21 N_B_c_12_p N_5_c_62_n 6.58693e-19 $X=0.109 $Y=0.162 $X2=0 $Y2=0
cc_22 N_B_M3_g N_5_c_63_n 3.37536e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_23 N_B_c_18_p N_5_c_63_n 5.57985e-19 $X=0.081 $Y=0.162 $X2=0 $Y2=0
cc_24 N_B_c_6_p N_5_c_63_n 0.00885372f $X=0.243 $Y=0.1575 $X2=0 $Y2=0
cc_25 N_B_M3_g N_5_c_66_n 2.23918e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_26 N_B_c_26_p N_5_c_66_n 9.91574e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_27 N_B_c_26_p N_5_c_68_n 0.00109779f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_28 N_B_c_26_p N_5_c_69_n 0.00109779f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_29 N_B_c_12_p N_7_M11_d 3.00753e-19 $X=0.109 $Y=0.162 $X2=0.135 $Y2=0.054
cc_30 N_B_c_30_p N_7_M11_d 2.63708e-19 $X=0.126 $Y=0.162 $X2=0.135 $Y2=0.054
cc_31 N_B_c_18_p N_7_M11_d 2.89529e-19 $X=0.081 $Y=0.162 $X2=0.135 $Y2=0.054
cc_32 N_B_c_6_p N_8_M13_s 4.94723e-19 $X=0.243 $Y=0.1575 $X2=0.135 $Y2=0.054
cc_33 N_A_M2_g N_5_M4_g 2.31381e-19 $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_34 N_A_c_47_p N_5_c_58_n 0.0241209f $X=0.126 $Y=0.072 $X2=0 $Y2=0
cc_35 N_A_c_48_p N_5_c_58_n 0.00176503f $X=0.11 $Y=0.072 $X2=0 $Y2=0
cc_36 N_A_c_39_n N_5_c_59_n 4.25003e-19 $X=0.189 $Y=0.108 $X2=0 $Y2=0
cc_37 N_A_M2_g N_5_c_61_n 3.6391e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_38 N_A_M1_g N_5_c_75_n 2.2474e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_39 N_A_c_48_p N_5_c_75_n 0.00448741f $X=0.11 $Y=0.072 $X2=0 $Y2=0
cc_40 N_A_c_39_n N_5_c_62_n 9.62587e-19 $X=0.189 $Y=0.108 $X2=0 $Y2=0
cc_41 N_A_M2_g N_5_c_63_n 3.96202e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_42 N_5_c_57_n N_Y_M5_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.054
cc_43 N_5_c_57_n N_Y_M7_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_44 N_5_c_57_n N_Y_M9_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_45 N_5_c_57_n N_Y_M15_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_46 N_5_c_57_n N_Y_c_114_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_47 N_5_c_68_n N_Y_c_114_n 8.262e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_48 N_5_c_57_n N_Y_M17_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0.234 $Y2=0.162
cc_49 N_5_c_57_n N_Y_c_117_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0.109 $Y2=0.162
cc_50 N_5_c_57_n N_Y_M19_d 3.80663e-19 $X=0.567 $Y=0.135 $X2=0.126 $Y2=0.162
cc_51 N_5_c_57_n N_Y_c_119_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0.081 $Y2=0.135
cc_52 N_5_M5_g N_Y_c_120_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_53 N_5_M6_g N_Y_c_120_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_54 N_5_M7_g N_Y_c_120_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_55 N_5_M8_g N_Y_c_120_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_56 N_5_M9_g N_Y_c_120_n 4.59284e-19 $X=0.567 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_57 N_5_M4_g N_Y_c_125_n 2.73951e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_5_c_57_n N_Y_c_125_n 0.0033353f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_59 N_5_c_96_p N_Y_c_125_n 0.00198751f $X=0.288 $Y=0.198 $X2=0 $Y2=0
cc_60 N_5_M5_g N_Y_c_128_n 4.59284e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_61 N_5_M6_g N_Y_c_128_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_62 N_5_M7_g N_Y_c_128_n 4.59284e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_63 N_5_M8_g N_Y_c_128_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_5_M9_g N_Y_c_128_n 4.59284e-19 $X=0.567 $Y=0.0675 $X2=0 $Y2=0
cc_65 N_5_c_57_n N_Y_c_128_n 0.00327571f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_66 N_5_c_61_n N_Y_c_128_n 4.25902e-19 $X=0.234 $Y=0.036 $X2=0 $Y2=0
cc_67 N_5_c_57_n N_Y_c_135_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0.243 $Y2=0.162
cc_68 N_5_c_105_p N_Y_c_135_n 7.00722e-19 $X=0.288 $Y=0.079 $X2=0.243 $Y2=0.162
cc_69 N_5_c_57_n N_Y_c_137_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_70 N_5_c_57_n N_Y_c_138_n 8.00061e-19 $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_71 N_5_c_57_n Y 0.0010162f $X=0.567 $Y=0.135 $X2=0 $Y2=0
cc_72 N_5_c_63_n N_8_M13_s 4.98974e-19 $X=0.252 $Y=0.198 $X2=0.081 $Y2=0.054

* END of "./OR2x6_ASAP7_75t_R.pex.sp.OR2X6_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: OR3x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:00:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OR3x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./OR3x1_ASAP7_75t_R.pex.sp.pex"
* File: OR3x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:00:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OR3X1_ASAP7_75T_R%A 2 5 7 10 VSS
c10 10 VSS 0.00209477f $X=0.081 $Y=0.134
c11 5 VSS 0.00225666f $X=0.081 $Y=0.1355
c12 2 VSS 0.0647772f $X=0.081 $Y=0.0675
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r14 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1355 $X2=0.081 $Y2=0.2025
r15 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.1355
.ends

.subckt PM_OR3X1_ASAP7_75T_R%B 2 5 7 10 VSS
c12 10 VSS 0.00163068f $X=0.136 $Y=0.134
c13 5 VSS 0.00104174f $X=0.135 $Y=0.1355
c14 2 VSS 0.0597304f $X=0.135 $Y=0.0675
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r16 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.2025
r17 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1355
.ends

.subckt PM_OR3X1_ASAP7_75T_R%C 2 5 7 10 VSS
c12 10 VSS 0.00120766f $X=0.187 $Y=0.134
c13 5 VSS 0.00128977f $X=0.189 $Y=0.1355
c14 2 VSS 0.0591499f $X=0.189 $Y=0.0675
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1355 $X2=0.189 $Y2=0.2025
r17 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.1355
.ends

.subckt PM_OR3X1_ASAP7_75T_R%6 2 5 7 9 14 15 19 22 24 27 31 33 35 37 44 45 46 47
+ 48 50 51 52 55 56 60 VSS
c32 63 VSS 1.83894e-19 $X=0.241 $Y=0.135
c33 62 VSS 1.75291e-19 $X=0.234 $Y=0.135
c34 60 VSS 8.02486e-19 $X=0.248 $Y=0.135
c35 56 VSS 3.99142e-19 $X=0.225 $Y=0.2
c36 55 VSS 0.0010825f $X=0.225 $Y=0.183
c37 54 VSS 7.38333e-19 $X=0.225 $Y=0.225
c38 52 VSS 5.63495e-19 $X=0.225 $Y=0.094
c39 51 VSS 8.71409e-19 $X=0.225 $Y=0.07
c40 50 VSS 9.66124e-19 $X=0.225 $Y=0.126
c41 48 VSS 0.00146362f $X=0.198 $Y=0.234
c42 47 VSS 0.00329896f $X=0.18 $Y=0.234
c43 46 VSS 0.00146362f $X=0.144 $Y=0.234
c44 45 VSS 0.00356618f $X=0.126 $Y=0.234
c45 44 VSS 0.00146362f $X=0.09 $Y=0.234
c46 43 VSS 0.00433575f $X=0.072 $Y=0.234
c47 38 VSS 0.00616571f $X=0.216 $Y=0.234
c48 37 VSS 0.00146362f $X=0.198 $Y=0.036
c49 36 VSS 0.00345005f $X=0.18 $Y=0.036
c50 35 VSS 0.00146362f $X=0.144 $Y=0.036
c51 34 VSS 0.00608953f $X=0.126 $Y=0.036
c52 33 VSS 0.00146362f $X=0.09 $Y=0.036
c53 32 VSS 0.00433548f $X=0.072 $Y=0.036
c54 31 VSS 0.0105179f $X=0.162 $Y=0.036
c55 27 VSS 0.00593593f $X=0.054 $Y=0.036
c56 24 VSS 0.00575397f $X=0.216 $Y=0.036
c57 22 VSS 0.00224171f $X=0.056 $Y=0.2025
c58 19 VSS 2.69461e-19 $X=0.071 $Y=0.2025
c59 14 VSS 5.38922e-19 $X=0.179 $Y=0.0675
c60 9 VSS 2.69461e-19 $X=0.071 $Y=0.0675
c61 5 VSS 0.00384897f $X=0.243 $Y=0.135
c62 2 VSS 0.0653035f $X=0.243 $Y=0.0675
r63 62 63 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.241 $Y2=0.135
r64 60 63 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.248
+ $Y=0.135 $X2=0.241 $Y2=0.135
r65 57 62 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.135 $X2=0.234 $Y2=0.135
r66 55 56 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.183 $X2=0.225 $Y2=0.2
r67 54 56 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.225 $X2=0.225 $Y2=0.2
r68 53 57 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.144 $X2=0.225 $Y2=0.135
r69 53 55 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.144 $X2=0.225 $Y2=0.183
r70 51 52 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.07 $X2=0.225 $Y2=0.094
r71 50 57 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r72 50 52 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.094
r73 49 51 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.07
r74 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r75 46 47 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.18 $Y2=0.234
r76 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r77 44 45 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.126 $Y2=0.234
r78 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.234 $X2=0.09 $Y2=0.234
r79 40 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.072 $Y2=0.234
r80 38 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.234 $X2=0.225 $Y2=0.225
r81 38 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.198 $Y2=0.234
r82 36 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r83 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r84 33 34 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.126 $Y2=0.036
r85 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r86 30 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r87 30 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.144 $Y2=0.036
r88 30 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r89 26 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.072 $Y2=0.036
r90 26 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r91 24 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.036 $X2=0.225 $Y2=0.045
r92 24 37 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.198 $Y2=0.036
r93 22 40 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r94 19 22 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r95 18 31 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.162
+ $Y=0.0675 $X2=0.162 $Y2=0.036
r96 15 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r97 14 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r98 12 27 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r99 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r100 5 60 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.248 $Y=0.135 $X2=0.248
+ $Y2=0.135
r101 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r102 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OR3X1_ASAP7_75T_R%Y 1 4 6 9 11 19 20 21 22 31 VSS
c10 31 VSS 0.0042631f $X=0.27 $Y=0.217
c11 28 VSS 3.40666e-19 $X=0.288 $Y=0.085
c12 27 VSS 5.8248e-20 $X=0.279 $Y=0.085
c13 26 VSS 0.00155357f $X=0.297 $Y=0.085
c14 22 VSS 9.50226e-20 $X=0.27 $Y=0.085
c15 21 VSS 7.43984e-19 $X=0.297 $Y=0.144
c16 20 VSS 0.00124704f $X=0.297 $Y=0.126
c17 19 VSS 0.00150883f $X=0.297 $Y=0.1475
c18 11 VSS 0.00237937f $X=0.27 $Y=0.076
c19 9 VSS 0.00596208f $X=0.268 $Y=0.2025
c20 4 VSS 0.00611016f $X=0.268 $Y=0.0675
r21 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.085 $X2=0.288 $Y2=0.085
r22 26 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.085 $X2=0.288 $Y2=0.085
r23 22 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.085 $X2=0.279 $Y2=0.085
r24 20 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.144
r25 19 21 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.1475 $X2=0.297 $Y2=0.144
r26 17 31 1.04762 $w=3.15e-08 $l=4.65833e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.297 $Y=0.183 $X2=0.27 $Y2=0.218
r27 17 19 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.183 $X2=0.297 $Y2=0.1475
r28 16 26 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.094 $X2=0.297 $Y2=0.085
r29 16 20 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.094 $X2=0.297 $Y2=0.126
r30 11 22 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.076 $X2=0.27 $Y2=0.085
r31 11 13 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.076 $X2=0.27 $Y2=0.06
r32 9 31 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.217 $X2=0.27
+ $Y2=0.217
r33 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.2025 $X2=0.268 $Y2=0.2025
r34 4 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.06 $X2=0.27
+ $Y2=0.06
r35 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.268 $Y2=0.0675
.ends

.subckt PM_OR3X1_ASAP7_75T_R%8 1 2 VSS
c1 1 VSS 0.00183233f $X=0.125 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends

.subckt PM_OR3X1_ASAP7_75T_R%9 1 2 VSS
c1 1 VSS 0.00183233f $X=0.179 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends


* END of "./OR3x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt OR3x1_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 VSS N_A_M0_g N_6_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_6_M1_d N_B_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 VSS N_C_M2_g N_6_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_6_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_8_M4_d N_A_M4_g N_6_M4_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M5 N_9_M5_d N_B_M5_g N_8_M5_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M6 VDD N_C_M6_g N_9_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M7 N_Y_M7_d N_6_M7_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
*
* 
* .include "OR3x1_ASAP7_75t_R.pex.sp.OR3X1_ASAP7_75T_R.pxi"
* BEGIN of "./OR3x1_ASAP7_75t_R.pex.sp.OR3X1_ASAP7_75T_R.pxi"
* File: OR3x1_ASAP7_75t_R.pex.sp.OR3X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:00:25 2017
* 
x_PM_OR3X1_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M4_g A VSS
+ PM_OR3X1_ASAP7_75T_R%A
x_PM_OR3X1_ASAP7_75T_R%B N_B_M1_g N_B_c_12_n N_B_M5_g B VSS
+ PM_OR3X1_ASAP7_75T_R%B
x_PM_OR3X1_ASAP7_75T_R%C N_C_M2_g N_C_c_25_n N_C_M6_g C VSS
+ PM_OR3X1_ASAP7_75T_R%C
x_PM_OR3X1_ASAP7_75T_R%6 N_6_M3_g N_6_c_48_n N_6_M7_g N_6_M0_s N_6_M2_s N_6_M1_d
+ N_6_M4_s N_6_c_35_n N_6_c_55_p N_6_c_36_n N_6_c_42_n N_6_c_37_n N_6_c_43_n
+ N_6_c_50_n N_6_c_39_n N_6_c_65_p N_6_c_45_n N_6_c_66_p N_6_c_52_n N_6_c_60_p
+ N_6_c_63_p N_6_c_54_n N_6_c_57_p N_6_c_64_p N_6_c_62_p VSS
+ PM_OR3X1_ASAP7_75T_R%6
x_PM_OR3X1_ASAP7_75T_R%Y N_Y_M3_d N_Y_c_67_n N_Y_M7_d N_Y_c_69_n N_Y_c_70_n Y
+ N_Y_c_72_n N_Y_c_73_n N_Y_c_75_n N_Y_c_76_n VSS PM_OR3X1_ASAP7_75T_R%Y
x_PM_OR3X1_ASAP7_75T_R%8 N_8_M5_s N_8_M4_d VSS PM_OR3X1_ASAP7_75T_R%8
x_PM_OR3X1_ASAP7_75T_R%9 N_9_M6_s N_9_M5_d VSS PM_OR3X1_ASAP7_75T_R%9
cc_1 N_A_M0_g N_B_M1_g 0.00327995f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_12_n 0.00153036f $X=0.081 $Y=0.1355 $X2=0.135 $Y2=0.1355
cc_3 A B 0.00581129f $X=0.081 $Y=0.134 $X2=0.136 $Y2=0.134
cc_4 N_A_M0_g N_C_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 A N_6_c_35_n 0.00165292f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_6 A N_6_c_36_n 6.98375e-19 $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_7 N_A_M0_g N_6_c_37_n 2.64276e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_8 A N_6_c_37_n 0.00125352f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_9 N_A_M0_g N_6_c_39_n 2.63936e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_10 A N_6_c_39_n 0.00125335f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_11 N_B_M1_g N_C_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_12 N_B_c_12_n N_C_c_25_n 0.00145605f $X=0.135 $Y=0.1355 $X2=0.081 $Y2=0.1355
cc_13 B C 0.00581378f $X=0.136 $Y=0.134 $X2=0.081 $Y2=0.134
cc_14 N_B_M1_g N_6_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_15 B N_6_c_42_n 0.00114532f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_16 N_B_M1_g N_6_c_43_n 2.64276e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_17 B N_6_c_43_n 0.00125352f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_18 N_B_M1_g N_6_c_45_n 3.48272e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_19 B N_6_c_45_n 0.00125335f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_20 N_C_M2_g N_6_M3_g 0.00284417f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_21 N_C_c_25_n N_6_c_48_n 0.00128448f $X=0.189 $Y=0.1355 $X2=0.081 $Y2=0.1355
cc_22 C N_6_c_42_n 0.00114532f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_23 N_C_M2_g N_6_c_50_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_24 C N_6_c_50_n 0.00125352f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_25 N_C_M2_g N_6_c_52_n 2.63936e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_26 C N_6_c_52_n 0.00125335f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_27 C N_6_c_54_n 0.0107657f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_28 N_6_c_55_p N_Y_c_67_n 0.0011977f $X=0.216 $Y=0.036 $X2=0.081 $Y2=0.1355
cc_29 N_6_c_42_n N_Y_c_67_n 3.23836e-19 $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.1355
cc_30 N_6_c_57_p N_Y_c_69_n 0.00126271f $X=0.225 $Y=0.183 $X2=0 $Y2=0
cc_31 N_6_c_55_p N_Y_c_70_n 0.00171688f $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_32 N_6_c_57_p Y 9.77772e-19 $X=0.225 $Y=0.183 $X2=0 $Y2=0
cc_33 N_6_c_60_p N_Y_c_72_n 8.44897e-19 $X=0.225 $Y=0.126 $X2=0 $Y2=0
cc_34 N_6_c_48_n N_Y_c_73_n 3.67758e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_35 N_6_c_62_p N_Y_c_73_n 0.0011714f $X=0.248 $Y=0.135 $X2=0 $Y2=0
cc_36 N_6_c_63_p N_Y_c_75_n 0.00171688f $X=0.225 $Y=0.07 $X2=0 $Y2=0
cc_37 N_6_c_64_p N_Y_c_76_n 0.00305095f $X=0.225 $Y=0.2 $X2=0 $Y2=0
cc_38 N_6_c_65_p N_8_M5_s 3.71563e-19 $X=0.126 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_39 N_6_c_66_p N_9_M6_s 3.71563e-19 $X=0.18 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./OR3x1_ASAP7_75t_R.pex.sp.OR3X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: OR3x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:00:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OR3x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./OR3x2_ASAP7_75t_R.pex.sp.pex"
* File: OR3x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:00:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OR3X2_ASAP7_75T_R%A 2 5 7 15 VSS
c12 15 VSS 0.012188f $X=0.081 $Y=0.134
c13 5 VSS 0.00277866f $X=0.081 $Y=0.1355
c14 2 VSS 0.0654935f $X=0.081 $Y=0.0675
r15 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r16 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1355 $X2=0.081 $Y2=0.2025
r17 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.1355
.ends

.subckt PM_OR3X2_ASAP7_75T_R%B 2 5 7 12 VSS
c15 12 VSS 0.00407422f $X=0.136 $Y=0.134
c16 5 VSS 0.00107816f $X=0.135 $Y=0.1355
c17 2 VSS 0.0600722f $X=0.135 $Y=0.0675
r18 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r19 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.2025
r20 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1355
.ends

.subckt PM_OR3X2_ASAP7_75T_R%C 2 5 7 10 VSS
c13 10 VSS 0.00129842f $X=0.187 $Y=0.134
c14 5 VSS 0.00112836f $X=0.189 $Y=0.1355
c15 2 VSS 0.0583806f $X=0.189 $Y=0.0675
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1355 $X2=0.189 $Y2=0.2025
r18 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.1355
.ends

.subckt PM_OR3X2_ASAP7_75T_R%6 2 7 10 13 15 17 22 23 27 30 32 34 35 41 42 44 47
+ 50 55 57 58 59 64 65 66 69 70 72 75 78 81 VSS
c44 81 VSS 1.74783e-19 $X=0.225 $Y=0.135
c45 78 VSS 1.31878e-20 $X=0.2655 $Y=0.135
c46 77 VSS 7.16223e-19 $X=0.261 $Y=0.135
c47 75 VSS 1.63496e-19 $X=0.27 $Y=0.135
c48 72 VSS 1.87382e-19 $X=0.225 $Y=0.216
c49 71 VSS 2.19263e-19 $X=0.225 $Y=0.207
c50 70 VSS 3.97206e-19 $X=0.225 $Y=0.2
c51 69 VSS 0.00112536f $X=0.225 $Y=0.184
c52 68 VSS 1.76972e-19 $X=0.225 $Y=0.225
c53 66 VSS 4.69579e-19 $X=0.225 $Y=0.106
c54 65 VSS 3.85466e-19 $X=0.225 $Y=0.086
c55 64 VSS 2.34472e-19 $X=0.225 $Y=0.07
c56 63 VSS 3.64354e-19 $X=0.225 $Y=0.063
c57 62 VSS 7.18445e-19 $X=0.225 $Y=0.126
c58 60 VSS 0.001912f $X=0.207 $Y=0.234
c59 59 VSS 0.00142296f $X=0.198 $Y=0.234
c60 58 VSS 0.00333599f $X=0.18 $Y=0.234
c61 57 VSS 0.00308768f $X=0.144 $Y=0.234
c62 56 VSS 0.0013368f $X=0.107 $Y=0.234
c63 55 VSS 0.00369436f $X=0.095 $Y=0.234
c64 50 VSS 0.00187843f $X=0.054 $Y=0.234
c65 48 VSS 0.00421964f $X=0.216 $Y=0.234
c66 47 VSS 0.00146362f $X=0.198 $Y=0.036
c67 46 VSS 0.00258415f $X=0.18 $Y=0.036
c68 45 VSS 8.80786e-19 $X=0.153 $Y=0.036
c69 44 VSS 0.00423484f $X=0.144 $Y=0.036
c70 43 VSS 0.00238018f $X=0.107 $Y=0.036
c71 42 VSS 0.00369338f $X=0.095 $Y=0.036
c72 41 VSS 0.0106914f $X=0.162 $Y=0.036
c73 35 VSS 0.00609534f $X=0.054 $Y=0.036
c74 34 VSS 0.00187843f $X=0.054 $Y=0.036
c75 32 VSS 0.00574233f $X=0.216 $Y=0.036
c76 30 VSS 0.00242916f $X=0.056 $Y=0.2025
c77 27 VSS 3.33606e-19 $X=0.071 $Y=0.2025
c78 22 VSS 5.38922e-19 $X=0.179 $Y=0.0675
c79 17 VSS 3.33606e-19 $X=0.071 $Y=0.0675
c80 13 VSS 0.00483852f $X=0.297 $Y=0.135
c81 10 VSS 0.0639847f $X=0.297 $Y=0.0675
c82 2 VSS 0.0613335f $X=0.243 $Y=0.0675
r83 77 78 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.135 $X2=0.2655 $Y2=0.135
r84 75 78 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.135 $X2=0.2655 $Y2=0.135
r85 75 76 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.27 $Y=0.135 $X2=0.27
+ $Y2=0.135
r86 73 81 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.225 $Y2=0.135
r87 73 77 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.261 $Y2=0.135
r88 71 72 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.207 $X2=0.225 $Y2=0.216
r89 70 71 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.2 $X2=0.225 $Y2=0.207
r90 69 70 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.184 $X2=0.225 $Y2=0.2
r91 68 72 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.225 $X2=0.225 $Y2=0.216
r92 67 81 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.144 $X2=0.225 $Y2=0.135
r93 67 69 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.144 $X2=0.225 $Y2=0.184
r94 65 66 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.086 $X2=0.225 $Y2=0.106
r95 64 65 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.07 $X2=0.225 $Y2=0.086
r96 63 64 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.063 $X2=0.225 $Y2=0.07
r97 62 81 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r98 62 66 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.106
r99 61 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.063
r100 59 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.207 $Y2=0.234
r101 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r102 57 58 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.18 $Y2=0.234
r103 56 57 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.234 $X2=0.144 $Y2=0.234
r104 55 56 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.234 $X2=0.107 $Y2=0.234
r105 50 55 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.095 $Y2=0.234
r106 48 68 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.234 $X2=0.225 $Y2=0.225
r107 48 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.207 $Y2=0.234
r108 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r109 44 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.153 $Y2=0.036
r110 43 44 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.036 $X2=0.144 $Y2=0.036
r111 42 43 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.036 $X2=0.107 $Y2=0.036
r112 40 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r113 40 45 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.153 $Y2=0.036
r114 40 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r115 34 42 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.095 $Y2=0.036
r116 34 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r117 32 61 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.036 $X2=0.225 $Y2=0.045
r118 32 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.198 $Y2=0.036
r119 30 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r120 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r121 26 41 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.162 $Y=0.0675 $X2=0.162 $Y2=0.036
r122 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r123 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r124 20 35 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.054 $Y=0.0675 $X2=0.054 $Y2=0.036
r125 17 20 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r126 13 76 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.27 $Y2=0.135
r127 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.135 $X2=0.297 $Y2=0.2025
r128 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.0675 $X2=0.297 $Y2=0.135
r129 5 76 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.27 $Y2=0.135
r130 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r131 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OR3X2_ASAP7_75T_R%Y 1 2 5 6 7 10 13 18 22 24 26 28 32 34 35 36 VSS
c17 38 VSS 0.00101302f $X=0.351 $Y=0.2045
c18 36 VSS 7.93583e-20 $X=0.351 $Y=0.14575
c19 35 VSS 7.60733e-19 $X=0.351 $Y=0.144
c20 34 VSS 0.00229014f $X=0.351 $Y=0.126
c21 33 VSS 0.00176873f $X=0.351 $Y=0.086
c22 32 VSS 0.00218466f $X=0.351 $Y=0.1475
c23 30 VSS 7.5805e-19 $X=0.351 $Y=0.225
c24 28 VSS 0.00318415f $X=0.313 $Y=0.234
c25 27 VSS 3.63468e-19 $X=0.284 $Y=0.234
c26 26 VSS 0.00201509f $X=0.279 $Y=0.234
c27 25 VSS 0.00755718f $X=0.342 $Y=0.234
c28 24 VSS 0.00318415f $X=0.313 $Y=0.036
c29 23 VSS 3.63468e-19 $X=0.284 $Y=0.036
c30 22 VSS 0.00201509f $X=0.279 $Y=0.036
c31 21 VSS 0.00755718f $X=0.342 $Y=0.036
c32 18 VSS 9.19783e-19 $X=0.27 $Y=0.198
c33 13 VSS 9.19783e-19 $X=0.27 $Y=0.072
c34 10 VSS 0.0108833f $X=0.27 $Y=0.2025
c35 6 VSS 5.81027e-19 $X=0.287 $Y=0.2025
c36 5 VSS 0.0110126f $X=0.27 $Y=0.0675
c37 1 VSS 5.81027e-19 $X=0.287 $Y=0.0675
r38 37 38 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.184 $X2=0.351 $Y2=0.2045
r39 35 36 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.144 $X2=0.351 $Y2=0.14575
r40 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.144
r41 33 34 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.086 $X2=0.351 $Y2=0.126
r42 32 37 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1475 $X2=0.351 $Y2=0.184
r43 32 36 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.1475 $X2=0.351 $Y2=0.14575
r44 30 38 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.2045
r45 29 33 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.086
r46 27 28 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.234 $X2=0.313 $Y2=0.234
r47 26 27 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.234 $X2=0.284 $Y2=0.234
r48 25 30 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.234 $X2=0.351 $Y2=0.225
r49 25 28 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.313 $Y2=0.234
r50 23 24 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.036 $X2=0.313 $Y2=0.036
r51 22 23 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.036 $X2=0.284 $Y2=0.036
r52 21 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.036 $X2=0.351 $Y2=0.045
r53 21 24 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.313 $Y2=0.036
r54 16 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.27 $Y=0.225 $X2=0.279 $Y2=0.234
r55 16 18 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.225 $X2=0.27 $Y2=0.198
r56 11 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.27 $Y=0.045 $X2=0.279 $Y2=0.036
r57 11 13 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.045 $X2=0.27 $Y2=0.072
r58 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.198 $X2=0.27
+ $Y2=0.198
r59 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r60 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r61 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.072 $X2=0.27
+ $Y2=0.072
r62 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
r63 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends

.subckt PM_OR3X2_ASAP7_75T_R%8 1 2 VSS
c0 1 VSS 0.00240443f $X=0.125 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends

.subckt PM_OR3X2_ASAP7_75T_R%9 1 2 VSS
c1 1 VSS 0.00183233f $X=0.179 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends


* END of "./OR3x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt OR3x2_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 VSS N_A_M0_g N_6_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_6_M1_d N_B_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 VSS N_C_M2_g N_6_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_6_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_6_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_8_M5_d N_A_M5_g N_6_M5_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M6 N_9_M6_d N_B_M6_g N_8_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 VDD N_C_M7_g N_9_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M8 N_Y_M8_d N_6_M8_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.162
M9 N_Y_M9_d N_6_M9_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
*
* 
* .include "OR3x2_ASAP7_75t_R.pex.sp.OR3X2_ASAP7_75T_R.pxi"
* BEGIN of "./OR3x2_ASAP7_75t_R.pex.sp.OR3X2_ASAP7_75T_R.pxi"
* File: OR3x2_ASAP7_75t_R.pex.sp.OR3X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:00:48 2017
* 
x_PM_OR3X2_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M5_g A VSS
+ PM_OR3X2_ASAP7_75T_R%A
x_PM_OR3X2_ASAP7_75T_R%B N_B_M1_g N_B_c_14_n N_B_M6_g B VSS
+ PM_OR3X2_ASAP7_75T_R%B
x_PM_OR3X2_ASAP7_75T_R%C N_C_M2_g N_C_c_30_n N_C_M7_g C VSS
+ PM_OR3X2_ASAP7_75T_R%C
x_PM_OR3X2_ASAP7_75T_R%6 N_6_M3_g N_6_M8_g N_6_M4_g N_6_c_60_n N_6_M9_g N_6_M0_s
+ N_6_M2_s N_6_M1_d N_6_M5_s N_6_c_41_n N_6_c_68_p N_6_c_42_n N_6_c_43_n
+ N_6_c_51_n N_6_c_44_n N_6_c_52_n N_6_c_62_n N_6_c_46_n N_6_c_47_n N_6_c_54_n
+ N_6_c_84_p N_6_c_64_n N_6_c_56_n N_6_c_66_n N_6_c_81_p N_6_c_71_p N_6_c_74_p
+ N_6_c_78_p N_6_c_82_p N_6_c_73_p N_6_c_57_n VSS PM_OR3X2_ASAP7_75T_R%6
x_PM_OR3X2_ASAP7_75T_R%Y N_Y_M4_d N_Y_M3_d N_Y_c_86_n N_Y_M9_d N_Y_M8_d
+ N_Y_c_89_n N_Y_c_90_n N_Y_c_92_n N_Y_c_94_n N_Y_c_95_n N_Y_c_96_n N_Y_c_97_n Y
+ N_Y_c_98_n N_Y_c_100_n N_Y_c_101_n VSS PM_OR3X2_ASAP7_75T_R%Y
x_PM_OR3X2_ASAP7_75T_R%8 N_8_M6_s N_8_M5_d VSS PM_OR3X2_ASAP7_75T_R%8
x_PM_OR3X2_ASAP7_75T_R%9 N_9_M7_s N_9_M6_d VSS PM_OR3X2_ASAP7_75T_R%9
cc_1 N_A_M0_g N_B_M1_g 0.00327995f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_14_n 0.00199416f $X=0.081 $Y=0.1355 $X2=0.135 $Y2=0.1355
cc_3 A B 0.00263946f $X=0.081 $Y=0.134 $X2=0.136 $Y2=0.134
cc_4 N_A_M0_g N_C_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 A N_6_c_41_n 0.00208198f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_6 A N_6_c_42_n 0.001197f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_7 A N_6_c_43_n 0.00201602f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_8 N_A_M0_g N_6_c_44_n 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_9 A N_6_c_44_n 2.98181e-19 $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_10 A N_6_c_46_n 0.00119636f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_11 N_A_M0_g N_6_c_47_n 4.27122e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_12 A N_6_c_47_n 2.97858e-19 $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_13 N_B_M1_g N_C_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_B_c_14_n N_C_c_30_n 0.00145605f $X=0.135 $Y=0.1355 $X2=0.081 $Y2=0.1355
cc_15 B C 0.00563872f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_16 N_B_M1_g N_6_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 B N_6_c_41_n 0.00137263f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_18 B N_6_c_51_n 0.00137531f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_19 N_B_M1_g N_6_c_52_n 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_20 B N_6_c_52_n 0.00375082f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_21 N_B_M1_g N_6_c_54_n 3.22617e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_22 B N_6_c_54_n 0.00398142f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_23 B N_6_c_56_n 2.74021e-19 $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_24 B N_6_c_57_n 2.74021e-19 $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_25 N_C_M2_g N_6_M3_g 0.00284417f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_26 N_C_M2_g N_6_M4_g 2.31381e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_C_c_30_n N_6_c_60_n 0.00125914f $X=0.189 $Y=0.1355 $X2=0 $Y2=0
cc_28 C N_6_c_51_n 0.00114532f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_29 N_C_M2_g N_6_c_62_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_30 C N_6_c_62_n 0.00125352f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_31 N_C_M2_g N_6_c_64_n 2.56604e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_32 C N_6_c_64_n 0.00123587f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_33 C N_6_c_66_n 0.0107608f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_34 N_6_c_60_n N_Y_M4_d 3.80351e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_35 N_6_c_68_p N_Y_c_86_n 0.00134941f $X=0.216 $Y=0.036 $X2=0.081 $Y2=0.1355
cc_36 N_6_c_51_n N_Y_c_86_n 3.14194e-19 $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.1355
cc_37 N_6_c_60_n N_Y_M9_d 3.80351e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_38 N_6_c_71_p N_Y_c_89_n 0.00134941f $X=0.225 $Y=0.184 $X2=0 $Y2=0
cc_39 N_6_c_56_n N_Y_c_90_n 0.00177067f $X=0.225 $Y=0.07 $X2=0 $Y2=0
cc_40 N_6_c_73_p N_Y_c_90_n 4.86094e-19 $X=0.2655 $Y=0.135 $X2=0 $Y2=0
cc_41 N_6_c_74_p N_Y_c_92_n 0.00177067f $X=0.225 $Y=0.2 $X2=0.081 $Y2=0.135
cc_42 N_6_c_73_p N_Y_c_92_n 4.86094e-19 $X=0.2655 $Y=0.135 $X2=0.081 $Y2=0.135
cc_43 N_6_c_68_p N_Y_c_94_n 0.00177067f $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_44 N_6_M4_g N_Y_c_95_n 2.89885e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_45 N_6_c_78_p N_Y_c_96_n 0.00177067f $X=0.225 $Y=0.216 $X2=0 $Y2=0
cc_46 N_6_M4_g N_Y_c_97_n 2.89885e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_6_c_60_n N_Y_c_98_n 4.52406e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_48 N_6_c_81_p N_Y_c_98_n 4.04965e-19 $X=0.225 $Y=0.106 $X2=0 $Y2=0
cc_49 N_6_c_82_p N_Y_c_100_n 4.01628e-19 $X=0.27 $Y=0.135 $X2=0 $Y2=0
cc_50 N_6_c_71_p N_Y_c_101_n 4.03366e-19 $X=0.225 $Y=0.184 $X2=0 $Y2=0
cc_51 N_6_c_84_p N_9_M7_s 3.56327e-19 $X=0.18 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./OR3x2_ASAP7_75t_R.pex.sp.OR3X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: OR3x4_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:01:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OR3x4_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./OR3x4_ASAP7_75t_R.pex.sp.pex"
* File: OR3x4_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:01:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OR3X4_ASAP7_75T_R%A 2 5 7 15 VSS
c12 15 VSS 0.012188f $X=0.081 $Y=0.134
c13 5 VSS 0.00277866f $X=0.081 $Y=0.1355
c14 2 VSS 0.0654935f $X=0.081 $Y=0.0675
r15 5 15 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r16 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.1355 $X2=0.081 $Y2=0.2025
r17 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.1355
.ends

.subckt PM_OR3X4_ASAP7_75T_R%B 2 5 7 12 VSS
c15 12 VSS 0.00407422f $X=0.136 $Y=0.134
c16 5 VSS 0.00107816f $X=0.135 $Y=0.1355
c17 2 VSS 0.0600722f $X=0.135 $Y=0.0675
r18 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r19 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.2025
r20 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.1355
.ends

.subckt PM_OR3X4_ASAP7_75T_R%C 2 5 7 10 VSS
c13 10 VSS 0.00129842f $X=0.187 $Y=0.134
c14 5 VSS 0.00112836f $X=0.189 $Y=0.1355
c15 2 VSS 0.0583806f $X=0.189 $Y=0.0675
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r17 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1355 $X2=0.189 $Y2=0.2025
r18 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.1355
.ends

.subckt PM_OR3X4_ASAP7_75T_R%6 2 7 10 15 18 23 26 29 31 33 38 39 43 46 48 50 51
+ 57 58 60 63 66 71 73 74 75 80 81 85 86 88 94 97 VSS
c53 97 VSS 1.74783e-19 $X=0.225 $Y=0.135
c54 94 VSS 1.31878e-20 $X=0.2655 $Y=0.135
c55 93 VSS 7.16223e-19 $X=0.261 $Y=0.135
c56 91 VSS 2.28939e-19 $X=0.27 $Y=0.135
c57 88 VSS 1.87382e-19 $X=0.225 $Y=0.216
c58 87 VSS 2.19263e-19 $X=0.225 $Y=0.207
c59 86 VSS 3.97206e-19 $X=0.225 $Y=0.2
c60 85 VSS 0.00114186f $X=0.225 $Y=0.184
c61 84 VSS 1.76972e-19 $X=0.225 $Y=0.225
c62 82 VSS 4.69579e-19 $X=0.225 $Y=0.106
c63 81 VSS 3.85466e-19 $X=0.225 $Y=0.086
c64 80 VSS 2.34472e-19 $X=0.225 $Y=0.07
c65 79 VSS 3.64354e-19 $X=0.225 $Y=0.063
c66 78 VSS 7.34955e-19 $X=0.225 $Y=0.126
c67 76 VSS 0.001912f $X=0.207 $Y=0.234
c68 75 VSS 0.00142296f $X=0.198 $Y=0.234
c69 74 VSS 0.00333599f $X=0.18 $Y=0.234
c70 73 VSS 0.00308768f $X=0.144 $Y=0.234
c71 72 VSS 0.0013368f $X=0.107 $Y=0.234
c72 71 VSS 0.00369436f $X=0.095 $Y=0.234
c73 66 VSS 0.00187843f $X=0.054 $Y=0.234
c74 64 VSS 0.00421964f $X=0.216 $Y=0.234
c75 63 VSS 0.00146362f $X=0.198 $Y=0.036
c76 62 VSS 0.00258415f $X=0.18 $Y=0.036
c77 61 VSS 8.80786e-19 $X=0.153 $Y=0.036
c78 60 VSS 0.00423484f $X=0.144 $Y=0.036
c79 59 VSS 0.00238018f $X=0.107 $Y=0.036
c80 58 VSS 0.00369338f $X=0.095 $Y=0.036
c81 57 VSS 0.0106914f $X=0.162 $Y=0.036
c82 51 VSS 0.00609534f $X=0.054 $Y=0.036
c83 50 VSS 0.00187843f $X=0.054 $Y=0.036
c84 48 VSS 0.00574233f $X=0.216 $Y=0.036
c85 46 VSS 0.00242916f $X=0.056 $Y=0.2025
c86 43 VSS 3.33606e-19 $X=0.071 $Y=0.2025
c87 38 VSS 5.38922e-19 $X=0.179 $Y=0.0675
c88 33 VSS 3.33606e-19 $X=0.071 $Y=0.0675
c89 29 VSS 0.0156502f $X=0.405 $Y=0.135
c90 26 VSS 0.0639847f $X=0.405 $Y=0.0675
c91 18 VSS 0.0638949f $X=0.351 $Y=0.0675
c92 10 VSS 0.0636879f $X=0.297 $Y=0.0675
c93 2 VSS 0.0611266f $X=0.243 $Y=0.0675
r94 93 94 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.135 $X2=0.2655 $Y2=0.135
r95 91 94 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.135 $X2=0.2655 $Y2=0.135
r96 91 92 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.27 $Y=0.135 $X2=0.27
+ $Y2=0.135
r97 89 97 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.225 $Y2=0.135
r98 89 93 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.135 $X2=0.261 $Y2=0.135
r99 87 88 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.207 $X2=0.225 $Y2=0.216
r100 86 87 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.2 $X2=0.225 $Y2=0.207
r101 85 86 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.184 $X2=0.225 $Y2=0.2
r102 84 88 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.225 $X2=0.225 $Y2=0.216
r103 83 97 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.144 $X2=0.225 $Y2=0.135
r104 83 85 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.144 $X2=0.225 $Y2=0.184
r105 81 82 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.086 $X2=0.225 $Y2=0.106
r106 80 81 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.07 $X2=0.225 $Y2=0.086
r107 79 80 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.063 $X2=0.225 $Y2=0.07
r108 78 97 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.135
r109 78 82 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.126 $X2=0.225 $Y2=0.106
r110 77 79 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.045 $X2=0.225 $Y2=0.063
r111 75 76 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.207 $Y2=0.234
r112 74 75 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.234 $X2=0.198 $Y2=0.234
r113 73 74 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.18 $Y2=0.234
r114 72 73 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.234 $X2=0.144 $Y2=0.234
r115 71 72 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.234 $X2=0.107 $Y2=0.234
r116 66 71 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.095 $Y2=0.234
r117 64 84 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.234 $X2=0.225 $Y2=0.225
r118 64 76 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.207 $Y2=0.234
r119 62 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r120 60 61 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.153 $Y2=0.036
r121 59 60 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.036 $X2=0.144 $Y2=0.036
r122 58 59 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.036 $X2=0.107 $Y2=0.036
r123 56 62 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r124 56 61 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.153 $Y2=0.036
r125 56 57 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r126 50 58 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.095 $Y2=0.036
r127 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r128 48 77 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.036 $X2=0.225 $Y2=0.045
r129 48 63 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.198 $Y2=0.036
r130 46 66 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r131 43 46 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r132 42 57 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.162 $Y=0.0675 $X2=0.162 $Y2=0.036
r133 39 42 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r134 38 42 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r135 36 51 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.054 $Y=0.0675 $X2=0.054 $Y2=0.036
r136 33 36 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r137 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r138 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r139 21 29 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r140 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r141 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r142 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r143 13 92 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.27 $Y2=0.135
r144 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.135 $X2=0.297 $Y2=0.2025
r145 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.297 $Y=0.0675 $X2=0.297 $Y2=0.135
r146 5 92 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.243
+ $Y=0.135 $X2=0.27 $Y2=0.135
r147 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r148 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OR3X4_ASAP7_75T_R%Y 1 2 5 6 7 10 11 12 15 16 17 20 23 28 31 32 34 35
+ 36 38 41 46 49 51 56 58 VSS
c26 64 VSS 0.00150149f $X=0.378 $Y=0.234
c27 63 VSS 0.00150149f $X=0.378 $Y=0.036
c28 62 VSS 0.00101302f $X=0.459 $Y=0.2045
c29 60 VSS 7.51787e-20 $X=0.459 $Y=0.14575
c30 59 VSS 8.67879e-19 $X=0.459 $Y=0.144
c31 58 VSS 0.00285296f $X=0.459 $Y=0.126
c32 57 VSS 0.00176873f $X=0.459 $Y=0.086
c33 56 VSS 0.00274913f $X=0.459 $Y=0.1475
c34 54 VSS 7.5805e-19 $X=0.459 $Y=0.225
c35 51 VSS 0.0112873f $X=0.45 $Y=0.234
c36 49 VSS 0.0112873f $X=0.45 $Y=0.036
c37 46 VSS 0.00117559f $X=0.378 $Y=0.198
c38 41 VSS 0.00117559f $X=0.378 $Y=0.072
c39 38 VSS 0.00525658f $X=0.3265 $Y=0.234
c40 37 VSS 3.63468e-19 $X=0.284 $Y=0.234
c41 36 VSS 0.0020097f $X=0.279 $Y=0.234
c42 35 VSS 0.00484981f $X=0.369 $Y=0.234
c43 34 VSS 0.00525658f $X=0.3265 $Y=0.036
c44 33 VSS 3.63468e-19 $X=0.284 $Y=0.036
c45 32 VSS 0.0020097f $X=0.279 $Y=0.036
c46 31 VSS 0.00484981f $X=0.369 $Y=0.036
c47 28 VSS 5.19852e-19 $X=0.27 $Y=0.198
c48 23 VSS 5.19852e-19 $X=0.27 $Y=0.072
c49 20 VSS 0.0105054f $X=0.378 $Y=0.2025
c50 16 VSS 5.38922e-19 $X=0.395 $Y=0.2025
c51 15 VSS 0.0108685f $X=0.27 $Y=0.2025
c52 11 VSS 5.81027e-19 $X=0.287 $Y=0.2025
c53 10 VSS 0.0105054f $X=0.378 $Y=0.0675
c54 6 VSS 5.38922e-19 $X=0.395 $Y=0.0675
c55 5 VSS 0.0109978f $X=0.27 $Y=0.0675
c56 1 VSS 5.81027e-19 $X=0.287 $Y=0.0675
r57 61 62 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.184 $X2=0.459 $Y2=0.2045
r58 59 60 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.144 $X2=0.459 $Y2=0.14575
r59 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.126 $X2=0.459 $Y2=0.144
r60 57 58 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.086 $X2=0.459 $Y2=0.126
r61 56 61 2.47839 $w=1.8e-08 $l=3.65e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.1475 $X2=0.459 $Y2=0.184
r62 56 60 0.118827 $w=1.8e-08 $l=1.75e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.1475 $X2=0.459 $Y2=0.14575
r63 54 62 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.2045
r64 53 57 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.086
r65 52 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.387
+ $Y=0.234 $X2=0.378 $Y2=0.234
r66 51 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r67 51 52 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.387 $Y2=0.234
r68 50 63 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.387
+ $Y=0.036 $X2=0.378 $Y2=0.036
r69 49 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r70 49 50 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.387 $Y2=0.036
r71 44 64 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.225 $X2=0.378 $Y2=0.234
r72 44 46 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.225 $X2=0.378 $Y2=0.198
r73 39 63 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.045 $X2=0.378 $Y2=0.036
r74 39 41 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.045 $X2=0.378 $Y2=0.072
r75 37 38 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.234 $X2=0.3265 $Y2=0.234
r76 36 37 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.234 $X2=0.284 $Y2=0.234
r77 35 64 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.369
+ $Y=0.234 $X2=0.378 $Y2=0.234
r78 35 38 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.369
+ $Y=0.234 $X2=0.3265 $Y2=0.234
r79 33 34 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.036 $X2=0.3265 $Y2=0.036
r80 32 33 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.036 $X2=0.284 $Y2=0.036
r81 31 63 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.369
+ $Y=0.036 $X2=0.378 $Y2=0.036
r82 31 34 2.8858 $w=1.8e-08 $l=4.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.369
+ $Y=0.036 $X2=0.3265 $Y2=0.036
r83 26 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.27 $Y=0.225 $X2=0.279 $Y2=0.234
r84 26 28 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.225 $X2=0.27 $Y2=0.198
r85 21 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.27 $Y=0.045 $X2=0.279 $Y2=0.036
r86 21 23 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.045 $X2=0.27 $Y2=0.072
r87 20 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.198 $X2=0.378
+ $Y2=0.198
r88 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r89 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r90 15 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.198 $X2=0.27
+ $Y2=0.198
r91 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r92 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r93 10 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.072 $X2=0.378
+ $Y2=0.072
r94 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.0675 $X2=0.378 $Y2=0.0675
r95 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.0675 $X2=0.378 $Y2=0.0675
r96 5 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.072 $X2=0.27
+ $Y2=0.072
r97 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
r98 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends

.subckt PM_OR3X4_ASAP7_75T_R%8 1 2 VSS
c0 1 VSS 0.00240443f $X=0.125 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends

.subckt PM_OR3X4_ASAP7_75T_R%9 1 2 VSS
c1 1 VSS 0.00183233f $X=0.179 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends


* END of "./OR3x4_ASAP7_75t_R.pex.sp.pex"
* 
.subckt OR3x4_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 VSS N_A_M0_g N_6_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_6_M1_d N_B_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 VSS N_C_M2_g N_6_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_6_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_Y_M4_d N_6_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_6_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_6_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_8_M7_d N_A_M7_g N_6_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M8 N_9_M8_d N_B_M8_g N_8_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M9 VDD N_C_M9_g N_9_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M10 N_Y_M10_d N_6_M10_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M11 N_Y_M11_d N_6_M11_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M12 N_Y_M12_d N_6_M12_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M13 N_Y_M13_d N_6_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
*
* 
* .include "OR3x4_ASAP7_75t_R.pex.sp.OR3X4_ASAP7_75T_R.pxi"
* BEGIN of "./OR3x4_ASAP7_75t_R.pex.sp.OR3X4_ASAP7_75T_R.pxi"
* File: OR3x4_ASAP7_75t_R.pex.sp.OR3X4_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:01:10 2017
* 
x_PM_OR3X4_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M7_g A VSS
+ PM_OR3X4_ASAP7_75T_R%A
x_PM_OR3X4_ASAP7_75T_R%B N_B_M1_g N_B_c_14_n N_B_M8_g B VSS
+ PM_OR3X4_ASAP7_75T_R%B
x_PM_OR3X4_ASAP7_75T_R%C N_C_M2_g N_C_c_30_n N_C_M9_g C VSS
+ PM_OR3X4_ASAP7_75T_R%C
x_PM_OR3X4_ASAP7_75T_R%6 N_6_M3_g N_6_M10_g N_6_M4_g N_6_M11_g N_6_M5_g
+ N_6_M12_g N_6_M6_g N_6_c_60_n N_6_M13_g N_6_M0_s N_6_M2_s N_6_M1_d N_6_M7_s
+ N_6_c_41_n N_6_c_68_p N_6_c_42_n N_6_c_43_n N_6_c_51_n N_6_c_44_n N_6_c_52_n
+ N_6_c_62_n N_6_c_46_n N_6_c_47_n N_6_c_54_n N_6_c_93_p N_6_c_64_n N_6_c_56_n
+ N_6_c_66_n N_6_c_73_p N_6_c_78_p N_6_c_85_p N_6_c_77_p N_6_c_57_n VSS
+ PM_OR3X4_ASAP7_75T_R%6
x_PM_OR3X4_ASAP7_75T_R%Y N_Y_M4_d N_Y_M3_d N_Y_c_95_n N_Y_M6_d N_Y_M5_d
+ N_Y_c_98_n N_Y_M11_d N_Y_M10_d N_Y_c_100_n N_Y_M13_d N_Y_M12_d N_Y_c_102_n
+ N_Y_c_103_n N_Y_c_105_n N_Y_c_107_n N_Y_c_108_n N_Y_c_109_n N_Y_c_111_n
+ N_Y_c_112_n N_Y_c_113_n N_Y_c_115_n N_Y_c_116_n N_Y_c_117_n N_Y_c_118_n Y
+ N_Y_c_119_n VSS PM_OR3X4_ASAP7_75T_R%Y
x_PM_OR3X4_ASAP7_75T_R%8 N_8_M8_s N_8_M7_d VSS PM_OR3X4_ASAP7_75T_R%8
x_PM_OR3X4_ASAP7_75T_R%9 N_9_M9_s N_9_M8_d VSS PM_OR3X4_ASAP7_75T_R%9
cc_1 N_A_M0_g N_B_M1_g 0.00327995f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_14_n 0.00199416f $X=0.081 $Y=0.1355 $X2=0.135 $Y2=0.1355
cc_3 A B 0.00263946f $X=0.081 $Y=0.134 $X2=0.136 $Y2=0.134
cc_4 N_A_M0_g N_C_M2_g 2.66145e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_5 A N_6_c_41_n 0.00208198f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_6 A N_6_c_42_n 0.001197f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_7 A N_6_c_43_n 0.00201602f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_8 N_A_M0_g N_6_c_44_n 4.28653e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_9 A N_6_c_44_n 2.98181e-19 $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_10 A N_6_c_46_n 0.00119636f $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_11 N_A_M0_g N_6_c_47_n 4.27122e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_12 A N_6_c_47_n 2.97858e-19 $X=0.081 $Y=0.134 $X2=0 $Y2=0
cc_13 N_B_M1_g N_C_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_14 N_B_c_14_n N_C_c_30_n 0.00145605f $X=0.135 $Y=0.1355 $X2=0.081 $Y2=0.1355
cc_15 B C 0.00563872f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_16 N_B_M1_g N_6_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_17 B N_6_c_41_n 0.00137263f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_18 B N_6_c_51_n 0.00137531f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_19 N_B_M1_g N_6_c_52_n 2.34993e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_20 B N_6_c_52_n 0.00375082f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_21 N_B_M1_g N_6_c_54_n 3.22617e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_22 B N_6_c_54_n 0.00398142f $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_23 B N_6_c_56_n 2.74021e-19 $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_24 B N_6_c_57_n 2.74021e-19 $X=0.136 $Y=0.134 $X2=0 $Y2=0
cc_25 N_C_M2_g N_6_M3_g 0.00284417f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_26 N_C_M2_g N_6_M4_g 2.31381e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_C_c_30_n N_6_c_60_n 0.00125078f $X=0.189 $Y=0.1355 $X2=0 $Y2=0
cc_28 C N_6_c_51_n 0.00114532f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_29 N_C_M2_g N_6_c_62_n 2.64276e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_30 C N_6_c_62_n 0.00125352f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_31 N_C_M2_g N_6_c_64_n 2.56604e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_32 C N_6_c_64_n 0.00123587f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_33 C N_6_c_66_n 0.0107608f $X=0.187 $Y=0.134 $X2=0 $Y2=0
cc_34 N_6_c_60_n N_Y_M4_d 3.80351e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_35 N_6_c_68_p N_Y_c_95_n 0.00112271f $X=0.216 $Y=0.036 $X2=0.081 $Y2=0.1355
cc_36 N_6_c_51_n N_Y_c_95_n 3.14194e-19 $X=0.162 $Y=0.036 $X2=0.081 $Y2=0.1355
cc_37 N_6_c_60_n N_Y_M6_d 3.80663e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_38 N_6_c_60_n N_Y_c_98_n 8.00061e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_39 N_6_c_60_n N_Y_M11_d 3.80351e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_40 N_6_c_73_p N_Y_c_100_n 0.00112271f $X=0.225 $Y=0.184 $X2=0.081 $Y2=0.134
cc_41 N_6_c_60_n N_Y_M13_d 3.80663e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_42 N_6_c_60_n N_Y_c_102_n 8.00061e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_43 N_6_c_56_n N_Y_c_103_n 0.00179666f $X=0.225 $Y=0.07 $X2=0 $Y2=0
cc_44 N_6_c_77_p N_Y_c_103_n 4.86094e-19 $X=0.2655 $Y=0.135 $X2=0 $Y2=0
cc_45 N_6_c_78_p N_Y_c_105_n 0.00179666f $X=0.225 $Y=0.2 $X2=0 $Y2=0
cc_46 N_6_c_77_p N_Y_c_105_n 4.86094e-19 $X=0.2655 $Y=0.135 $X2=0 $Y2=0
cc_47 N_6_M5_g N_Y_c_107_n 2.89885e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_48 N_6_c_68_p N_Y_c_108_n 0.00179666f $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_49 N_6_M4_g N_Y_c_109_n 2.89885e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_50 N_6_c_60_n N_Y_c_109_n 7.93486e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_51 N_6_M5_g N_Y_c_111_n 2.89885e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_52 N_6_c_85_p N_Y_c_112_n 0.00179666f $X=0.225 $Y=0.216 $X2=0 $Y2=0
cc_53 N_6_M4_g N_Y_c_113_n 2.89885e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_54 N_6_c_60_n N_Y_c_113_n 7.93486e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_55 N_6_c_60_n N_Y_c_115_n 2.47493e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_56 N_6_c_60_n N_Y_c_116_n 2.47493e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_57 N_6_M6_g N_Y_c_117_n 2.89885e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_58 N_6_M6_g N_Y_c_118_n 2.89885e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_59 N_6_c_60_n N_Y_c_119_n 9.12721e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_60 N_6_c_93_p N_9_M9_s 3.56327e-19 $X=0.18 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./OR3x4_ASAP7_75t_R.pex.sp.OR3X4_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: OR4x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:01:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OR4x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./OR4x1_ASAP7_75t_R.pex.sp.pex"
* File: OR4x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:01:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OR4X1_ASAP7_75T_R%3 2 5 7 9 10 14 15 19 22 26 27 28 29 30 33 35 38 40
+ 45 46 48 51 58 59 63 65 66 73 VSS
c36 73 VSS 0.00417997f $X=0.342 $Y=0.234
c37 72 VSS 0.00278493f $X=0.351 $Y=0.234
c38 66 VSS 1.79388e-19 $X=0.068 $Y=0.135
c39 65 VSS 3.47369e-19 $X=0.063 $Y=0.135
c40 63 VSS 8.71424e-19 $X=0.081 $Y=0.135
c41 59 VSS 4.30865e-19 $X=0.351 $Y=0.2125
c42 58 VSS 0.0057844f $X=0.351 $Y=0.2
c43 57 VSS 4.01444e-19 $X=0.351 $Y=0.07
c44 56 VSS 0.00108941f $X=0.351 $Y=0.063
c45 55 VSS 8.62726e-19 $X=0.351 $Y=0.225
c46 53 VSS 0.00289269f $X=0.326 $Y=0.036
c47 52 VSS 3.40854e-19 $X=0.31 $Y=0.036
c48 51 VSS 0.00146362f $X=0.306 $Y=0.036
c49 50 VSS 0.0027713f $X=0.288 $Y=0.036
c50 49 VSS 9.5272e-19 $X=0.261 $Y=0.036
c51 48 VSS 0.00142296f $X=0.252 $Y=0.036
c52 47 VSS 0.00678169f $X=0.234 $Y=0.036
c53 46 VSS 0.00286574f $X=0.198 $Y=0.036
c54 45 VSS 0.0104492f $X=0.27 $Y=0.036
c55 41 VSS 0.00169362f $X=0.161 $Y=0.036
c56 40 VSS 0.00146362f $X=0.144 $Y=0.036
c57 39 VSS 0.00149782f $X=0.126 $Y=0.036
c58 38 VSS 0.0103752f $X=0.162 $Y=0.036
c59 35 VSS 0.00329991f $X=0.117 $Y=0.036
c60 34 VSS 0.00586463f $X=0.342 $Y=0.036
c61 33 VSS 6.41935e-19 $X=0.108 $Y=0.063
c62 31 VSS 0.00126924f $X=0.096 $Y=0.072
c63 30 VSS 1.4325e-20 $X=0.068 $Y=0.072
c64 29 VSS 5.64827e-20 $X=0.063 $Y=0.072
c65 28 VSS 0.0018601f $X=0.099 $Y=0.072
c66 27 VSS 1.71598e-19 $X=0.054 $Y=0.116
c67 26 VSS 4.86765e-19 $X=0.054 $Y=0.106
c68 25 VSS 1.7063e-19 $X=0.054 $Y=0.126
c69 22 VSS 0.00369079f $X=0.322 $Y=0.2025
c70 14 VSS 6.1012e-19 $X=0.287 $Y=0.0675
c71 9 VSS 6.55441e-19 $X=0.179 $Y=0.0675
c72 5 VSS 0.00217304f $X=0.081 $Y=0.135
c73 2 VSS 0.0651846f $X=0.081 $Y=0.0675
r74 73 74 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.3465 $Y2=0.234
r75 72 74 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.234 $X2=0.3465 $Y2=0.234
r76 69 73 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.342 $Y2=0.234
r77 65 66 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.135 $X2=0.068 $Y2=0.135
r78 63 66 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.068 $Y2=0.135
r79 60 65 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.135 $X2=0.063 $Y2=0.135
r80 58 59 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.2 $X2=0.351 $Y2=0.2125
r81 57 58 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.07 $X2=0.351 $Y2=0.2
r82 56 57 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.063 $X2=0.351 $Y2=0.07
r83 55 72 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.234
r84 55 59 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.225 $X2=0.351 $Y2=0.2125
r85 54 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.045 $X2=0.351 $Y2=0.063
r86 52 53 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.31
+ $Y=0.036 $X2=0.326 $Y2=0.036
r87 51 52 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.31 $Y2=0.036
r88 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r89 48 49 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.261 $Y2=0.036
r90 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r91 46 47 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.234 $Y2=0.036
r92 44 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.288 $Y2=0.036
r93 44 49 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.261 $Y2=0.036
r94 44 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r95 41 42 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.161
+ $Y=0.036 $X2=0.1615 $Y2=0.036
r96 40 41 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.161 $Y2=0.036
r97 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r98 37 46 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.198 $Y2=0.036
r99 37 42 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.1615 $Y2=0.036
r100 37 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r101 35 39 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.036 $X2=0.126 $Y2=0.036
r102 34 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.036 $X2=0.351 $Y2=0.045
r103 34 53 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.326 $Y2=0.036
r104 32 35 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.108 $Y=0.045 $X2=0.117 $Y2=0.036
r105 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.045 $X2=0.108 $Y2=0.063
r106 30 31 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.068
+ $Y=0.072 $X2=0.096 $Y2=0.072
r107 29 30 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.072 $X2=0.068 $Y2=0.072
r108 28 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.099 $Y=0.072 $X2=0.108 $Y2=0.063
r109 28 31 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.072 $X2=0.096 $Y2=0.072
r110 26 27 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.106 $X2=0.054 $Y2=0.116
r111 25 60 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.126 $X2=0.054 $Y2=0.135
r112 25 27 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.126 $X2=0.054 $Y2=0.116
r113 24 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.054 $Y=0.081 $X2=0.063 $Y2=0.072
r114 24 26 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.081 $X2=0.054 $Y2=0.106
r115 22 69 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234
+ $X2=0.324 $Y2=0.234
r116 19 22 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.2025 $X2=0.322 $Y2=0.2025
r117 18 45 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r118 15 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r119 14 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r120 13 38 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.162 $Y=0.0675 $X2=0.162 $Y2=0.036
r121 10 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.162 $Y2=0.0675
r122 9 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.0675 $X2=0.162 $Y2=0.0675
r123 5 63 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r124 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r125 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OR4X1_ASAP7_75T_R%D 2 5 7 11 VSS
c11 11 VSS 0.0046622f $X=0.135 $Y=0.132
c12 5 VSS 0.00117848f $X=0.135 $Y=0.135
c13 2 VSS 0.0594773f $X=0.135 $Y=0.0675
r14 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r15 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r16 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_OR4X1_ASAP7_75T_R%C 2 5 7 12 VSS
c14 12 VSS 0.00782796f $X=0.189 $Y=0.132
c15 5 VSS 0.00165807f $X=0.189 $Y=0.135
c16 2 VSS 0.0598363f $X=0.189 $Y=0.0675
r17 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OR4X1_ASAP7_75T_R%B 2 5 7 10 VSS
c13 10 VSS 0.00272832f $X=0.243 $Y=0.132
c14 5 VSS 0.00115441f $X=0.243 $Y=0.135
c15 2 VSS 0.060052f $X=0.243 $Y=0.0675
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OR4X1_ASAP7_75T_R%A 2 5 7 10 VSS
c9 10 VSS 0.00227875f $X=0.297 $Y=0.132
c10 5 VSS 0.00229951f $X=0.297 $Y=0.135
c11 2 VSS 0.0641834f $X=0.297 $Y=0.0675
r12 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OR4X1_ASAP7_75T_R%Y 1 6 14 16 18 23 24 26 30 33 VSS
c16 33 VSS 3.47399e-19 $X=0.0495 $Y=0.234
c17 32 VSS 0.00216674f $X=0.045 $Y=0.234
c18 30 VSS 0.00248716f $X=0.054 $Y=0.234
c19 28 VSS 0.00317012f $X=0.027 $Y=0.234
c20 26 VSS 3.3597e-19 $X=0.0495 $Y=0.036
c21 25 VSS 0.00216674f $X=0.045 $Y=0.036
c22 24 VSS 0.00627446f $X=0.054 $Y=0.036
c23 23 VSS 0.00218773f $X=0.054 $Y=0.036
c24 21 VSS 0.00318295f $X=0.027 $Y=0.036
c25 20 VSS 4.26553e-19 $X=0.018 $Y=0.216
c26 19 VSS 9.0411e-19 $X=0.018 $Y=0.207
c27 18 VSS 0.00222465f $X=0.018 $Y=0.189
c28 16 VSS 0.00131588f $X=0.018 $Y=0.0975
c29 15 VSS 8.54366e-19 $X=0.018 $Y=0.063
c30 14 VSS 0.00182881f $X=0.016 $Y=0.132
c31 12 VSS 4.02856e-19 $X=0.018 $Y=0.225
c32 9 VSS 0.00560367f $X=0.056 $Y=0.2025
c33 6 VSS 3.68013e-19 $X=0.071 $Y=0.2025
c34 1 VSS 3.75928e-19 $X=0.071 $Y=0.0675
r35 32 33 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.045
+ $Y=0.234 $X2=0.0495 $Y2=0.234
r36 30 33 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.0495 $Y2=0.234
r37 28 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.045 $Y2=0.234
r38 25 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.045
+ $Y=0.036 $X2=0.0495 $Y2=0.036
r39 23 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.0495 $Y2=0.036
r40 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r41 21 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.045 $Y2=0.036
r42 19 20 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.207 $X2=0.018 $Y2=0.216
r43 18 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.207
r44 17 18 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.189
r45 15 16 2.34259 $w=1.8e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.0975
r46 14 17 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.132 $X2=0.018 $Y2=0.144
r47 14 16 2.34259 $w=1.8e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.132 $X2=0.018 $Y2=0.0975
r48 12 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r49 12 20 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.216
r50 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r51 11 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r52 9 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r53 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
r54 4 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r55 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends

.subckt PM_OR4X1_ASAP7_75T_R%9 1 2 VSS
c1 1 VSS 0.00214488f $X=0.179 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends

.subckt PM_OR4X1_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00228146f $X=0.233 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.199 $Y2=0.2025
.ends

.subckt PM_OR4X1_ASAP7_75T_R%11 1 2 VSS
c0 1 VSS 0.00228146f $X=0.287 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.253 $Y2=0.2025
.ends


* END of "./OR4x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt OR4x1_ASAP7_75t_R  VSS VDD D C B A Y
* 
* Y	Y
* A	A
* B	B
* C	C
* D	D
M0 VSS N_3_M0_g N_Y_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_3_M1_d N_D_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 VSS N_C_M2_g N_3_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_3_M3_d N_B_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 VSS N_A_M4_g N_3_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 VDD N_3_M5_g N_Y_M5_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M6 N_9_M6_d N_D_M6_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M7 N_10_M7_d N_C_M7_g N_9_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M8 N_11_M8_d N_B_M8_g N_10_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M9 N_3_M9_d N_A_M9_g N_11_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
*
* 
* .include "OR4x1_ASAP7_75t_R.pex.sp.OR4X1_ASAP7_75T_R.pxi"
* BEGIN of "./OR4x1_ASAP7_75t_R.pex.sp.OR4X1_ASAP7_75T_R.pxi"
* File: OR4x1_ASAP7_75t_R.pex.sp.OR4X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:01:33 2017
* 
x_PM_OR4X1_ASAP7_75T_R%3 N_3_M0_g N_3_c_3_p N_3_M5_g N_3_M2_s N_3_M1_d N_3_M4_s
+ N_3_M3_d N_3_M9_d N_3_c_13_p N_3_c_28_p N_3_c_4_p N_3_c_9_p N_3_c_25_p
+ N_3_c_26_p N_3_c_32_p N_3_c_27_p N_3_c_10_p N_3_c_2_p N_3_c_14_p N_3_c_8_p
+ N_3_c_12_p N_3_c_18_p N_3_c_22_p N_3_c_16_p N_3_c_6_p N_3_c_36_p N_3_c_35_p
+ N_3_c_17_p VSS PM_OR4X1_ASAP7_75T_R%3
x_PM_OR4X1_ASAP7_75T_R%D N_D_M1_g N_D_c_39_n N_D_M6_g D VSS
+ PM_OR4X1_ASAP7_75T_R%D
x_PM_OR4X1_ASAP7_75T_R%C N_C_M2_g N_C_c_54_n N_C_M7_g C VSS
+ PM_OR4X1_ASAP7_75T_R%C
x_PM_OR4X1_ASAP7_75T_R%B N_B_M3_g N_B_c_70_n N_B_M8_g B VSS
+ PM_OR4X1_ASAP7_75T_R%B
x_PM_OR4X1_ASAP7_75T_R%A N_A_M4_g N_A_c_82_n N_A_M9_g A VSS
+ PM_OR4X1_ASAP7_75T_R%A
x_PM_OR4X1_ASAP7_75T_R%Y N_Y_M0_s N_Y_M5_s Y N_Y_c_86_n N_Y_c_98_n N_Y_c_87_n
+ N_Y_c_89_n N_Y_c_95_n N_Y_c_96_n N_Y_c_97_n VSS PM_OR4X1_ASAP7_75T_R%Y
x_PM_OR4X1_ASAP7_75T_R%9 N_9_M7_s N_9_M6_d VSS PM_OR4X1_ASAP7_75T_R%9
x_PM_OR4X1_ASAP7_75T_R%10 N_10_M8_s N_10_M7_d VSS PM_OR4X1_ASAP7_75T_R%10
x_PM_OR4X1_ASAP7_75T_R%11 N_11_M9_s N_11_M8_d VSS PM_OR4X1_ASAP7_75T_R%11
cc_1 N_3_M0_g N_D_M1_g 0.00284417f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_3_c_2_p N_D_M1_g 3.59101e-19 $X=0.144 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_3 N_3_c_3_p N_D_c_39_n 9.86475e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_3_c_4_p D 5.52051e-19 $X=0.054 $Y=0.116 $X2=0.135 $Y2=0.132
cc_5 N_3_c_2_p D 5.39549e-19 $X=0.144 $Y=0.036 $X2=0.135 $Y2=0.132
cc_6 N_3_c_6_p D 8.96322e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.132
cc_7 N_3_M0_g N_C_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_8 N_3_c_8_p N_C_M2_g 2.35421e-19 $X=0.198 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_9 N_3_c_9_p C 4.85889e-19 $X=0.099 $Y=0.072 $X2=0 $Y2=0
cc_10 N_3_c_10_p C 0.00210911f $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_11 N_3_c_8_p C 0.00373267f $X=0.198 $Y=0.036 $X2=0 $Y2=0
cc_12 N_3_c_12_p N_B_M3_g 2.57255e-19 $X=0.252 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_13 N_3_c_13_p B 4.68998e-19 $X=0.322 $Y=0.2025 $X2=0 $Y2=0
cc_14 N_3_c_14_p B 0.00114532f $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_15 N_3_c_12_p B 0.00123937f $X=0.252 $Y=0.036 $X2=0 $Y2=0
cc_16 N_3_c_16_p B 2.69891e-19 $X=0.351 $Y=0.2125 $X2=0 $Y2=0
cc_17 N_3_c_17_p B 4.44922e-19 $X=0.342 $Y=0.234 $X2=0 $Y2=0
cc_18 N_3_c_18_p N_A_M4_g 2.64924e-19 $X=0.306 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_19 N_3_c_13_p A 0.0013295f $X=0.322 $Y=0.2025 $X2=0 $Y2=0
cc_20 N_3_c_14_p A 0.00114532f $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_21 N_3_c_18_p A 0.00125383f $X=0.306 $Y=0.036 $X2=0 $Y2=0
cc_22 N_3_c_22_p A 0.00499854f $X=0.351 $Y=0.2 $X2=0 $Y2=0
cc_23 N_3_c_3_p Y 2.37651e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_24 N_3_c_4_p Y 0.00364616f $X=0.054 $Y=0.116 $X2=0 $Y2=0
cc_25 N_3_c_25_p N_Y_c_86_n 0.00364616f $X=0.063 $Y=0.072 $X2=0.135 $Y2=0.135
cc_26 N_3_c_26_p N_Y_c_87_n 8.91894e-19 $X=0.068 $Y=0.072 $X2=0 $Y2=0
cc_27 N_3_c_27_p N_Y_c_87_n 9.22842e-19 $X=0.117 $Y=0.036 $X2=0 $Y2=0
cc_28 N_3_c_28_p N_Y_c_89_n 0.00136707f $X=0.054 $Y=0.106 $X2=0 $Y2=0
cc_29 N_3_c_4_p N_Y_c_89_n 6.1755e-19 $X=0.054 $Y=0.116 $X2=0 $Y2=0
cc_30 N_3_c_25_p N_Y_c_89_n 0.0011724f $X=0.063 $Y=0.072 $X2=0 $Y2=0
cc_31 N_3_c_26_p N_Y_c_89_n 5.48981e-19 $X=0.068 $Y=0.072 $X2=0 $Y2=0
cc_32 N_3_c_32_p N_Y_c_89_n 2.94367e-19 $X=0.108 $Y=0.063 $X2=0 $Y2=0
cc_33 N_3_c_10_p N_Y_c_89_n 2.28909e-19 $X=0.162 $Y=0.036 $X2=0 $Y2=0
cc_34 N_3_c_25_p N_Y_c_95_n 8.91894e-19 $X=0.063 $Y=0.072 $X2=0 $Y2=0
cc_35 N_3_c_35_p N_Y_c_96_n 2.48124e-19 $X=0.068 $Y=0.135 $X2=0 $Y2=0
cc_36 N_3_c_36_p N_Y_c_97_n 2.48124e-19 $X=0.063 $Y=0.135 $X2=0 $Y2=0
cc_37 N_D_M1_g N_C_M2_g 0.00344695f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_38 N_D_c_39_n N_C_c_54_n 7.51247e-19 $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_39 D C 0.00489513f $X=0.135 $Y=0.132 $X2=0 $Y2=0
cc_40 N_D_M1_g N_B_M3_g 2.66145e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_41 D N_Y_c_98_n 4.90231e-19 $X=0.135 $Y=0.132 $X2=0.27 $Y2=0.0675
cc_42 N_C_M2_g N_B_M3_g 0.00327995f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_43 N_C_c_54_n N_B_c_70_n 7.51247e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_44 C B 0.00749132f $X=0.189 $Y=0.132 $X2=0.145 $Y2=0.0675
cc_45 N_C_M2_g N_A_M4_g 2.71887e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_46 C N_Y_c_96_n 2.2335e-19 $X=0.189 $Y=0.132 $X2=0.068 $Y2=0.072
cc_47 C N_9_M7_s 2.91005e-19 $X=0.189 $Y=0.132 $X2=0.081 $Y2=0.0675
cc_48 N_B_M3_g N_A_M4_g 0.00357042f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_49 N_B_c_70_n N_A_c_82_n 7.51046e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_50 B A 0.0057113f $X=0.243 $Y=0.132 $X2=0.145 $Y2=0.0675

* END of "./OR4x1_ASAP7_75t_R.pex.sp.OR4X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: OR4x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:01:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OR4x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./OR4x2_ASAP7_75t_R.pex.sp.pex"
* File: OR4x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:01:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OR4X2_ASAP7_75T_R%3 2 5 7 10 13 15 17 18 22 23 27 30 34 35 36 37 38
+ 43 46 48 53 54 56 59 66 67 73 76 78 86 VSS
c38 86 VSS 0.00417997f $X=0.396 $Y=0.234
c39 85 VSS 0.00278493f $X=0.405 $Y=0.234
c40 79 VSS 1.14182e-19 $X=0.122 $Y=0.135
c41 78 VSS 5.32186e-20 $X=0.117 $Y=0.135
c42 76 VSS 8.74201e-19 $X=0.135 $Y=0.135
c43 73 VSS 8.11001e-19 $X=0.099 $Y=0.135
c44 67 VSS 4.30865e-19 $X=0.405 $Y=0.2125
c45 66 VSS 0.0057844f $X=0.405 $Y=0.2
c46 65 VSS 4.01444e-19 $X=0.405 $Y=0.07
c47 64 VSS 0.00108941f $X=0.405 $Y=0.063
c48 63 VSS 8.62726e-19 $X=0.405 $Y=0.225
c49 61 VSS 0.00289269f $X=0.38 $Y=0.036
c50 60 VSS 3.40854e-19 $X=0.364 $Y=0.036
c51 59 VSS 0.00146362f $X=0.36 $Y=0.036
c52 58 VSS 0.0027713f $X=0.342 $Y=0.036
c53 57 VSS 9.5272e-19 $X=0.315 $Y=0.036
c54 56 VSS 0.00142296f $X=0.306 $Y=0.036
c55 55 VSS 0.00678169f $X=0.288 $Y=0.036
c56 54 VSS 0.00286574f $X=0.252 $Y=0.036
c57 53 VSS 0.0104492f $X=0.324 $Y=0.036
c58 49 VSS 0.00169362f $X=0.215 $Y=0.036
c59 48 VSS 0.00146362f $X=0.198 $Y=0.036
c60 47 VSS 0.00149782f $X=0.18 $Y=0.036
c61 46 VSS 0.0103752f $X=0.216 $Y=0.036
c62 43 VSS 0.00318678f $X=0.171 $Y=0.036
c63 42 VSS 0.00586463f $X=0.396 $Y=0.036
c64 41 VSS 6.41935e-19 $X=0.162 $Y=0.063
c65 39 VSS 0.00126924f $X=0.15 $Y=0.072
c66 38 VSS 1.4325e-20 $X=0.122 $Y=0.072
c67 37 VSS 1.44778e-19 $X=0.117 $Y=0.072
c68 36 VSS 0.0018601f $X=0.153 $Y=0.072
c69 35 VSS 2.28583e-19 $X=0.108 $Y=0.116
c70 34 VSS 6.20372e-19 $X=0.108 $Y=0.106
c71 33 VSS 2.29406e-19 $X=0.108 $Y=0.126
c72 30 VSS 0.00369079f $X=0.376 $Y=0.2025
c73 22 VSS 6.1012e-19 $X=0.341 $Y=0.0675
c74 17 VSS 6.55441e-19 $X=0.233 $Y=0.0675
c75 13 VSS 0.00128354f $X=0.135 $Y=0.135
c76 10 VSS 0.0612145f $X=0.135 $Y=0.0675
c77 5 VSS 0.00228311f $X=0.081 $Y=0.135
c78 2 VSS 0.0640029f $X=0.081 $Y=0.0675
r79 86 87 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.4005 $Y2=0.234
r80 85 87 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.234 $X2=0.4005 $Y2=0.234
r81 82 86 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.396 $Y2=0.234
r82 78 79 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.135 $X2=0.122 $Y2=0.135
r83 76 79 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.122 $Y2=0.135
r84 73 74 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.135 $X2=0.1035 $Y2=0.135
r85 72 78 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.135 $X2=0.117 $Y2=0.135
r86 72 74 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.135 $X2=0.1035 $Y2=0.135
r87 69 73 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.099 $Y2=0.135
r88 66 67 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.2 $X2=0.405 $Y2=0.2125
r89 65 66 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.07 $X2=0.405 $Y2=0.2
r90 64 65 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.063 $X2=0.405 $Y2=0.07
r91 63 85 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.234
r92 63 67 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.2125
r93 62 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.063
r94 60 61 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.364
+ $Y=0.036 $X2=0.38 $Y2=0.036
r95 59 60 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.036 $X2=0.364 $Y2=0.036
r96 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.36 $Y2=0.036
r97 56 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.036 $X2=0.315 $Y2=0.036
r98 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.306 $Y2=0.036
r99 54 55 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.036 $X2=0.288 $Y2=0.036
r100 52 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.342 $Y2=0.036
r101 52 57 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.315 $Y2=0.036
r102 52 53 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036
+ $X2=0.324 $Y2=0.036
r103 49 50 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.215
+ $Y=0.036 $X2=0.2155 $Y2=0.036
r104 48 49 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.215 $Y2=0.036
r105 47 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r106 45 54 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.252 $Y2=0.036
r107 45 50 0.0339506 $w=1.8e-08 $l=5e-10 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.2155 $Y2=0.036
r108 45 46 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036
+ $X2=0.216 $Y2=0.036
r109 43 47 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.036 $X2=0.18 $Y2=0.036
r110 42 62 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r111 42 61 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.38 $Y2=0.036
r112 40 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.045 $X2=0.171 $Y2=0.036
r113 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.045 $X2=0.162 $Y2=0.063
r114 38 39 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.122
+ $Y=0.072 $X2=0.15 $Y2=0.072
r115 37 38 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.117
+ $Y=0.072 $X2=0.122 $Y2=0.072
r116 36 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.153 $Y=0.072 $X2=0.162 $Y2=0.063
r117 36 39 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.153
+ $Y=0.072 $X2=0.15 $Y2=0.072
r118 34 35 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.106 $X2=0.108 $Y2=0.116
r119 33 72 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.126 $X2=0.108 $Y2=0.135
r120 33 35 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.126 $X2=0.108 $Y2=0.116
r121 32 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.108 $Y=0.081 $X2=0.117 $Y2=0.072
r122 32 34 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.081 $X2=0.108 $Y2=0.106
r123 30 82 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234
+ $X2=0.378 $Y2=0.234
r124 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.376 $Y2=0.2025
r125 26 53 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.324 $Y=0.0675 $X2=0.324 $Y2=0.036
r126 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.307 $Y=0.0675 $X2=0.324 $Y2=0.0675
r127 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.324 $Y2=0.0675
r128 21 46 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.216 $Y=0.0675 $X2=0.216 $Y2=0.036
r129 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r130 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r131 13 76 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r132 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r133 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r134 5 69 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r135 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r136 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_OR4X2_ASAP7_75T_R%D 2 5 7 11 VSS
c12 11 VSS 0.00473567f $X=0.189 $Y=0.132
c13 5 VSS 0.00107966f $X=0.189 $Y=0.135
c14 2 VSS 0.058708f $X=0.189 $Y=0.0675
r15 5 11 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r16 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r17 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_OR4X2_ASAP7_75T_R%C 2 5 7 12 VSS
c14 12 VSS 0.00782796f $X=0.243 $Y=0.132
c15 5 VSS 0.00165807f $X=0.243 $Y=0.135
c16 2 VSS 0.0598363f $X=0.243 $Y=0.0675
r17 5 12 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r18 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r19 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_OR4X2_ASAP7_75T_R%B 2 5 7 10 VSS
c13 10 VSS 0.00272832f $X=0.297 $Y=0.132
c14 5 VSS 0.00115441f $X=0.297 $Y=0.135
c15 2 VSS 0.060052f $X=0.297 $Y=0.0675
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r17 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r18 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_OR4X2_ASAP7_75T_R%A 2 5 7 10 VSS
c9 10 VSS 0.00227875f $X=0.351 $Y=0.132
c10 5 VSS 0.00229951f $X=0.351 $Y=0.135
c11 2 VSS 0.0641834f $X=0.351 $Y=0.0675
r12 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r13 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r14 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OR4X2_ASAP7_75T_R%Y 1 2 6 7 14 16 18 23 24 26 30 33 VSS
c17 33 VSS 0.00181175f $X=0.0875 $Y=0.234
c18 32 VSS 0.00725385f $X=0.067 $Y=0.234
c19 30 VSS 0.00377177f $X=0.108 $Y=0.234
c20 28 VSS 0.00320021f $X=0.027 $Y=0.234
c21 26 VSS 0.00273081f $X=0.099 $Y=0.036
c22 25 VSS 0.00725385f $X=0.067 $Y=0.036
c23 24 VSS 0.0101755f $X=0.108 $Y=0.036
c24 23 VSS 0.00252755f $X=0.108 $Y=0.036
c25 21 VSS 0.00320021f $X=0.027 $Y=0.036
c26 20 VSS 4.26553e-19 $X=0.018 $Y=0.216
c27 19 VSS 9.72017e-19 $X=0.018 $Y=0.207
c28 18 VSS 0.00260161f $X=0.018 $Y=0.189
c29 16 VSS 0.00320213f $X=0.018 $Y=0.126
c30 15 VSS 8.29409e-19 $X=0.018 $Y=0.063
c31 14 VSS 7.10225e-19 $X=0.018 $Y=0.132
c32 12 VSS 4.02856e-19 $X=0.018 $Y=0.225
c33 10 VSS 0.00865473f $X=0.108 $Y=0.2025
c34 6 VSS 7.01619e-19 $X=0.125 $Y=0.2025
c35 1 VSS 7.09533e-19 $X=0.125 $Y=0.0675
r36 32 33 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.067
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r37 30 33 1.39198 $w=1.8e-08 $l=2.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.0875 $Y2=0.234
r38 28 32 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.067 $Y2=0.234
r39 25 26 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.067
+ $Y=0.036 $X2=0.099 $Y2=0.036
r40 23 26 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.099 $Y2=0.036
r41 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r42 21 25 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.067 $Y2=0.036
r43 19 20 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.207 $X2=0.018 $Y2=0.216
r44 18 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.207
r45 17 18 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.189
r46 15 16 4.27778 $w=1.8e-08 $l=6.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.126
r47 14 17 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.132 $X2=0.018 $Y2=0.144
r48 14 16 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.132 $X2=0.018 $Y2=0.126
r49 12 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r50 12 20 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.216
r51 11 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r52 11 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r53 10 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r54 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r55 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r56 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r57 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r58 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends

.subckt PM_OR4X2_ASAP7_75T_R%9 1 2 VSS
c1 1 VSS 0.00214488f $X=0.233 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.199 $Y2=0.2025
.ends

.subckt PM_OR4X2_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00228146f $X=0.287 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.253 $Y2=0.2025
.ends

.subckt PM_OR4X2_ASAP7_75T_R%11 1 2 VSS
c0 1 VSS 0.00228146f $X=0.341 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.341
+ $Y=0.2025 $X2=0.307 $Y2=0.2025
.ends


* END of "./OR4x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt OR4x2_ASAP7_75t_R  VSS VDD D C B A Y
* 
* Y	Y
* A	A
* B	B
* C	C
* D	D
M0 N_Y_M0_d N_3_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_Y_M1_d N_3_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_3_M2_d N_D_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 VSS N_C_M3_g N_3_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 N_3_M4_d N_B_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 VSS N_A_M5_g N_3_M5_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_3_M6_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M7 N_Y_M7_d N_3_M7_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M8 N_9_M8_d N_D_M8_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M9 N_10_M9_d N_C_M9_g N_9_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 N_11_M10_d N_B_M10_g N_10_M10_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.287 $Y=0.162
M11 N_3_M11_d N_A_M11_g N_11_M11_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
*
* 
* .include "OR4x2_ASAP7_75t_R.pex.sp.OR4X2_ASAP7_75T_R.pxi"
* BEGIN of "./OR4x2_ASAP7_75t_R.pex.sp.OR4X2_ASAP7_75T_R.pxi"
* File: OR4x2_ASAP7_75t_R.pex.sp.OR4X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:01:55 2017
* 
x_PM_OR4X2_ASAP7_75T_R%3 N_3_M0_g N_3_c_24_p N_3_M6_g N_3_M1_g N_3_c_4_p
+ N_3_M7_g N_3_M3_s N_3_M2_d N_3_M5_s N_3_M4_d N_3_M11_d N_3_c_14_p N_3_c_29_p
+ N_3_c_5_p N_3_c_10_p N_3_c_26_p N_3_c_32_p N_3_c_28_p N_3_c_11_p N_3_c_3_p
+ N_3_c_15_p N_3_c_9_p N_3_c_13_p N_3_c_19_p N_3_c_23_p N_3_c_17_p N_3_c_25_p
+ N_3_c_7_p N_3_c_36_p N_3_c_18_p VSS PM_OR4X2_ASAP7_75T_R%3
x_PM_OR4X2_ASAP7_75T_R%D N_D_M2_g N_D_c_42_n N_D_M8_g D VSS
+ PM_OR4X2_ASAP7_75T_R%D
x_PM_OR4X2_ASAP7_75T_R%C N_C_M3_g N_C_c_57_n N_C_M9_g C VSS
+ PM_OR4X2_ASAP7_75T_R%C
x_PM_OR4X2_ASAP7_75T_R%B N_B_M4_g N_B_c_73_n N_B_M10_g B VSS
+ PM_OR4X2_ASAP7_75T_R%B
x_PM_OR4X2_ASAP7_75T_R%A N_A_M5_g N_A_c_85_n N_A_M11_g A VSS
+ PM_OR4X2_ASAP7_75T_R%A
x_PM_OR4X2_ASAP7_75T_R%Y N_Y_M1_d N_Y_M0_d N_Y_M7_d N_Y_M6_d Y N_Y_c_89_n
+ N_Y_c_102_n N_Y_c_90_n N_Y_c_92_n N_Y_c_97_n N_Y_c_99_n N_Y_c_100_n VSS
+ PM_OR4X2_ASAP7_75T_R%Y
x_PM_OR4X2_ASAP7_75T_R%9 N_9_M9_s N_9_M8_d VSS PM_OR4X2_ASAP7_75T_R%9
x_PM_OR4X2_ASAP7_75T_R%10 N_10_M10_s N_10_M9_d VSS PM_OR4X2_ASAP7_75T_R%10
x_PM_OR4X2_ASAP7_75T_R%11 N_11_M11_s N_11_M10_d VSS PM_OR4X2_ASAP7_75T_R%11
cc_1 N_3_M0_g N_D_M2_g 2.31381e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_3_M1_g N_D_M2_g 0.00284417f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_3_c_3_p N_D_M2_g 3.59101e-19 $X=0.198 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_4 N_3_c_4_p N_D_c_42_n 9.51968e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_5 N_3_c_5_p D 5.61145e-19 $X=0.108 $Y=0.116 $X2=0.189 $Y2=0.132
cc_6 N_3_c_3_p D 5.39549e-19 $X=0.198 $Y=0.036 $X2=0.189 $Y2=0.132
cc_7 N_3_c_7_p D 9.06205e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.132
cc_8 N_3_M1_g N_C_M3_g 2.31381e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_9 N_3_c_9_p N_C_M3_g 2.35421e-19 $X=0.252 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_10 N_3_c_10_p C 4.85889e-19 $X=0.153 $Y=0.072 $X2=0 $Y2=0
cc_11 N_3_c_11_p C 0.00210911f $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_12 N_3_c_9_p C 0.00373267f $X=0.252 $Y=0.036 $X2=0 $Y2=0
cc_13 N_3_c_13_p N_B_M4_g 2.57255e-19 $X=0.306 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_14 N_3_c_14_p B 4.68998e-19 $X=0.376 $Y=0.2025 $X2=0 $Y2=0
cc_15 N_3_c_15_p B 0.00114532f $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_16 N_3_c_13_p B 0.00123937f $X=0.306 $Y=0.036 $X2=0 $Y2=0
cc_17 N_3_c_17_p B 2.69891e-19 $X=0.405 $Y=0.2125 $X2=0 $Y2=0
cc_18 N_3_c_18_p B 4.44922e-19 $X=0.396 $Y=0.234 $X2=0 $Y2=0
cc_19 N_3_c_19_p N_A_M5_g 2.64924e-19 $X=0.36 $Y=0.036 $X2=0.189 $Y2=0.0675
cc_20 N_3_c_14_p A 0.0013295f $X=0.376 $Y=0.2025 $X2=0 $Y2=0
cc_21 N_3_c_15_p A 0.00114532f $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_22 N_3_c_19_p A 0.00125383f $X=0.36 $Y=0.036 $X2=0 $Y2=0
cc_23 N_3_c_23_p A 0.00499854f $X=0.405 $Y=0.2 $X2=0 $Y2=0
cc_24 N_3_c_24_p Y 2.59855e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_25 N_3_c_25_p Y 8.19699e-19 $X=0.099 $Y=0.135 $X2=0 $Y2=0
cc_26 N_3_c_26_p N_Y_c_89_n 0.00101189f $X=0.117 $Y=0.072 $X2=0.189 $Y2=0.135
cc_27 N_3_c_26_p N_Y_c_90_n 0.00178379f $X=0.117 $Y=0.072 $X2=0 $Y2=0
cc_28 N_3_c_28_p N_Y_c_90_n 9.64215e-19 $X=0.171 $Y=0.036 $X2=0 $Y2=0
cc_29 N_3_c_29_p N_Y_c_92_n 0.00145159f $X=0.108 $Y=0.106 $X2=0 $Y2=0
cc_30 N_3_c_5_p N_Y_c_92_n 6.24449e-19 $X=0.108 $Y=0.116 $X2=0 $Y2=0
cc_31 N_3_c_26_p N_Y_c_92_n 0.00118866f $X=0.117 $Y=0.072 $X2=0 $Y2=0
cc_32 N_3_c_32_p N_Y_c_92_n 5.48981e-19 $X=0.122 $Y=0.072 $X2=0 $Y2=0
cc_33 N_3_c_11_p N_Y_c_92_n 2.28909e-19 $X=0.216 $Y=0.036 $X2=0 $Y2=0
cc_34 N_3_M0_g N_Y_c_97_n 4.31632e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_3_c_25_p N_Y_c_97_n 5.89897e-19 $X=0.099 $Y=0.135 $X2=0 $Y2=0
cc_36 N_3_c_36_p N_Y_c_99_n 5.30962e-19 $X=0.117 $Y=0.135 $X2=0 $Y2=0
cc_37 N_3_M0_g N_Y_c_100_n 3.34515e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_38 N_3_c_25_p N_Y_c_100_n 5.30962e-19 $X=0.099 $Y=0.135 $X2=0 $Y2=0
cc_39 N_D_M2_g N_C_M3_g 0.00344695f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_40 N_D_c_42_n N_C_c_57_n 7.51247e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_41 D C 0.00489513f $X=0.189 $Y=0.132 $X2=0.135 $Y2=0.135
cc_42 N_D_M2_g N_B_M4_g 2.66145e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_43 D N_Y_c_102_n 2.67769e-19 $X=0.189 $Y=0.132 $X2=0.199 $Y2=0.0675
cc_44 N_C_M3_g N_B_M4_g 0.00327995f $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_45 N_C_c_57_n N_B_c_73_n 7.51247e-19 $X=0.243 $Y=0.135 $X2=0.081 $Y2=0.135
cc_46 C B 0.00749132f $X=0.243 $Y=0.132 $X2=0.135 $Y2=0.0675
cc_47 N_C_M3_g N_A_M5_g 2.71887e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_48 C N_Y_c_99_n 2.28048e-19 $X=0.243 $Y=0.132 $X2=0.376 $Y2=0.2025
cc_49 C N_9_M9_s 2.91005e-19 $X=0.243 $Y=0.132 $X2=0.081 $Y2=0.0675
cc_50 N_B_M4_g N_A_M5_g 0.00357042f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_51 N_B_c_73_n N_A_c_85_n 7.51046e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_52 B A 0.0057113f $X=0.297 $Y=0.132 $X2=0.135 $Y2=0.0675

* END of "./OR4x2_ASAP7_75t_R.pex.sp.OR4X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: OR5x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:02:17 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OR5x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./OR5x1_ASAP7_75t_R.pex.sp.pex"
* File: OR5x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:02:17 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OR5X1_ASAP7_75T_R%A 2 5 7 10 VSS
c10 10 VSS 0.00172694f $X=0.081 $Y=0.135
c11 5 VSS 0.00325747f $X=0.081 $Y=0.136
c12 2 VSS 0.0653596f $X=0.081 $Y=0.054
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.136 $X2=0.081
+ $Y2=0.136
r14 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.136 $X2=0.081 $Y2=0.2025
r15 2 5 307.213 $w=2e-08 $l=8.2e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.136
.ends

.subckt PM_OR5X1_ASAP7_75T_R%B 2 5 7 10 VSS
c12 10 VSS 0.0024522f $X=0.135 $Y=0.135
c13 5 VSS 0.0017107f $X=0.135 $Y=0.1355
c14 2 VSS 0.0604599f $X=0.135 $Y=0.054
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.136 $X2=0.135
+ $Y2=0.136
r16 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.2025
r17 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.1355
.ends

.subckt PM_OR5X1_ASAP7_75T_R%C 2 5 7 10 VSS
c11 10 VSS 0.00209947f $X=0.189 $Y=0.135
c12 5 VSS 0.00160244f $X=0.189 $Y=0.1355
c13 2 VSS 0.0597904f $X=0.189 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.136 $X2=0.189
+ $Y2=0.136
r15 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1355 $X2=0.189 $Y2=0.2025
r16 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.1355
.ends

.subckt PM_OR5X1_ASAP7_75T_R%D 2 5 7 10 VSS
c13 10 VSS 0.0024709f $X=0.243 $Y=0.135
c14 5 VSS 0.00160623f $X=0.243 $Y=0.1355
c15 2 VSS 0.059515f $X=0.243 $Y=0.054
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.136 $X2=0.243
+ $Y2=0.136
r17 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1355 $X2=0.243 $Y2=0.2025
r18 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.1355
.ends

.subckt PM_OR5X1_ASAP7_75T_R%E 2 5 7 10 VSS
c10 10 VSS 0.00305094f $X=0.297 $Y=0.135
c11 5 VSS 0.00162408f $X=0.297 $Y=0.1355
c12 2 VSS 0.0594813f $X=0.297 $Y=0.054
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.136 $X2=0.297
+ $Y2=0.136
r14 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.1355 $X2=0.297 $Y2=0.2025
r15 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.1355
.ends

.subckt PM_OR5X1_ASAP7_75T_R%8 2 5 7 9 12 14 15 18 19 20 23 24 27 32 33 43 45 51
+ 53 56 61 62 65 67 68 VSS
c32 68 VSS 1.69937e-19 $X=0.351 $Y=0.121
c33 67 VSS 9.91953e-19 $X=0.351 $Y=0.106
c34 65 VSS 2.89334e-19 $X=0.351 $Y=0.136
c35 62 VSS 1.69932e-19 $X=0.306 $Y=0.072
c36 61 VSS 0.00394258f $X=0.342 $Y=0.072
c37 60 VSS 8.65169e-19 $X=0.297 $Y=0.063
c38 56 VSS 0.00545273f $X=0.054 $Y=0.234
c39 54 VSS 0.00317163f $X=0.027 $Y=0.234
c40 53 VSS 0.00146362f $X=0.252 $Y=0.036
c41 52 VSS 0.00631462f $X=0.234 $Y=0.036
c42 51 VSS 0.00146362f $X=0.198 $Y=0.036
c43 50 VSS 0.00284382f $X=0.18 $Y=0.036
c44 46 VSS 9.64186e-19 $X=0.153 $Y=0.036
c45 45 VSS 0.00142296f $X=0.144 $Y=0.036
c46 44 VSS 0.00636214f $X=0.126 $Y=0.036
c47 43 VSS 0.00142296f $X=0.09 $Y=0.036
c48 42 VSS 1.68773e-19 $X=0.072 $Y=0.036
c49 41 VSS 0.00470185f $X=0.07 $Y=0.036
c50 34 VSS 0.0032477f $X=0.027 $Y=0.036
c51 33 VSS 0.0066498f $X=0.288 $Y=0.036
c52 32 VSS 0.00607891f $X=0.018 $Y=0.2
c53 31 VSS 9.13166e-19 $X=0.018 $Y=0.07
c54 30 VSS 0.00117262f $X=0.018 $Y=0.225
c55 27 VSS 0.00244555f $X=0.056 $Y=0.2025
c56 24 VSS 4.49354e-19 $X=0.071 $Y=0.2025
c57 23 VSS 0.00838562f $X=0.27 $Y=0.054
c58 19 VSS 5.3314e-19 $X=0.287 $Y=0.054
c59 18 VSS 0.00791982f $X=0.162 $Y=0.054
c60 14 VSS 5.3314e-19 $X=0.179 $Y=0.054
c61 12 VSS 0.00523518f $X=0.056 $Y=0.054
c62 9 VSS 2.53241e-19 $X=0.071 $Y=0.054
c63 5 VSS 0.00201427f $X=0.351 $Y=0.1355
c64 2 VSS 0.064696f $X=0.351 $Y=0.0675
r65 67 68 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.106 $X2=0.351 $Y2=0.121
r66 65 68 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.136 $X2=0.351 $Y2=0.121
r67 63 67 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.106
r68 61 63 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.072 $X2=0.351 $Y2=0.081
r69 61 62 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.072 $X2=0.306 $Y2=0.072
r70 60 62 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.297 $Y=0.063 $X2=0.306 $Y2=0.072
r71 59 60 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.063
r72 54 56 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.054 $Y2=0.234
r73 52 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r74 51 52 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.234 $Y2=0.036
r75 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r76 48 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.252 $Y2=0.036
r77 45 46 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.153 $Y2=0.036
r78 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r79 43 44 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.126 $Y2=0.036
r80 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r81 41 42 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.07
+ $Y=0.036 $X2=0.072 $Y2=0.036
r82 39 50 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r83 39 46 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.153 $Y2=0.036
r84 36 41 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.07 $Y2=0.036
r85 34 36 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.054 $Y2=0.036
r86 33 59 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r87 33 48 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.27 $Y2=0.036
r88 31 32 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.2
r89 30 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r90 30 32 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2
r91 29 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r92 29 31 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r93 27 56 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r94 24 27 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r95 23 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r96 20 23 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.054 $X2=0.27 $Y2=0.054
r97 19 23 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.054 $X2=0.27 $Y2=0.054
r98 18 39 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036 $X2=0.162
+ $Y2=0.036
r99 15 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.162 $Y2=0.054
r100 14 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.054 $X2=0.162 $Y2=0.054
r101 12 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r102 9 12 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r103 5 65 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.136 $X2=0.351
+ $Y2=0.136
r104 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.1355 $X2=0.351 $Y2=0.2025
r105 2 5 254.762 $w=2e-08 $l=6.8e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.1355
.ends

.subckt PM_OR5X1_ASAP7_75T_R%Y 1 6 13 14 20 28 30 32 VSS
c10 32 VSS 0.00163763f $X=0.405 $Y=0.1895
c11 30 VSS 0.00130271f $X=0.405 $Y=0.096
c12 29 VSS 8.85605e-19 $X=0.405 $Y=0.063
c13 28 VSS 0.00260206f $X=0.409 $Y=0.129
c14 26 VSS 0.00156079f $X=0.405 $Y=0.225
c15 20 VSS 0.00269153f $X=0.378 $Y=0.234
c16 18 VSS 0.00601235f $X=0.396 $Y=0.234
c17 14 VSS 0.00638782f $X=0.378 $Y=0.036
c18 13 VSS 0.00275846f $X=0.378 $Y=0.036
c19 11 VSS 0.00601314f $X=0.396 $Y=0.036
c20 9 VSS 0.00639685f $X=0.376 $Y=0.2025
c21 4 VSS 2.69461e-19 $X=0.376 $Y=0.0675
r22 31 32 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.154 $X2=0.405 $Y2=0.1895
r23 29 30 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.063 $X2=0.405 $Y2=0.096
r24 28 31 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.129 $X2=0.405 $Y2=0.154
r25 28 30 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.129 $X2=0.405 $Y2=0.096
r26 26 32 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.225 $X2=0.405 $Y2=0.1895
r27 25 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.045 $X2=0.405 $Y2=0.063
r28 18 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.234 $X2=0.405 $Y2=0.225
r29 18 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.234 $X2=0.378 $Y2=0.234
r30 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r31 11 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.036 $X2=0.405 $Y2=0.045
r32 11 13 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.378 $Y2=0.036
r33 9 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r34 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.2025 $X2=0.376 $Y2=0.2025
r35 4 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r36 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.0675 $X2=0.376 $Y2=0.0675
.ends

.subckt PM_OR5X1_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00228332f $X=0.125 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends

.subckt PM_OR5X1_ASAP7_75T_R%11 1 2 VSS
c0 1 VSS 0.00228332f $X=0.179 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends

.subckt PM_OR5X1_ASAP7_75T_R%12 1 2 VSS
c0 1 VSS 0.00228332f $X=0.233 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.199 $Y2=0.2025
.ends

.subckt PM_OR5X1_ASAP7_75T_R%13 1 2 VSS
c0 1 VSS 0.00228332f $X=0.287 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.253 $Y2=0.2025
.ends


* END of "./OR5x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt OR5x1_ASAP7_75t_R  VSS VDD A B C D E Y
* 
* Y	Y
* E	E
* D	D
* C	C
* B	B
* A	A
M0 VSS N_A_M0_g N_8_M0_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_8_M1_d N_B_M1_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_C_M2_g N_8_M2_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 N_8_M3_d N_D_M3_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 VSS N_E_M4_g N_8_M4_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_8_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_10_M6_d N_A_M6_g N_8_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M7 N_11_M7_d N_B_M7_g N_10_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M8 N_12_M8_d N_C_M8_g N_11_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M9 N_13_M9_d N_D_M9_g N_12_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M10 VDD N_E_M10_g N_13_M10_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 N_Y_M11_d N_8_M11_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
*
* 
* .include "OR5x1_ASAP7_75t_R.pex.sp.OR5X1_ASAP7_75T_R.pxi"
* BEGIN of "./OR5x1_ASAP7_75t_R.pex.sp.OR5X1_ASAP7_75T_R.pxi"
* File: OR5x1_ASAP7_75t_R.pex.sp.OR5X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:02:17 2017
* 
x_PM_OR5X1_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M6_g A VSS
+ PM_OR5X1_ASAP7_75T_R%A
x_PM_OR5X1_ASAP7_75T_R%B N_B_M1_g N_B_c_12_n N_B_M7_g B VSS
+ PM_OR5X1_ASAP7_75T_R%B
x_PM_OR5X1_ASAP7_75T_R%C N_C_M2_g N_C_c_25_n N_C_M8_g C VSS
+ PM_OR5X1_ASAP7_75T_R%C
x_PM_OR5X1_ASAP7_75T_R%D N_D_M3_g N_D_c_36_n N_D_M9_g D VSS
+ PM_OR5X1_ASAP7_75T_R%D
x_PM_OR5X1_ASAP7_75T_R%E N_E_M4_g N_E_c_49_n N_E_M10_g E VSS
+ PM_OR5X1_ASAP7_75T_R%E
x_PM_OR5X1_ASAP7_75T_R%8 N_8_M5_g N_8_c_78_n N_8_M11_g N_8_M0_s N_8_c_57_n
+ N_8_M2_s N_8_M1_d N_8_c_63_n N_8_M4_s N_8_M3_d N_8_c_72_n N_8_M6_s N_8_c_58_n
+ N_8_c_60_n N_8_c_82_p N_8_c_61_n N_8_c_65_n N_8_c_69_n N_8_c_73_n N_8_c_67_n
+ N_8_c_83_p N_8_c_75_n N_8_c_86_p N_8_c_76_n N_8_c_80_n VSS
+ PM_OR5X1_ASAP7_75T_R%8
x_PM_OR5X1_ASAP7_75T_R%Y N_Y_M5_d N_Y_M11_d N_Y_c_91_n N_Y_c_94_n N_Y_c_89_n Y
+ N_Y_c_98_n N_Y_c_90_n VSS PM_OR5X1_ASAP7_75T_R%Y
x_PM_OR5X1_ASAP7_75T_R%10 N_10_M7_s N_10_M6_d VSS PM_OR5X1_ASAP7_75T_R%10
x_PM_OR5X1_ASAP7_75T_R%11 N_11_M8_s N_11_M7_d VSS PM_OR5X1_ASAP7_75T_R%11
x_PM_OR5X1_ASAP7_75T_R%12 N_12_M9_s N_12_M8_d VSS PM_OR5X1_ASAP7_75T_R%12
x_PM_OR5X1_ASAP7_75T_R%13 N_13_M10_s N_13_M9_d VSS PM_OR5X1_ASAP7_75T_R%13
cc_1 N_A_M0_g N_B_M1_g 0.00333077f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A_c_2_p N_B_c_12_n 7.98811e-19 $X=0.081 $Y=0.136 $X2=0.135 $Y2=0.1355
cc_3 A B 0.00621434f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A_M0_g N_C_M2_g 2.71887e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 A N_8_c_57_n 3.52002e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.136
cc_6 N_A_c_2_p N_8_c_58_n 3.06446e-19 $X=0.081 $Y=0.136 $X2=0 $Y2=0
cc_7 A N_8_c_58_n 0.00134508f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_8 A N_8_c_60_n 0.00436697f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_A_M0_g N_8_c_61_n 2.57864e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_10 A N_8_c_61_n 0.00123648f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 N_B_M1_g N_C_M2_g 0.00357042f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_12 N_B_c_12_n N_C_c_25_n 7.92653e-19 $X=0.135 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_13 B C 0.00817592f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 N_B_M1_g N_D_M3_g 2.71887e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_15 B N_8_c_63_n 3.31541e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_16 B N_8_c_58_n 5.56013e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_17 N_B_M1_g N_8_c_65_n 2.57565e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_18 B N_8_c_65_n 0.00123952f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_19 B N_8_c_67_n 4.64233e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_20 N_C_M2_g N_D_M3_g 0.00327995f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_21 N_C_c_25_n N_D_c_36_n 7.90494e-19 $X=0.189 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_22 C D 0.00817682f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 N_C_M2_g N_E_M4_g 2.66145e-19 $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_24 C N_8_c_63_n 3.31541e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_25 N_C_M2_g N_8_c_69_n 2.64924e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_26 C N_8_c_69_n 0.00125705f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_27 N_D_M3_g N_E_M4_g 0.00344695f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_28 N_D_c_36_n N_E_c_49_n 7.90494e-19 $X=0.243 $Y=0.1355 $X2=0.135 $Y2=0.1355
cc_29 D E 0.00646431f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_30 N_D_M3_g N_8_M5_g 2.31381e-19 $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_31 D N_8_c_72_n 3.24828e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_32 N_D_M3_g N_8_c_73_n 2.64924e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_33 D N_8_c_73_n 0.00125705f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_34 D N_8_c_75_n 4.59663e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_35 D N_8_c_76_n 2.69033e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_36 N_E_M4_g N_8_M5_g 0.00284417f $X=0.297 $Y=0.054 $X2=0.189 $Y2=0.054
cc_37 N_E_c_49_n N_8_c_78_n 8.31912e-19 $X=0.297 $Y=0.1355 $X2=0.189 $Y2=0.1355
cc_38 E N_8_c_75_n 0.00135016f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_39 E N_8_c_80_n 0.00215339f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_40 E N_Y_c_89_n 3.55123e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_41 E N_Y_c_90_n 4.73275e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_42 N_8_M5_g N_Y_c_91_n 2.56972e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.136
cc_43 N_8_c_82_p N_Y_c_91_n 5.2369e-19 $X=0.288 $Y=0.036 $X2=0.081 $Y2=0.136
cc_44 N_8_c_83_p N_Y_c_91_n 0.00100131f $X=0.342 $Y=0.072 $X2=0.081 $Y2=0.136
cc_45 N_8_c_83_p N_Y_c_94_n 0.00135705f $X=0.342 $Y=0.072 $X2=0 $Y2=0
cc_46 N_8_M5_g N_Y_c_89_n 3.02028e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_8_c_86_p N_Y_c_89_n 2.49025e-19 $X=0.351 $Y=0.136 $X2=0 $Y2=0
cc_48 N_8_c_80_n Y 0.00186022f $X=0.351 $Y=0.121 $X2=0 $Y2=0
cc_49 N_8_c_83_p N_Y_c_98_n 0.00186022f $X=0.342 $Y=0.072 $X2=0 $Y2=0

* END of "./OR5x1_ASAP7_75t_R.pex.sp.OR5X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: OR5x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:02:40 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "OR5x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./OR5x2_ASAP7_75t_R.pex.sp.pex"
* File: OR5x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:02:40 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_OR5X2_ASAP7_75T_R%A 2 5 7 10 VSS
c10 10 VSS 0.00172694f $X=0.081 $Y=0.135
c11 5 VSS 0.00325747f $X=0.081 $Y=0.136
c12 2 VSS 0.0653596f $X=0.081 $Y=0.054
r13 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.136 $X2=0.081
+ $Y2=0.136
r14 5 7 249.142 $w=2e-08 $l=6.65e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.136 $X2=0.081 $Y2=0.2025
r15 2 5 307.213 $w=2e-08 $l=8.2e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.136
.ends

.subckt PM_OR5X2_ASAP7_75T_R%B 2 5 7 10 VSS
c12 10 VSS 0.0024522f $X=0.135 $Y=0.135
c13 5 VSS 0.0017107f $X=0.135 $Y=0.1355
c14 2 VSS 0.0604599f $X=0.135 $Y=0.054
r15 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.136 $X2=0.135
+ $Y2=0.136
r16 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.1355 $X2=0.135 $Y2=0.2025
r17 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.1355
.ends

.subckt PM_OR5X2_ASAP7_75T_R%C 2 5 7 10 VSS
c11 10 VSS 0.00209947f $X=0.189 $Y=0.135
c12 5 VSS 0.00160244f $X=0.189 $Y=0.1355
c13 2 VSS 0.0597904f $X=0.189 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.136 $X2=0.189
+ $Y2=0.136
r15 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.1355 $X2=0.189 $Y2=0.2025
r16 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.054 $X2=0.189 $Y2=0.1355
.ends

.subckt PM_OR5X2_ASAP7_75T_R%D 2 5 7 10 VSS
c13 10 VSS 0.00246323f $X=0.243 $Y=0.135
c14 5 VSS 0.00160828f $X=0.243 $Y=0.1355
c15 2 VSS 0.059515f $X=0.243 $Y=0.054
r16 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.136 $X2=0.243
+ $Y2=0.136
r17 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.1355 $X2=0.243 $Y2=0.2025
r18 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.054 $X2=0.243 $Y2=0.1355
.ends

.subckt PM_OR5X2_ASAP7_75T_R%E 2 5 7 10 VSS
c11 10 VSS 0.00347535f $X=0.297 $Y=0.135
c12 5 VSS 0.00152014f $X=0.297 $Y=0.1355
c13 2 VSS 0.0587069f $X=0.297 $Y=0.054
r14 5 10 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.136 $X2=0.297
+ $Y2=0.136
r15 5 7 251.016 $w=2e-08 $l=6.7e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.1355 $X2=0.297 $Y2=0.2025
r16 2 5 305.34 $w=2e-08 $l=8.15e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.054 $X2=0.297 $Y2=0.1355
.ends

.subckt PM_OR5X2_ASAP7_75T_R%8 2 7 10 13 15 17 20 22 23 26 27 28 31 32 35 40 41
+ 51 53 59 61 64 69 70 75 76 VSS
c40 76 VSS 1.76122e-19 $X=0.351 $Y=0.121
c41 75 VSS 9.91953e-19 $X=0.351 $Y=0.106
c42 73 VSS 4.38495e-19 $X=0.351 $Y=0.136
c43 70 VSS 1.69932e-19 $X=0.306 $Y=0.072
c44 69 VSS 0.00373357f $X=0.342 $Y=0.072
c45 68 VSS 8.65169e-19 $X=0.297 $Y=0.063
c46 64 VSS 0.00545273f $X=0.054 $Y=0.234
c47 62 VSS 0.00317163f $X=0.027 $Y=0.234
c48 61 VSS 0.00146362f $X=0.252 $Y=0.036
c49 60 VSS 0.00631462f $X=0.234 $Y=0.036
c50 59 VSS 0.00146362f $X=0.198 $Y=0.036
c51 58 VSS 0.00284382f $X=0.18 $Y=0.036
c52 54 VSS 9.64186e-19 $X=0.153 $Y=0.036
c53 53 VSS 0.00142296f $X=0.144 $Y=0.036
c54 52 VSS 0.00636214f $X=0.126 $Y=0.036
c55 51 VSS 0.00142296f $X=0.09 $Y=0.036
c56 50 VSS 1.68773e-19 $X=0.072 $Y=0.036
c57 49 VSS 0.00470185f $X=0.07 $Y=0.036
c58 42 VSS 0.0032477f $X=0.027 $Y=0.036
c59 41 VSS 0.00660869f $X=0.288 $Y=0.036
c60 40 VSS 0.00607891f $X=0.018 $Y=0.2
c61 39 VSS 9.13166e-19 $X=0.018 $Y=0.07
c62 38 VSS 0.00117262f $X=0.018 $Y=0.225
c63 35 VSS 0.00244555f $X=0.056 $Y=0.2025
c64 32 VSS 4.49354e-19 $X=0.071 $Y=0.2025
c65 31 VSS 0.00836246f $X=0.27 $Y=0.054
c66 27 VSS 5.3314e-19 $X=0.287 $Y=0.054
c67 26 VSS 0.00791982f $X=0.162 $Y=0.054
c68 22 VSS 5.3314e-19 $X=0.179 $Y=0.054
c69 20 VSS 0.00523518f $X=0.056 $Y=0.054
c70 17 VSS 2.53241e-19 $X=0.071 $Y=0.054
c71 13 VSS 0.0040976f $X=0.405 $Y=0.135
c72 10 VSS 0.0639847f $X=0.405 $Y=0.0675
c73 2 VSS 0.060828f $X=0.351 $Y=0.0675
r74 75 76 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.106 $X2=0.351 $Y2=0.121
r75 73 76 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.136 $X2=0.351 $Y2=0.121
r76 71 75 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.106
r77 69 71 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.072 $X2=0.351 $Y2=0.081
r78 69 70 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.072 $X2=0.306 $Y2=0.072
r79 68 70 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.297 $Y=0.063 $X2=0.306 $Y2=0.072
r80 67 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.045 $X2=0.297 $Y2=0.063
r81 62 64 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.054 $Y2=0.234
r82 60 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.036 $X2=0.252 $Y2=0.036
r83 59 60 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.036 $X2=0.234 $Y2=0.036
r84 58 59 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.198 $Y2=0.036
r85 56 61 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.252 $Y2=0.036
r86 53 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.153 $Y2=0.036
r87 52 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r88 51 52 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.126 $Y2=0.036
r89 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r90 49 50 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.07
+ $Y=0.036 $X2=0.072 $Y2=0.036
r91 47 58 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r92 47 54 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.153 $Y2=0.036
r93 44 49 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.07 $Y2=0.036
r94 42 44 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.054 $Y2=0.036
r95 41 67 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.288 $Y=0.036 $X2=0.297 $Y2=0.045
r96 41 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.036 $X2=0.27 $Y2=0.036
r97 39 40 8.82716 $w=1.8e-08 $l=1.3e-07 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.07 $X2=0.018 $Y2=0.2
r98 38 62 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r99 38 40 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.2
r100 37 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r101 37 39 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.07
r102 35 64 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r103 32 35 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r104 31 56 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r105 28 31 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.054 $X2=0.27 $Y2=0.054
r106 27 31 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.054 $X2=0.27 $Y2=0.054
r107 26 47 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.162 $Y=0.036
+ $X2=0.162 $Y2=0.036
r108 23 26 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.054 $X2=0.162 $Y2=0.054
r109 22 26 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.179 $Y=0.054 $X2=0.162 $Y2=0.054
r110 20 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036
+ $X2=0.054 $Y2=0.036
r111 17 20 11.1111 $w=5.4e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.054 $X2=0.056 $Y2=0.054
r112 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r113 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r114 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.405 $Y2=0.135
r115 5 73 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.136 $X2=0.351
+ $Y2=0.136
r116 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r117 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_OR5X2_ASAP7_75T_R%Y 1 2 6 7 10 11 13 14 18 26 28 30 VSS
c17 30 VSS 0.0022158f $X=0.459 $Y=0.1895
c18 28 VSS 0.00230667f $X=0.459 $Y=0.10525
c19 27 VSS 8.85605e-19 $X=0.459 $Y=0.063
c20 26 VSS 0.00238564f $X=0.459 $Y=0.1475
c21 24 VSS 0.00189369f $X=0.459 $Y=0.225
c22 18 VSS 0.0146644f $X=0.45 $Y=0.234
c23 14 VSS 0.0104099f $X=0.378 $Y=0.036
c24 13 VSS 0.00285686f $X=0.378 $Y=0.036
c25 11 VSS 0.0135753f $X=0.45 $Y=0.036
c26 10 VSS 0.00904301f $X=0.378 $Y=0.2025
c27 6 VSS 5.72268e-19 $X=0.395 $Y=0.2025
c28 1 VSS 5.25448e-19 $X=0.395 $Y=0.0675
r29 29 30 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.154 $X2=0.459 $Y2=0.1895
r30 27 28 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.063 $X2=0.459 $Y2=0.10525
r31 26 29 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.1475 $X2=0.459 $Y2=0.154
r32 26 28 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.1475 $X2=0.459 $Y2=0.10525
r33 24 30 2.41049 $w=1.8e-08 $l=3.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.1895
r34 23 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.063
r35 18 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r36 18 20 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.378 $Y2=0.234
r37 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r38 11 23 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r39 11 13 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.378 $Y2=0.036
r40 10 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r41 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r42 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r43 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r44 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.0675 $X2=0.378 $Y2=0.0675
r45 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.378 $Y2=0.0675
.ends

.subckt PM_OR5X2_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00228332f $X=0.125 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends

.subckt PM_OR5X2_ASAP7_75T_R%11 1 2 VSS
c0 1 VSS 0.00228332f $X=0.179 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends

.subckt PM_OR5X2_ASAP7_75T_R%12 1 2 VSS
c0 1 VSS 0.00228332f $X=0.233 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.199 $Y2=0.2025
.ends

.subckt PM_OR5X2_ASAP7_75T_R%13 1 2 VSS
c0 1 VSS 0.00228332f $X=0.287 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.253 $Y2=0.2025
.ends


* END of "./OR5x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt OR5x2_ASAP7_75t_R  VSS VDD A B C D E Y
* 
* Y	Y
* E	E
* D	D
* C	C
* B	B
* A	A
M0 VSS N_A_M0_g N_8_M0_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 N_8_M1_d N_B_M1_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 VSS N_C_M2_g N_8_M2_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.179 $Y=0.027
M3 N_8_M3_d N_D_M3_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.233 $Y=0.027
M4 VSS N_E_M4_g N_8_M4_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_8_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_8_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_10_M7_d N_A_M7_g N_8_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M8 N_11_M8_d N_B_M8_g N_10_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M9 N_12_M9_d N_C_M9_g N_11_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M10 N_13_M10_d N_D_M10_g N_12_M10_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M11 VDD N_E_M11_g N_13_M11_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M12 N_Y_M12_d N_8_M12_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M13 N_Y_M13_d N_8_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
*
* 
* .include "OR5x2_ASAP7_75t_R.pex.sp.OR5X2_ASAP7_75T_R.pxi"
* BEGIN of "./OR5x2_ASAP7_75t_R.pex.sp.OR5X2_ASAP7_75T_R.pxi"
* File: OR5x2_ASAP7_75t_R.pex.sp.OR5X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:02:40 2017
* 
x_PM_OR5X2_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M7_g A VSS
+ PM_OR5X2_ASAP7_75T_R%A
x_PM_OR5X2_ASAP7_75T_R%B N_B_M1_g N_B_c_12_n N_B_M8_g B VSS
+ PM_OR5X2_ASAP7_75T_R%B
x_PM_OR5X2_ASAP7_75T_R%C N_C_M2_g N_C_c_25_n N_C_M9_g C VSS
+ PM_OR5X2_ASAP7_75T_R%C
x_PM_OR5X2_ASAP7_75T_R%D N_D_M3_g N_D_c_36_n N_D_M10_g D VSS
+ PM_OR5X2_ASAP7_75T_R%D
x_PM_OR5X2_ASAP7_75T_R%E N_E_M4_g N_E_c_49_n N_E_M11_g E VSS
+ PM_OR5X2_ASAP7_75T_R%E
x_PM_OR5X2_ASAP7_75T_R%8 N_8_M5_g N_8_M12_g N_8_M6_g N_8_c_80_n N_8_M13_g
+ N_8_M0_s N_8_c_58_n N_8_M2_s N_8_M1_d N_8_c_64_n N_8_M4_s N_8_M3_d N_8_c_73_n
+ N_8_M7_s N_8_c_59_n N_8_c_61_n N_8_c_89_p N_8_c_62_n N_8_c_66_n N_8_c_70_n
+ N_8_c_74_n N_8_c_68_n N_8_c_90_p N_8_c_76_n N_8_c_77_n N_8_c_82_n VSS
+ PM_OR5X2_ASAP7_75T_R%8
x_PM_OR5X2_ASAP7_75T_R%Y N_Y_M6_d N_Y_M5_d N_Y_M13_d N_Y_M12_d N_Y_c_102_n
+ N_Y_c_103_n N_Y_c_104_n N_Y_c_108_n N_Y_c_98_n Y N_Y_c_114_n N_Y_c_99_n VSS
+ PM_OR5X2_ASAP7_75T_R%Y
x_PM_OR5X2_ASAP7_75T_R%10 N_10_M8_s N_10_M7_d VSS PM_OR5X2_ASAP7_75T_R%10
x_PM_OR5X2_ASAP7_75T_R%11 N_11_M9_s N_11_M8_d VSS PM_OR5X2_ASAP7_75T_R%11
x_PM_OR5X2_ASAP7_75T_R%12 N_12_M10_s N_12_M9_d VSS PM_OR5X2_ASAP7_75T_R%12
x_PM_OR5X2_ASAP7_75T_R%13 N_13_M11_s N_13_M10_d VSS PM_OR5X2_ASAP7_75T_R%13
cc_1 N_A_M0_g N_B_M1_g 0.00333077f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A_c_2_p N_B_c_12_n 7.98811e-19 $X=0.081 $Y=0.136 $X2=0.135 $Y2=0.1355
cc_3 A B 0.00621434f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_A_M0_g N_C_M2_g 2.71887e-19 $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_5 A N_8_c_58_n 3.52002e-19 $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_6 N_A_c_2_p N_8_c_59_n 3.06446e-19 $X=0.081 $Y=0.136 $X2=0 $Y2=0
cc_7 A N_8_c_59_n 0.00134508f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_8 A N_8_c_61_n 0.00436697f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_9 N_A_M0_g N_8_c_62_n 2.57864e-19 $X=0.081 $Y=0.054 $X2=0 $Y2=0
cc_10 A N_8_c_62_n 0.00123648f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_11 N_B_M1_g N_C_M2_g 0.00357042f $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_12 N_B_c_12_n N_C_c_25_n 7.92653e-19 $X=0.135 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_13 B C 0.00817592f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_14 N_B_M1_g N_D_M3_g 2.71887e-19 $X=0.135 $Y=0.054 $X2=0.081 $Y2=0.054
cc_15 B N_8_c_64_n 3.31541e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_16 B N_8_c_59_n 5.56013e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_17 N_B_M1_g N_8_c_66_n 2.57565e-19 $X=0.135 $Y=0.054 $X2=0 $Y2=0
cc_18 B N_8_c_66_n 0.00123952f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_19 B N_8_c_68_n 4.64233e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_20 N_C_M2_g N_D_M3_g 0.00327995f $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_21 N_C_c_25_n N_D_c_36_n 7.90494e-19 $X=0.189 $Y=0.1355 $X2=0.081 $Y2=0.136
cc_22 C D 0.00817682f $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 N_C_M2_g N_E_M4_g 2.66145e-19 $X=0.189 $Y=0.054 $X2=0.081 $Y2=0.054
cc_24 C N_8_c_64_n 3.31541e-19 $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_25 N_C_M2_g N_8_c_70_n 2.64924e-19 $X=0.189 $Y=0.054 $X2=0 $Y2=0
cc_26 C N_8_c_70_n 0.00125705f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_27 N_D_M3_g N_E_M4_g 0.00344695f $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_28 N_D_c_36_n N_E_c_49_n 7.90494e-19 $X=0.243 $Y=0.1355 $X2=0.135 $Y2=0.1355
cc_29 D E 0.00646361f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_30 N_D_M3_g N_8_M5_g 2.31381e-19 $X=0.243 $Y=0.054 $X2=0.135 $Y2=0.054
cc_31 D N_8_c_73_n 3.24828e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_32 N_D_M3_g N_8_c_74_n 2.64924e-19 $X=0.243 $Y=0.054 $X2=0 $Y2=0
cc_33 D N_8_c_74_n 0.00125705f $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_34 D N_8_c_76_n 4.59663e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_35 D N_8_c_77_n 2.69033e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_36 N_E_M4_g N_8_M5_g 0.00284417f $X=0.297 $Y=0.054 $X2=0.189 $Y2=0.054
cc_37 N_E_M4_g N_8_M6_g 2.31381e-19 $X=0.297 $Y=0.054 $X2=0.189 $Y2=0.135
cc_38 N_E_c_49_n N_8_c_80_n 8.36511e-19 $X=0.297 $Y=0.1355 $X2=0.189 $Y2=0.136
cc_39 E N_8_c_76_n 0.00135016f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_40 E N_8_c_82_n 0.00213556f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_41 E N_Y_c_98_n 2.63055e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_42 E N_Y_c_99_n 2.15095e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_43 N_8_c_80_n N_Y_M6_d 3.80663e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.054
cc_44 N_8_c_80_n N_Y_M13_d 3.80663e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_45 N_8_c_80_n N_Y_c_102_n 8.00061e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_46 N_8_M6_g N_Y_c_103_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_8_M5_g N_Y_c_104_n 2.30014e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.136
cc_48 N_8_c_80_n N_Y_c_104_n 6.10804e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.136
cc_49 N_8_c_89_p N_Y_c_104_n 6.57712e-19 $X=0.288 $Y=0.036 $X2=0.081 $Y2=0.136
cc_50 N_8_c_90_p N_Y_c_104_n 0.0015537f $X=0.342 $Y=0.072 $X2=0.081 $Y2=0.136
cc_51 N_8_c_80_n N_Y_c_108_n 8.00061e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_52 N_8_c_90_p N_Y_c_108_n 0.00157502f $X=0.342 $Y=0.072 $X2=0 $Y2=0
cc_53 N_8_M6_g N_Y_c_98_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_54 N_8_c_80_n N_Y_c_98_n 5.51214e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_55 N_8_c_80_n Y 4.10099e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_56 N_8_c_82_n Y 5.62507e-19 $X=0.351 $Y=0.121 $X2=0 $Y2=0
cc_57 N_8_c_90_p N_Y_c_114_n 5.62507e-19 $X=0.342 $Y=0.072 $X2=0 $Y2=0

* END of "./OR5x2_ASAP7_75t_R.pex.sp.OR5X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: XOR2x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:07:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "XOR2x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./XOR2x1_ASAP7_75t_R.pex.sp.pex"
* File: XOR2x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:07:55 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_XOR2X1_ASAP7_75T_R%A 2 5 7 10 13 15 18 21 23 37 41 45 46 47 48 49 50
+ 52 53 54 56 59 60 61 63 66 72 73 84 91 VSS
c65 91 VSS 5.91166e-19 $X=0.513 $Y=0.169
c66 84 VSS 2.50262e-19 $X=0.513 $Y=0.135
c67 73 VSS 0.0018565f $X=0.513 $Y=0.189
c68 72 VSS 0.00559832f $X=0.513 $Y=0.189
c69 66 VSS 0.00766534f $X=0.018 $Y=0.135
c70 63 VSS 6.41874e-19 $X=0.351 $Y=0.135
c71 61 VSS 1.40425e-19 $X=0.323 $Y=0.135
c72 60 VSS 0.00120624f $X=0.314 $Y=0.175
c73 59 VSS 2.5887e-19 $X=0.314 $Y=0.149
c74 58 VSS 0.00219751f $X=0.314 $Y=0.185
c75 56 VSS 1.57364e-19 $X=0.2805 $Y=0.194
c76 55 VSS 0.00137179f $X=0.256 $Y=0.194
c77 54 VSS 3.88371e-19 $X=0.231 $Y=0.194
c78 53 VSS 1.68167e-19 $X=0.305 $Y=0.194
c79 52 VSS 2.80979e-20 $X=0.222 $Y=0.225
c80 50 VSS 0.00102062f $X=0.2025 $Y=0.234
c81 49 VSS 0.00132447f $X=0.192 $Y=0.234
c82 48 VSS 0.00269371f $X=0.174 $Y=0.234
c83 47 VSS 0.00142972f $X=0.144 $Y=0.234
c84 46 VSS 0.00192708f $X=0.126 $Y=0.234
c85 45 VSS 0.00156636f $X=0.107 $Y=0.234
c86 44 VSS 0.00122076f $X=0.092 $Y=0.234
c87 43 VSS 0.0075732f $X=0.078 $Y=0.234
c88 42 VSS 0.00323226f $X=0.027 $Y=0.234
c89 41 VSS 0.00322347f $X=0.213 $Y=0.234
c90 37 VSS 0.00238557f $X=0.06 $Y=0.134
c91 34 VSS 0.00210073f $X=0.018 $Y=0.188
c92 33 VSS 1.95142e-19 $X=0.018 $Y=0.149
c93 32 VSS 0.00169007f $X=0.018 $Y=0.225
c94 21 VSS 0.00101384f $X=0.513 $Y=0.135
c95 18 VSS 0.0608664f $X=0.513 $Y=0.0675
c96 13 VSS 0.0014355f $X=0.351 $Y=0.135
c97 10 VSS 0.0612409f $X=0.351 $Y=0.0675
c98 5 VSS 0.0062617f $X=0.081 $Y=0.135
c99 2 VSS 0.0638905f $X=0.081 $Y=0.0675
r100 90 91 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.149 $X2=0.513 $Y2=0.169
r101 84 90 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.149
r102 73 91 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.189 $X2=0.513 $Y2=0.169
r103 72 73 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.189 $X2=0.513
+ $Y2=0.189
r104 68 72 13.5123 $w=1.8e-08 $l=1.99e-07 $layer=M2 $thickness=3.6e-08 $X=0.314
+ $Y=0.189 $X2=0.513 $Y2=0.189
r105 68 69 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.314 $Y=0.189 $X2=0.314
+ $Y2=0.189
r106 61 63 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.323
+ $Y=0.135 $X2=0.351 $Y2=0.135
r107 59 60 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.314
+ $Y=0.149 $X2=0.314 $Y2=0.175
r108 58 69 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.314
+ $Y=0.185 $X2=0.314 $Y2=0.194
r109 58 60 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.314
+ $Y=0.185 $X2=0.314 $Y2=0.175
r110 57 61 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.314 $Y=0.144 $X2=0.323 $Y2=0.135
r111 57 59 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.314
+ $Y=0.144 $X2=0.314 $Y2=0.149
r112 55 56 1.66358 $w=1.8e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.194 $X2=0.2805 $Y2=0.194
r113 54 55 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.231
+ $Y=0.194 $X2=0.256 $Y2=0.194
r114 53 69 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.305
+ $Y=0.194 $X2=0.314 $Y2=0.194
r115 53 56 1.66358 $w=1.8e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.305
+ $Y=0.194 $X2=0.2805 $Y2=0.194
r116 51 54 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.222 $Y=0.203 $X2=0.231 $Y2=0.194
r117 51 52 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.222
+ $Y=0.203 $X2=0.222 $Y2=0.225
r118 49 50 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.192
+ $Y=0.234 $X2=0.2025 $Y2=0.234
r119 48 49 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.174
+ $Y=0.234 $X2=0.192 $Y2=0.234
r120 47 48 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.174 $Y2=0.234
r121 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.144 $Y2=0.234
r122 45 46 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.234 $X2=0.126 $Y2=0.234
r123 44 45 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.092
+ $Y=0.234 $X2=0.107 $Y2=0.234
r124 43 44 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.234 $X2=0.092 $Y2=0.234
r125 42 43 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.078 $Y2=0.234
r126 41 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.213 $Y=0.234 $X2=0.222 $Y2=0.225
r127 41 50 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.213
+ $Y=0.234 $X2=0.2025 $Y2=0.234
r128 37 39 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r129 35 66 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r130 35 37 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.06 $Y2=0.135
r131 33 34 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.149 $X2=0.018 $Y2=0.188
r132 32 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r133 32 34 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.188
r134 31 66 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r135 31 33 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.149
r136 21 84 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r137 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r138 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r139 13 63 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r140 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r141 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r142 5 39 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r143 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r144 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_XOR2X1_ASAP7_75T_R%B 2 7 10 13 15 18 21 23 33 36 38 39 40 41 45 51 56
+ 57 62 63 VSS
c65 63 VSS 1.32738e-19 $X=0.567 $Y=0.1265
c66 62 VSS 7.53013e-19 $X=0.567 $Y=0.118
c67 57 VSS 7.29302e-20 $X=0.135 $Y=0.1305
c68 56 VSS 0.00125411f $X=0.135 $Y=0.126
c69 51 VSS 8.08201e-20 $X=0.567 $Y=0.135
c70 45 VSS 1.6751e-19 $X=0.135 $Y=0.135
c71 41 VSS 0.00555131f $X=0.527 $Y=0.081
c72 40 VSS 0.00750485f $X=0.298 $Y=0.081
c73 39 VSS 6.93547e-19 $X=0.567 $Y=0.081
c74 38 VSS 0.00230547f $X=0.567 $Y=0.081
c75 33 VSS 0.00106687f $X=0.135 $Y=0.081
c76 21 VSS 0.00214349f $X=0.567 $Y=0.135
c77 18 VSS 0.0661718f $X=0.567 $Y=0.0675
c78 13 VSS 0.0184971f $X=0.297 $Y=0.135
c79 10 VSS 0.065697f $X=0.297 $Y=0.0675
c80 2 VSS 0.0639533f $X=0.135 $Y=0.0675
r81 62 63 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.118 $X2=0.567 $Y2=0.1265
r82 56 57 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.1305
r83 51 63 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.1265
r84 45 57 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.1305
r85 40 41 15.5494 $w=1.8e-08 $l=2.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.298
+ $Y=0.081 $X2=0.527 $Y2=0.081
r86 39 62 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.567 $Y2=0.118
r87 38 41 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.081 $X2=0.527 $Y2=0.081
r88 38 39 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.567 $Y=0.081 $X2=0.567
+ $Y2=0.081
r89 36 40 5.6358 $w=1.8e-08 $l=8.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.215
+ $Y=0.081 $X2=0.298 $Y2=0.081
r90 33 56 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.081 $X2=0.135 $Y2=0.126
r91 32 36 5.4321 $w=1.8e-08 $l=8e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.081 $X2=0.215 $Y2=0.081
r92 32 33 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.135 $Y=0.081 $X2=0.135
+ $Y2=0.081
r93 21 51 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r94 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r95 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r96 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r97 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r98 5 13 202.5 $w=1.6e-08 $l=1.62e-07 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.297 $Y2=0.135
r99 5 45 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r100 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r101 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_XOR2X1_ASAP7_75T_R%5 2 7 10 13 15 17 18 22 27 30 34 35 37 40 41 42 43
+ 46 48 49 50 51 54 56 57 60 VSS
c65 60 VSS 0.0012649f $X=0.1835 $Y=0.072
c66 57 VSS 2.07023e-20 $X=0.405 $Y=0.1305
c67 56 VSS 0.00144893f $X=0.405 $Y=0.126
c68 54 VSS 3.04905e-19 $X=0.405 $Y=0.135
c69 51 VSS 1.01588e-19 $X=0.365 $Y=0.072
c70 50 VSS 3.21516e-19 $X=0.305 $Y=0.072
c71 49 VSS 0.00264353f $X=0.256 $Y=0.072
c72 48 VSS 0.00102041f $X=0.213 $Y=0.072
c73 46 VSS 0.00225686f $X=0.396 $Y=0.072
c74 43 VSS 1.76975e-19 $X=0.183 $Y=0.149
c75 42 VSS 0.0015758f $X=0.183 $Y=0.126
c76 41 VSS 0.0131572f $X=0.183 $Y=0.174
c77 40 VSS 0.00153513f $X=0.183 $Y=0.174
c78 37 VSS 7.86306e-19 $X=0.1835 $Y=0.063
c79 35 VSS 0.0024907f $X=0.159 $Y=0.036
c80 34 VSS 0.00300662f $X=0.144 $Y=0.036
c81 30 VSS 0.0102544f $X=0.108 $Y=0.036
c82 29 VSS 0.00277426f $X=0.108 $Y=0.036
c83 27 VSS 0.00524826f $X=0.174 $Y=0.036
c84 25 VSS 4.79275e-19 $X=0.16 $Y=0.2025
c85 17 VSS 5.72255e-19 $X=0.125 $Y=0.0675
c86 13 VSS 0.00334187f $X=0.459 $Y=0.135
c87 10 VSS 0.0624922f $X=0.459 $Y=0.0675
c88 2 VSS 0.0619049f $X=0.405 $Y=0.0675
r89 56 57 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.126 $X2=0.405 $Y2=0.1305
r90 54 57 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.1305
r91 52 56 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.081 $X2=0.405 $Y2=0.126
r92 50 51 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.305
+ $Y=0.072 $X2=0.365 $Y2=0.072
r93 49 50 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.072 $X2=0.305 $Y2=0.072
r94 48 49 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.213
+ $Y=0.072 $X2=0.256 $Y2=0.072
r95 47 60 0.144403 $w=3.7e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.193
+ $Y=0.072 $X2=0.1835 $Y2=0.072
r96 47 48 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.193
+ $Y=0.072 $X2=0.213 $Y2=0.072
r97 46 52 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.072 $X2=0.405 $Y2=0.081
r98 46 51 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.072 $X2=0.365 $Y2=0.072
r99 42 43 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.183
+ $Y=0.126 $X2=0.183 $Y2=0.149
r100 40 43 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.183
+ $Y=0.174 $X2=0.183 $Y2=0.149
r101 40 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.183 $Y=0.174
+ $X2=0.183 $Y2=0.174
r102 38 60 0.505846 $w=1.9e-08 $l=9.24662e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.183 $Y=0.081 $X2=0.1835 $Y2=0.072
r103 38 42 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.183
+ $Y=0.081 $X2=0.183 $Y2=0.126
r104 37 60 0.505846 $w=1.9e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1835
+ $Y=0.063 $X2=0.1835 $Y2=0.072
r105 36 37 1.14327 $w=1.9e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1835
+ $Y=0.045 $X2=0.1835 $Y2=0.063
r106 34 35 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.159 $Y2=0.036
r107 29 34 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.144 $Y2=0.036
r108 29 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036
+ $X2=0.108 $Y2=0.036
r109 27 36 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.174 $Y=0.036 $X2=0.1835 $Y2=0.045
r110 27 35 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.174
+ $Y=0.036 $X2=0.159 $Y2=0.036
r111 25 41 11.8071 $w=5e-08 $l=2.85e-08 $layer=LISD $thickness=2.8e-08 $X=0.175
+ $Y=0.2025 $X2=0.175 $Y2=0.174
r112 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.16 $Y2=0.2025
r113 21 30 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.108 $Y=0.0675 $X2=0.108 $Y2=0.036
r114 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r115 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r116 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r117 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r118 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r119 5 54 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r120 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r121 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_XOR2X1_ASAP7_75T_R%Y 1 6 7 11 16 17 24 28 29 30 32 34 36 38 42 43 44
+ 46 51 53 54 VSS
c51 57 VSS 0.00176645f $X=0.459 $Y=0.036
c52 54 VSS 4.50279e-19 $X=0.45 $Y=0.184
c53 53 VSS 2.6023e-19 $X=0.459 $Y=0.184
c54 51 VSS 0.0032764f $X=0.432 $Y=0.184
c55 46 VSS 0.00439799f $X=0.576 $Y=0.036
c56 45 VSS 4.0861e-19 $X=0.526 $Y=0.036
c57 44 VSS 0.00147038f $X=0.522 $Y=0.036
c58 43 VSS 0.0062512f $X=0.504 $Y=0.036
c59 42 VSS 0.00359087f $X=0.594 $Y=0.036
c60 41 VSS 0.00513487f $X=0.594 $Y=0.036
c61 38 VSS 1.37072e-19 $X=0.459 $Y=0.149
c62 36 VSS 6.99723e-19 $X=0.459 $Y=0.081
c63 35 VSS 8.65169e-19 $X=0.459 $Y=0.063
c64 34 VSS 0.0010647f $X=0.457 $Y=0.092
c65 32 VSS 4.74957e-19 $X=0.459 $Y=0.175
c66 30 VSS 5.32692e-19 $X=0.418 $Y=0.036
c67 29 VSS 0.0161907f $X=0.414 $Y=0.036
c68 28 VSS 0.011938f $X=0.432 $Y=0.036
c69 24 VSS 0.00600583f $X=0.27 $Y=0.036
c70 21 VSS 0.00269031f $X=0.45 $Y=0.036
c71 16 VSS 5.83596e-19 $X=0.449 $Y=0.2025
c72 14 VSS 2.69461e-19 $X=0.592 $Y=0.0675
c73 6 VSS 5.25448e-19 $X=0.449 $Y=0.0675
c74 1 VSS 4.39464e-19 $X=0.287 $Y=0.0675
r75 54 55 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.184 $X2=0.4545 $Y2=0.184
r76 53 55 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.184 $X2=0.4545 $Y2=0.184
r77 50 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.184 $X2=0.45 $Y2=0.184
r78 50 51 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.184 $X2=0.432
+ $Y2=0.184
r79 45 46 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.526
+ $Y=0.036 $X2=0.576 $Y2=0.036
r80 44 45 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.036 $X2=0.526 $Y2=0.036
r81 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.036 $X2=0.522 $Y2=0.036
r82 41 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.036 $X2=0.576 $Y2=0.036
r83 41 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.036 $X2=0.594
+ $Y2=0.036
r84 39 57 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.459 $Y2=0.036
r85 39 43 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.504 $Y2=0.036
r86 37 38 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.118 $X2=0.459 $Y2=0.149
r87 35 36 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.063 $X2=0.459 $Y2=0.081
r88 34 37 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.092 $X2=0.459 $Y2=0.118
r89 34 36 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.092 $X2=0.459 $Y2=0.081
r90 32 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.175 $X2=0.459 $Y2=0.184
r91 32 38 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.175 $X2=0.459 $Y2=0.149
r92 31 57 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r93 31 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.063
r94 29 30 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.418 $Y2=0.036
r95 27 30 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.418 $Y2=0.036
r96 27 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r97 23 29 9.77778 $w=1.8e-08 $l=1.44e-07 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.414 $Y2=0.036
r98 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r99 21 57 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.459 $Y2=0.036
r100 21 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.432 $Y2=0.036
r101 20 51 15.9673 $w=2.4e-08 $l=1.85e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.2025 $X2=0.432 $Y2=0.184
r102 17 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r103 16 20 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r104 14 42 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.594 $Y=0.0675 $X2=0.594 $Y2=0.036
r105 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.0675 $X2=0.592 $Y2=0.0675
r106 10 28 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.432 $Y=0.0675 $X2=0.432 $Y2=0.036
r107 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r108 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
r109 4 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r110 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.272 $Y2=0.0675
.ends

.subckt PM_XOR2X1_ASAP7_75T_R%10 1 2 VSS
c2 1 VSS 0.00180539f $X=0.125 $Y=0.2025
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends


* END of "./XOR2x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt XOR2x1_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 N_5_M0_d N_A_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 VSS N_B_M1_g N_5_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_Y_M2_d N_B_M2_g noxref_8 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 noxref_8 N_A_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M4 N_Y_M4_d N_5_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M5 N_Y_M5_d N_5_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M6 noxref_9 N_A_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M7 N_Y_M7_d N_B_M7_g noxref_9 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M8 N_10_M8_d N_A_M8_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M9 N_5_M9_d N_B_M9_g N_10_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M10 VDD N_B_M10_g noxref_6 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 noxref_6 N_A_M11_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M12 N_Y_M12_d N_5_M12_g noxref_6 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M13 N_Y_M13_d N_5_M13_g noxref_6 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M14 noxref_6 N_A_M14_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M15 VDD N_B_M15_g noxref_6 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
*
* 
* .include "XOR2x1_ASAP7_75t_R.pex.sp.XOR2X1_ASAP7_75T_R.pxi"
* BEGIN of "./XOR2x1_ASAP7_75t_R.pex.sp.XOR2X1_ASAP7_75T_R.pxi"
* File: XOR2x1_ASAP7_75t_R.pex.sp.XOR2X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:07:55 2017
* 
x_PM_XOR2X1_ASAP7_75T_R%A N_A_M0_g N_A_c_6_p N_A_M8_g N_A_M3_g N_A_c_7_p
+ N_A_M11_g N_A_M6_g N_A_c_12_p N_A_M14_g A N_A_c_47_p N_A_c_64_p N_A_c_65_p
+ N_A_c_2_p N_A_c_8_p N_A_c_27_p N_A_c_31_p N_A_c_40_p N_A_c_4_p N_A_c_9_p
+ N_A_c_35_p N_A_c_55_p N_A_c_5_p N_A_c_10_p N_A_c_38_p N_A_c_18_p N_A_c_16_p
+ N_A_c_53_p N_A_c_20_p N_A_c_46_p VSS PM_XOR2X1_ASAP7_75T_R%A
x_PM_XOR2X1_ASAP7_75T_R%B N_B_M1_g N_B_M9_g N_B_M2_g N_B_c_71_n N_B_M10_g
+ N_B_M7_g N_B_c_77_n N_B_M15_g N_B_c_89_p B N_B_c_124_p N_B_c_122_p N_B_c_78_n
+ N_B_c_80_n N_B_c_82_n N_B_c_114_p N_B_c_83_n N_B_c_84_n N_B_c_121_p N_B_c_85_n
+ VSS PM_XOR2X1_ASAP7_75T_R%B
x_PM_XOR2X1_ASAP7_75T_R%5 N_5_M4_g N_5_M12_g N_5_M5_g N_5_c_135_n N_5_M13_g
+ N_5_M1_s N_5_M0_d N_5_M9_d N_5_c_186_p N_5_c_152_n N_5_c_154_n N_5_c_156_n
+ N_5_c_180_p N_5_c_137_n N_5_c_139_n N_5_c_159_n N_5_c_143_n N_5_c_163_n
+ N_5_c_164_n N_5_c_144_n N_5_c_145_n N_5_c_146_n N_5_c_175_p N_5_c_170_n
+ N_5_c_148_n N_5_c_171_n VSS PM_XOR2X1_ASAP7_75T_R%5
x_PM_XOR2X1_ASAP7_75T_R%Y N_Y_M2_d N_Y_M5_d N_Y_M4_d N_Y_M7_d N_Y_M13_d
+ N_Y_M12_d N_Y_c_205_n N_Y_c_207_n N_Y_c_196_n N_Y_c_209_n N_Y_c_197_n Y
+ N_Y_c_212_n N_Y_c_199_n N_Y_c_214_n N_Y_c_216_n N_Y_c_200_n N_Y_c_217_n
+ N_Y_c_236_n N_Y_c_202_n N_Y_c_204_n VSS PM_XOR2X1_ASAP7_75T_R%Y
x_PM_XOR2X1_ASAP7_75T_R%10 N_10_M9_s N_10_M8_d VSS PM_XOR2X1_ASAP7_75T_R%10
cc_1 N_A_M0_g N_B_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_M1_g 3.72893e-19 $X=0.144 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_3 N_A_M3_g N_B_M2_g 0.00323392f $X=0.351 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_4 N_A_c_4_p N_B_M2_g 3.987e-19 $X=0.305 $Y=0.194 $X2=0.297 $Y2=0.0675
cc_5 N_A_c_5_p N_B_M2_g 3.81992e-19 $X=0.314 $Y=0.175 $X2=0.297 $Y2=0.0675
cc_6 N_A_c_6_p N_B_c_71_n 8.12544e-19 $X=0.081 $Y=0.135 $X2=0.297 $Y2=0.135
cc_7 N_A_c_7_p N_B_c_71_n 0.00113906f $X=0.351 $Y=0.135 $X2=0.297 $Y2=0.135
cc_8 N_A_c_8_p N_B_c_71_n 2.65814e-19 $X=0.174 $Y=0.234 $X2=0.297 $Y2=0.135
cc_9 N_A_c_9_p N_B_c_71_n 0.0010895f $X=0.231 $Y=0.194 $X2=0.297 $Y2=0.135
cc_10 N_A_c_10_p N_B_c_71_n 0.00113991f $X=0.323 $Y=0.135 $X2=0.297 $Y2=0.135
cc_11 N_A_M6_g N_B_M7_g 0.00323392f $X=0.513 $Y=0.0675 $X2=0.567 $Y2=0.0675
cc_12 N_A_c_12_p N_B_c_77_n 9.33263e-19 $X=0.513 $Y=0.135 $X2=0.567 $Y2=0.135
cc_13 N_A_c_8_p N_B_c_78_n 2.55398e-19 $X=0.174 $Y=0.234 $X2=0.298 $Y2=0.081
cc_14 N_A_c_9_p N_B_c_78_n 9.35543e-19 $X=0.231 $Y=0.194 $X2=0.298 $Y2=0.081
cc_15 N_A_c_10_p N_B_c_80_n 3.08473e-19 $X=0.323 $Y=0.135 $X2=0.527 $Y2=0.081
cc_16 N_A_c_16_p N_B_c_80_n 0.00480718f $X=0.513 $Y=0.189 $X2=0.527 $Y2=0.081
cc_17 N_A_c_2_p N_B_c_82_n 3.94969e-19 $X=0.144 $Y=0.234 $X2=0.135 $Y2=0.135
cc_18 N_A_c_18_p N_B_c_83_n 4.8829e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.126
cc_19 A N_B_c_84_n 4.29558e-19 $X=0.06 $Y=0.134 $X2=0.135 $Y2=0.1305
cc_20 N_A_c_20_p N_B_c_85_n 0.00129773f $X=0.513 $Y=0.135 $X2=0.567 $Y2=0.1265
cc_21 N_A_M3_g N_5_M4_g 0.00323392f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_22 N_A_M6_g N_5_M4_g 2.69148e-19 $X=0.513 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_23 N_A_M3_g N_5_M5_g 2.69148e-19 $X=0.351 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_24 N_A_M6_g N_5_M5_g 0.00323392f $X=0.513 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_25 N_A_c_7_p N_5_c_135_n 0.00118234f $X=0.351 $Y=0.135 $X2=0.297 $Y2=0.135
cc_26 N_A_c_12_p N_5_c_135_n 9.33059e-19 $X=0.513 $Y=0.135 $X2=0.297 $Y2=0.135
cc_27 N_A_c_27_p N_5_c_137_n 6.81694e-19 $X=0.192 $Y=0.234 $X2=0.298 $Y2=0.081
cc_28 N_A_c_5_p N_5_c_137_n 2.53521e-19 $X=0.314 $Y=0.175 $X2=0.298 $Y2=0.081
cc_29 N_A_c_8_p N_5_c_139_n 0.00258171f $X=0.174 $Y=0.234 $X2=0.527 $Y2=0.081
cc_30 N_A_c_27_p N_5_c_139_n 0.00116706f $X=0.192 $Y=0.234 $X2=0.527 $Y2=0.081
cc_31 N_A_c_31_p N_5_c_139_n 8.50062e-19 $X=0.2025 $Y=0.234 $X2=0.527 $Y2=0.081
cc_32 N_A_c_9_p N_5_c_139_n 0.00100151f $X=0.231 $Y=0.194 $X2=0.527 $Y2=0.081
cc_33 N_A_c_10_p N_5_c_143_n 2.53521e-19 $X=0.323 $Y=0.135 $X2=0.135 $Y2=0.135
cc_34 N_A_c_9_p N_5_c_144_n 3.73122e-19 $X=0.231 $Y=0.194 $X2=0 $Y2=0
cc_35 N_A_c_35_p N_5_c_145_n 3.73122e-19 $X=0.2805 $Y=0.194 $X2=0.567 $Y2=0.135
cc_36 N_A_M3_g N_5_c_146_n 3.36975e-19 $X=0.351 $Y=0.0675 $X2=0.567 $Y2=0.135
cc_37 N_A_c_10_p N_5_c_146_n 0.00215596f $X=0.323 $Y=0.135 $X2=0.567 $Y2=0.135
cc_38 N_A_c_38_p N_5_c_148_n 8.71544e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.1305
cc_39 VSS N_A_c_35_p 2.87556e-19 $X=0.2805 $Y=0.194 $X2=0.135 $Y2=0.0675
cc_40 VSS N_A_c_40_p 9.1988e-19 $X=0.222 $Y=0.225 $X2=0.135 $Y2=0.135
cc_41 VSS N_A_c_4_p 4.50928e-19 $X=0.305 $Y=0.194 $X2=0.135 $Y2=0.135
cc_42 VSS N_A_c_35_p 0.00191341f $X=0.2805 $Y=0.194 $X2=0.135 $Y2=0.135
cc_43 VSS N_A_c_5_p 5.25032e-19 $X=0.314 $Y=0.175 $X2=0.135 $Y2=0.135
cc_44 VSS N_A_c_16_p 3.98572e-19 $X=0.513 $Y=0.189 $X2=0.297 $Y2=0.0675
cc_45 VSS N_A_c_16_p 2.66313e-19 $X=0.513 $Y=0.189 $X2=0.297 $Y2=0.2025
cc_46 VSS N_A_c_46_p 0.00100232f $X=0.513 $Y=0.169 $X2=0.297 $Y2=0.2025
cc_47 VSS N_A_c_47_p 0.00162699f $X=0.213 $Y=0.234 $X2=0 $Y2=0
cc_48 VSS N_A_c_35_p 0.00468689f $X=0.2805 $Y=0.194 $X2=0 $Y2=0
cc_49 VSS N_A_M3_g 4.26368e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_50 VSS N_A_c_38_p 4.87592e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_51 VSS N_A_c_16_p 0.00261669f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_52 VSS N_A_M6_g 2.63086e-19 $X=0.513 $Y=0.0675 $X2=0.527 $Y2=0.081
cc_53 VSS N_A_c_53_p 0.00133331f $X=0.513 $Y=0.189 $X2=0.527 $Y2=0.081
cc_54 N_A_M3_g N_Y_c_196_n 2.63664e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_55 N_A_c_55_p N_Y_c_197_n 2.51979e-19 $X=0.314 $Y=0.149 $X2=0.135 $Y2=0.081
cc_56 N_A_c_46_p N_Y_c_197_n 0.00102489f $X=0.513 $Y=0.169 $X2=0.135 $Y2=0.081
cc_57 N_A_c_20_p N_Y_c_199_n 0.00102489f $X=0.513 $Y=0.135 $X2=0.567 $Y2=0.081
cc_58 N_A_M6_g N_Y_c_200_n 3.7388e-19 $X=0.513 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_59 N_A_c_20_p N_Y_c_200_n 2.45728e-19 $X=0.513 $Y=0.135 $X2=0.135 $Y2=0.135
cc_60 N_A_c_16_p N_Y_c_202_n 6.12216e-19 $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_61 N_A_c_53_p N_Y_c_202_n 0.00102489f $X=0.513 $Y=0.189 $X2=0 $Y2=0
cc_62 N_A_c_16_p N_Y_c_204_n 6.55744e-19 $X=0.513 $Y=0.189 $X2=0.135 $Y2=0.081
cc_63 VSS N_A_c_10_p 5.39108e-19 $X=0.323 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_64 N_A_c_64_p N_10_M9_s 2.09605e-19 $X=0.107 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_65 N_A_c_65_p N_10_M9_s 2.34185e-19 $X=0.126 $Y=0.234 $X2=0.135 $Y2=0.0675
cc_66 N_B_M2_g N_5_M4_g 2.34385e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_67 N_B_M7_g N_5_M5_g 2.34385e-19 $X=0.567 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_68 N_B_c_80_n N_5_c_135_n 2.36611e-19 $X=0.527 $Y=0.081 $X2=0.351 $Y2=0.135
cc_69 N_B_c_89_p N_5_c_152_n 0.00122578f $X=0.135 $Y=0.081 $X2=0 $Y2=0
cc_70 N_B_c_83_n N_5_c_152_n 8.28374e-19 $X=0.135 $Y=0.126 $X2=0 $Y2=0
cc_71 N_B_M1_g N_5_c_154_n 2.34628e-19 $X=0.135 $Y=0.0675 $X2=0.018 $Y2=0.188
cc_72 N_B_c_89_p N_5_c_154_n 0.00367716f $X=0.135 $Y=0.081 $X2=0.018 $Y2=0.188
cc_73 N_B_c_71_n N_5_c_156_n 3.48111e-19 $X=0.297 $Y=0.135 $X2=0.027 $Y2=0.135
cc_74 N_B_c_78_n N_5_c_156_n 3.78066e-19 $X=0.298 $Y=0.081 $X2=0.027 $Y2=0.135
cc_75 N_B_c_71_n N_5_c_139_n 0.00247099f $X=0.297 $Y=0.135 $X2=0.213 $Y2=0.234
cc_76 N_B_c_78_n N_5_c_159_n 5.35839e-19 $X=0.298 $Y=0.081 $X2=0.027 $Y2=0.234
cc_77 N_B_c_83_n N_5_c_159_n 0.00160818f $X=0.135 $Y=0.126 $X2=0.027 $Y2=0.234
cc_78 N_B_c_71_n N_5_c_143_n 0.00210929f $X=0.297 $Y=0.135 $X2=0.078 $Y2=0.234
cc_79 N_B_c_82_n N_5_c_143_n 0.00148426f $X=0.135 $Y=0.135 $X2=0.078 $Y2=0.234
cc_80 N_B_c_80_n N_5_c_163_n 0.00133833f $X=0.527 $Y=0.081 $X2=0.126 $Y2=0.234
cc_81 N_B_c_71_n N_5_c_164_n 9.68215e-19 $X=0.297 $Y=0.135 $X2=0.174 $Y2=0.234
cc_82 N_B_c_78_n N_5_c_164_n 5.10242e-19 $X=0.298 $Y=0.081 $X2=0.174 $Y2=0.234
cc_83 N_B_c_78_n N_5_c_144_n 0.001214f $X=0.298 $Y=0.081 $X2=0.192 $Y2=0.234
cc_84 N_B_M2_g N_5_c_145_n 4.31042e-19 $X=0.297 $Y=0.0675 $X2=0.2025 $Y2=0.234
cc_85 N_B_c_78_n N_5_c_145_n 0.00109315f $X=0.298 $Y=0.081 $X2=0.2025 $Y2=0.234
cc_86 N_B_c_80_n N_5_c_146_n 0.00150184f $X=0.527 $Y=0.081 $X2=0.222 $Y2=0.203
cc_87 N_B_c_80_n N_5_c_170_n 7.13114e-19 $X=0.527 $Y=0.081 $X2=0.2805 $Y2=0.194
cc_88 N_B_c_89_p N_5_c_171_n 0.00148426f $X=0.135 $Y=0.081 $X2=0.314 $Y2=0.175
cc_89 N_B_c_78_n N_5_c_171_n 3.03428e-19 $X=0.298 $Y=0.081 $X2=0.314 $Y2=0.175
cc_90 VSS N_B_c_71_n 6.8292e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_91 VSS N_B_M2_g 2.82011e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_92 VSS N_B_c_80_n 3.45043e-19 $X=0.527 $Y=0.081 $X2=0.078 $Y2=0.234
cc_93 VSS N_B_M7_g 3.69259e-19 $X=0.567 $Y=0.0675 $X2=0.092 $Y2=0.234
cc_94 VSS N_B_c_114_p 3.92849e-19 $X=0.567 $Y=0.135 $X2=0.092 $Y2=0.234
cc_95 N_B_c_71_n N_Y_c_205_n 6.8292e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_96 N_B_c_78_n N_Y_c_205_n 4.64672e-19 $X=0.298 $Y=0.081 $X2=0 $Y2=0
cc_97 N_B_c_80_n N_Y_c_207_n 3.14976e-19 $X=0.527 $Y=0.081 $X2=0 $Y2=0
cc_98 N_B_M2_g N_Y_c_196_n 2.64369e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_99 N_B_c_80_n N_Y_c_209_n 4.77607e-19 $X=0.527 $Y=0.081 $X2=0 $Y2=0
cc_100 N_B_c_80_n Y 7.65288e-19 $X=0.527 $Y=0.081 $X2=0.018 $Y2=0.188
cc_101 N_B_c_121_p Y 5.08627e-19 $X=0.567 $Y=0.118 $X2=0.018 $Y2=0.188
cc_102 N_B_c_122_p N_Y_c_212_n 3.83522e-19 $X=0.567 $Y=0.081 $X2=0.06 $Y2=0.135
cc_103 N_B_c_80_n N_Y_c_212_n 4.49897e-19 $X=0.527 $Y=0.081 $X2=0.06 $Y2=0.135
cc_104 N_B_c_124_p N_Y_c_214_n 3.10247e-19 $X=0.567 $Y=0.081 $X2=0.027 $Y2=0.234
cc_105 N_B_c_122_p N_Y_c_214_n 0.00127078f $X=0.567 $Y=0.081 $X2=0.027 $Y2=0.234
cc_106 N_B_c_80_n N_Y_c_216_n 9.16084e-19 $X=0.527 $Y=0.081 $X2=0.078 $Y2=0.234
cc_107 N_B_M7_g N_Y_c_217_n 2.37298e-19 $X=0.567 $Y=0.0675 $X2=0.126 $Y2=0.234
cc_108 N_B_c_122_p N_Y_c_217_n 0.00506289f $X=0.567 $Y=0.081 $X2=0.126 $Y2=0.234
cc_109 N_B_c_80_n N_Y_c_204_n 2.40707e-19 $X=0.527 $Y=0.081 $X2=0.231 $Y2=0.194
cc_110 VSS N_B_c_122_p 3.03729e-19 $X=0.567 $Y=0.081 $X2=0.081 $Y2=0.0675
cc_111 VSS N_5_c_139_n 0.00251508f $X=0.183 $Y=0.174 $X2=0.081 $Y2=0.135
cc_112 VSS N_5_M4_g 3.77795e-19 $X=0.405 $Y=0.0675 $X2=0.018 $Y2=0.188
cc_113 VSS N_5_c_175_p 2.31252e-19 $X=0.405 $Y=0.135 $X2=0.018 $Y2=0.188
cc_114 VSS N_5_M5_g 2.86067e-19 $X=0.459 $Y=0.0675 $X2=0.06 $Y2=0.135
cc_115 N_5_c_145_n N_Y_M2_d 3.26345e-19 $X=0.305 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_116 N_5_c_135_n N_Y_M5_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_117 N_5_c_135_n N_Y_M13_d 4.0989e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_118 N_5_c_180_p N_Y_c_205_n 3.59575e-19 $X=0.1835 $Y=0.063 $X2=0 $Y2=0
cc_119 N_5_c_159_n N_Y_c_205_n 3.69284e-19 $X=0.183 $Y=0.126 $X2=0 $Y2=0
cc_120 N_5_c_145_n N_Y_c_205_n 0.00279801f $X=0.305 $Y=0.072 $X2=0 $Y2=0
cc_121 N_5_c_135_n N_Y_c_207_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_122 N_5_c_163_n N_Y_c_207_n 0.00107773f $X=0.396 $Y=0.072 $X2=0 $Y2=0
cc_123 N_5_M4_g N_Y_c_196_n 2.34002e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_124 N_5_c_186_p N_Y_c_196_n 6.66585e-19 $X=0.174 $Y=0.036 $X2=0 $Y2=0
cc_125 N_5_c_145_n N_Y_c_196_n 0.0130846f $X=0.305 $Y=0.072 $X2=0 $Y2=0
cc_126 N_5_M5_g Y 3.07672e-19 $X=0.459 $Y=0.0675 $X2=0.018 $Y2=0.188
cc_127 N_5_c_170_n Y 0.00120079f $X=0.405 $Y=0.126 $X2=0.018 $Y2=0.188
cc_128 N_5_c_163_n N_Y_c_212_n 0.00120079f $X=0.396 $Y=0.072 $X2=0.06 $Y2=0.135
cc_129 N_5_c_135_n N_Y_c_199_n 0.00230686f $X=0.459 $Y=0.135 $X2=0.064 $Y2=0.135
cc_130 N_5_c_175_p N_Y_c_199_n 0.00120079f $X=0.405 $Y=0.135 $X2=0.064 $Y2=0.135
cc_131 N_5_c_135_n N_Y_c_236_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.222 $Y2=0.203
cc_132 N_5_c_135_n N_Y_c_204_n 4.91185e-19 $X=0.459 $Y=0.135 $X2=0.231 $Y2=0.194
cc_133 VSS N_5_c_146_n 4.42394e-19 $X=0.365 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_134 VSS N_Y_c_205_n 0.00169333f $X=0.272 $Y=0.2025 $X2=0 $Y2=0
cc_135 VSS N_Y_c_197_n 6.21879e-19 $X=0.486 $Y=0.2025 $X2=0.018 $Y2=0.225
cc_136 VSS N_Y_c_214_n 0.00107252f $X=0.592 $Y=0.2025 $X2=0.027 $Y2=0.234
cc_137 VSS N_Y_c_236_n 0.0038608f $X=0.378 $Y=0.2025 $X2=0.222 $Y2=0.203
cc_138 VSS N_Y_c_236_n 0.00387022f $X=0.486 $Y=0.2025 $X2=0.222 $Y2=0.203
cc_139 VSS N_Y_c_236_n 0.00263673f $X=0.468 $Y=0.234 $X2=0.222 $Y2=0.203
cc_140 VSS N_Y_c_204_n 2.19246e-19 $X=0.378 $Y=0.2025 $X2=0.231 $Y2=0.194
cc_141 VSS N_Y_c_204_n 0.00238589f $X=0.468 $Y=0.234 $X2=0.231 $Y2=0.194
cc_142 VSS N_Y_c_196_n 3.19084e-19 $X=0.414 $Y=0.036 $X2=0.081 $Y2=0.0675

* END of "./XOR2x1_ASAP7_75t_R.pex.sp.XOR2X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: XOR2x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:08:17 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "XOR2x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./XOR2x2_ASAP7_75t_R.pex.sp.pex"
* File: XOR2x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:08:17 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_XOR2X2_ASAP7_75T_R%3 2 5 7 9 12 14 15 18 21 25 27 30 31 32 34 40 43
+ 45 46 VSS
c36 50 VSS 0.00179571f $X=0.311 $Y=0.198
c37 46 VSS 7.99121e-21 $X=0.36 $Y=0.198
c38 45 VSS 0.00213751f $X=0.342 $Y=0.198
c39 43 VSS 6.88106e-19 $X=0.378 $Y=0.198
c40 40 VSS 6.20662e-19 $X=0.311 $Y=0.163
c41 34 VSS 0.00174874f $X=0.311 $Y=0.09
c42 32 VSS 6.14081e-19 $X=0.311 $Y=0.189
c43 31 VSS 0.00208239f $X=0.279 $Y=0.198
c44 30 VSS 8.46035e-21 $X=0.144 $Y=0.198
c45 29 VSS 0.00220046f $X=0.126 $Y=0.198
c46 28 VSS 1.81812e-19 $X=0.099 $Y=0.198
c47 27 VSS 4.67334e-20 $X=0.09 $Y=0.198
c48 26 VSS 3.79585e-19 $X=0.302 $Y=0.198
c49 25 VSS 6.92425e-19 $X=0.081 $Y=0.1695
c50 21 VSS 4.12414e-19 $X=0.081 $Y=0.135
c51 19 VSS 9.17737e-19 $X=0.081 $Y=0.189
c52 18 VSS 0.024763f $X=0.378 $Y=0.216
c53 14 VSS 5.52978e-19 $X=0.395 $Y=0.216
c54 12 VSS 0.0143648f $X=0.326 $Y=0.0675
c55 9 VSS 4.79903e-19 $X=0.341 $Y=0.0675
c56 5 VSS 0.00172642f $X=0.081 $Y=0.135
c57 2 VSS 0.0664606f $X=0.081 $Y=0.0675
r58 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r59 43 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.198 $X2=0.36 $Y2=0.198
r60 41 50 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.32
+ $Y=0.198 $X2=0.311 $Y2=0.198
r61 41 45 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.32
+ $Y=0.198 $X2=0.342 $Y2=0.198
r62 39 40 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.15 $X2=0.311 $Y2=0.163
r63 34 39 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.09 $X2=0.311 $Y2=0.15
r64 32 50 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.189 $X2=0.311 $Y2=0.198
r65 32 40 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.189 $X2=0.311 $Y2=0.163
r66 30 31 9.16667 $w=1.8e-08 $l=1.35e-07 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.198 $X2=0.279 $Y2=0.198
r67 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.198 $X2=0.144 $Y2=0.198
r68 28 29 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.198 $X2=0.126 $Y2=0.198
r69 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.198 $X2=0.099 $Y2=0.198
r70 26 50 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.302
+ $Y=0.198 $X2=0.311 $Y2=0.198
r71 26 31 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.302
+ $Y=0.198 $X2=0.279 $Y2=0.198
r72 24 25 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.15 $X2=0.081 $Y2=0.1695
r73 21 24 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.15
r74 19 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.189 $X2=0.09 $Y2=0.198
r75 19 25 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.189 $X2=0.081 $Y2=0.1695
r76 18 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.198 $X2=0.378
+ $Y2=0.198
r77 15 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.216 $X2=0.378 $Y2=0.216
r78 14 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.216 $X2=0.378 $Y2=0.216
r79 12 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.311 $Y=0.09 $X2=0.311
+ $Y2=0.09
r80 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.0675 $X2=0.326 $Y2=0.0675
r81 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r82 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r83 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_XOR2X2_ASAP7_75T_R%B 2 5 7 10 13 15 19 22 24 25 26 30 31 32 33 34 35
+ 36 37 43 44 45 50 VSS
c45 50 VSS 0.00219816f $X=0.429 $Y=0.135
c46 45 VSS 4.62983e-20 $X=0.431 $Y=0.1225
c47 44 VSS 0.00266656f $X=0.431 $Y=0.119
c48 43 VSS 0.00109749f $X=0.431 $Y=0.081
c49 42 VSS 9.62667e-19 $X=0.431 $Y=0.063
c50 41 VSS 1.23361e-19 $X=0.431 $Y=0.126
c51 39 VSS 0.00128265f $X=0.4065 $Y=0.036
c52 38 VSS 0.00120569f $X=0.391 $Y=0.036
c53 37 VSS 0.00322944f $X=0.38 $Y=0.036
c54 36 VSS 0.00199133f $X=0.342 $Y=0.036
c55 35 VSS 0.00134741f $X=0.32 $Y=0.036
c56 34 VSS 0.00205247f $X=0.302 $Y=0.036
c57 33 VSS 0.00231441f $X=0.279 $Y=0.036
c58 32 VSS 0.00518759f $X=0.422 $Y=0.036
c59 31 VSS 5.2764e-21 $X=0.27 $Y=0.066
c60 30 VSS 6.78204e-20 $X=0.27 $Y=0.063
c61 29 VSS 4.397e-21 $X=0.27 $Y=0.069
c62 27 VSS 8.52667e-19 $X=0.2455 $Y=0.078
c63 26 VSS 0.00320415f $X=0.23 $Y=0.078
c64 25 VSS 5.19699e-20 $X=0.144 $Y=0.078
c65 24 VSS 9.86545e-19 $X=0.261 $Y=0.078
c66 22 VSS 3.81104e-19 $X=0.135 $Y=0.128
c67 21 VSS 0.00125483f $X=0.135 $Y=0.121
c68 19 VSS 5.20634e-20 $X=0.135 $Y=0.135
c69 13 VSS 0.00157266f $X=0.405 $Y=0.135
c70 10 VSS 0.0593607f $X=0.405 $Y=0.0675
c71 5 VSS 0.00145372f $X=0.135 $Y=0.135
c72 2 VSS 0.0618866f $X=0.135 $Y=0.0675
r73 50 51 0.0987654 $w=2.475e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.429
+ $Y=0.144 $X2=0.431 $Y2=0.144
r74 47 50 1.18519 $w=2.475e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.144 $X2=0.429 $Y2=0.144
r75 44 45 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.119 $X2=0.431 $Y2=0.1225
r76 43 44 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.081 $X2=0.431 $Y2=0.119
r77 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.063 $X2=0.431 $Y2=0.081
r78 41 51 0.260825 $w=2.475e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.126 $X2=0.431 $Y2=0.144
r79 41 45 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.126 $X2=0.431 $Y2=0.1225
r80 40 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.045 $X2=0.431 $Y2=0.063
r81 38 39 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.391
+ $Y=0.036 $X2=0.4065 $Y2=0.036
r82 37 38 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.38
+ $Y=0.036 $X2=0.391 $Y2=0.036
r83 36 37 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.38 $Y2=0.036
r84 35 36 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.32
+ $Y=0.036 $X2=0.342 $Y2=0.036
r85 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.302
+ $Y=0.036 $X2=0.32 $Y2=0.036
r86 33 34 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.036 $X2=0.302 $Y2=0.036
r87 32 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.422 $Y=0.036 $X2=0.431 $Y2=0.045
r88 32 39 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.422
+ $Y=0.036 $X2=0.4065 $Y2=0.036
r89 30 31 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.063 $X2=0.27 $Y2=0.066
r90 29 31 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.069 $X2=0.27 $Y2=0.066
r91 28 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.27 $Y=0.045 $X2=0.279 $Y2=0.036
r92 28 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.045 $X2=0.27 $Y2=0.063
r93 26 27 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.078 $X2=0.2455 $Y2=0.078
r94 25 26 5.83951 $w=1.8e-08 $l=8.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.078 $X2=0.23 $Y2=0.078
r95 24 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.261 $Y=0.078 $X2=0.27 $Y2=0.069
r96 24 27 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.078 $X2=0.2455 $Y2=0.078
r97 21 22 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.121 $X2=0.135 $Y2=0.128
r98 19 22 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.128
r99 17 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.087 $X2=0.144 $Y2=0.078
r100 17 21 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.087 $X2=0.135 $Y2=0.121
r101 13 47 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r102 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.216
r103 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r104 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r105 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r106 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_XOR2X2_ASAP7_75T_R%A 2 7 10 13 15 19 21 24 VSS
c33 24 VSS 1.44512e-20 $X=0.351 $Y=0.1305
c34 21 VSS 2.12541e-19 $X=0.351 $Y=0.135
c35 19 VSS 0.00136948f $X=0.351 $Y=0.102
c36 13 VSS 0.0161676f $X=0.351 $Y=0.135
c37 10 VSS 0.0634112f $X=0.351 $Y=0.0675
c38 2 VSS 0.0655165f $X=0.189 $Y=0.0675
r39 23 24 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.126 $X2=0.351 $Y2=0.1305
r40 21 24 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.1305
r41 19 23 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.102 $X2=0.351 $Y2=0.126
r42 13 21 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r43 13 15 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.216
r44 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r45 5 13 202.5 $w=1.6e-08 $l=1.62e-07 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.351 $Y2=0.135
r46 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r47 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_XOR2X2_ASAP7_75T_R%6 2 7 10 13 15 17 22 25 27 30 35 36 38 48 49 52 53
+ 55 56 58 62 66 67 VSS
c45 69 VSS 9.17717e-19 $X=0.045 $Y=0.036
c46 68 VSS 0.00328948f $X=0.036 $Y=0.036
c47 67 VSS 0.002959f $X=0.054 $Y=0.036
c48 66 VSS 0.0023031f $X=0.054 $Y=0.036
c49 62 VSS 2.80912e-19 $X=0.486 $Y=0.176
c50 58 VSS 9.45598e-19 $X=0.486 $Y=0.135
c51 56 VSS 2.70108e-19 $X=0.486 $Y=0.189
c52 55 VSS 5.06567e-20 $X=0.4745 $Y=0.198
c53 54 VSS 0.00185179f $X=0.472 $Y=0.198
c54 53 VSS 0.00117446f $X=0.441 $Y=0.198
c55 52 VSS 1.3551e-19 $X=0.477 $Y=0.198
c56 51 VSS 6.41935e-19 $X=0.432 $Y=0.225
c57 49 VSS 0.00308828f $X=0.422 $Y=0.234
c58 48 VSS 0.0323459f $X=0.392 $Y=0.234
c59 47 VSS 8.76814e-19 $X=0.072 $Y=0.234
c60 46 VSS 0.00270525f $X=0.063 $Y=0.234
c61 39 VSS 0.00341041f $X=0.036 $Y=0.234
c62 38 VSS 0.00309411f $X=0.423 $Y=0.234
c63 37 VSS 2.98008e-19 $X=0.027 $Y=0.216
c64 36 VSS 0.00366991f $X=0.027 $Y=0.207
c65 35 VSS 0.00237432f $X=0.027 $Y=0.121
c66 34 VSS 7.78132e-19 $X=0.027 $Y=0.069
c67 33 VSS 2.81452e-19 $X=0.027 $Y=0.225
c68 30 VSS 0.00549743f $X=0.214 $Y=0.2025
c69 25 VSS 0.00677526f $X=0.056 $Y=0.2025
c70 22 VSS 2.69461e-19 $X=0.071 $Y=0.2025
c71 17 VSS 3.25039e-19 $X=0.071 $Y=0.0675
c72 13 VSS 0.00427912f $X=0.513 $Y=0.135
c73 10 VSS 0.0639847f $X=0.513 $Y=0.0675
c74 2 VSS 0.0613093f $X=0.459 $Y=0.0675
r75 68 69 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.045 $Y2=0.036
r76 66 69 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.045 $Y2=0.036
r77 66 67 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r78 63 68 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.036 $Y2=0.036
r79 61 62 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.163 $X2=0.486 $Y2=0.176
r80 58 61 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.135 $X2=0.486 $Y2=0.163
r81 58 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.486 $Y=0.135 $X2=0.486
+ $Y2=0.135
r82 56 62 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.189 $X2=0.486 $Y2=0.176
r83 54 55 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.472
+ $Y=0.198 $X2=0.4745 $Y2=0.198
r84 53 54 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.441
+ $Y=0.198 $X2=0.472 $Y2=0.198
r85 52 56 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.477 $Y=0.198 $X2=0.486 $Y2=0.189
r86 52 55 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.477
+ $Y=0.198 $X2=0.4745 $Y2=0.198
r87 50 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.432 $Y=0.207 $X2=0.441 $Y2=0.198
r88 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.207 $X2=0.432 $Y2=0.225
r89 48 49 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.392
+ $Y=0.234 $X2=0.422 $Y2=0.234
r90 46 47 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.234 $X2=0.072 $Y2=0.234
r91 44 48 11.9506 $w=1.8e-08 $l=1.76e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.392 $Y2=0.234
r92 44 47 9.77778 $w=1.8e-08 $l=1.44e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.234 $X2=0.072 $Y2=0.234
r93 41 46 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.063 $Y2=0.234
r94 39 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.054 $Y2=0.234
r95 38 51 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.423 $Y=0.234 $X2=0.432 $Y2=0.225
r96 38 49 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.423
+ $Y=0.234 $X2=0.422 $Y2=0.234
r97 36 37 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.207 $X2=0.027 $Y2=0.216
r98 35 36 5.83951 $w=1.8e-08 $l=8.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.121 $X2=0.027 $Y2=0.207
r99 34 35 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.069 $X2=0.027 $Y2=0.121
r100 33 39 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.225 $X2=0.036 $Y2=0.234
r101 33 37 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.216
r102 32 63 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.036
r103 32 34 1.62963 $w=1.8e-08 $l=2.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.069
r104 30 44 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.234
+ $X2=0.216 $Y2=0.234
r105 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.214 $Y2=0.2025
r106 25 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r107 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r108 20 67 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.054 $Y=0.0675 $X2=0.054 $Y2=0.036
r109 17 20 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r110 13 59 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.486 $Y2=0.135
r111 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r112 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r113 5 59 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.486 $Y2=0.135
r114 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r115 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_XOR2X2_ASAP7_75T_R%Y 1 2 6 7 10 13 14 19 25 26 30 31 32 VSS
c21 34 VSS 4.55454e-19 $X=0.567 $Y=0.216
c22 32 VSS 6.60149e-19 $X=0.567 $Y=0.13325
c23 31 VSS 0.00413443f $X=0.567 $Y=0.119
c24 30 VSS 0.00358963f $X=0.567 $Y=0.1475
c25 28 VSS 4.30151e-19 $X=0.567 $Y=0.225
c26 26 VSS 0.00278214f $X=0.5265 $Y=0.234
c27 25 VSS 0.00252246f $X=0.495 $Y=0.234
c28 20 VSS 0.00875248f $X=0.558 $Y=0.234
c29 19 VSS 0.00278214f $X=0.5265 $Y=0.036
c30 18 VSS 0.00107061f $X=0.495 $Y=0.036
c31 14 VSS 0.00915654f $X=0.486 $Y=0.036
c32 13 VSS 0.00154248f $X=0.486 $Y=0.036
c33 11 VSS 0.00875248f $X=0.558 $Y=0.036
c34 10 VSS 0.0108098f $X=0.486 $Y=0.2025
c35 6 VSS 6.04166e-19 $X=0.503 $Y=0.2025
c36 1 VSS 5.72268e-19 $X=0.503 $Y=0.0675
r37 33 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.207 $X2=0.567 $Y2=0.216
r38 31 32 0.967593 $w=1.8e-08 $l=1.425e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.119 $X2=0.567 $Y2=0.13325
r39 30 33 4.04012 $w=1.8e-08 $l=5.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.1475 $X2=0.567 $Y2=0.207
r40 30 32 0.967593 $w=1.8e-08 $l=1.425e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.1475 $X2=0.567 $Y2=0.13325
r41 28 34 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.225 $X2=0.567 $Y2=0.216
r42 27 31 5.02469 $w=1.8e-08 $l=7.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.045 $X2=0.567 $Y2=0.119
r43 25 26 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.234 $X2=0.5265 $Y2=0.234
r44 22 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.495 $Y2=0.234
r45 20 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.234 $X2=0.567 $Y2=0.225
r46 20 26 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.5265 $Y2=0.234
r47 18 19 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.036 $X2=0.5265 $Y2=0.036
r48 13 18 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.495 $Y2=0.036
r49 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036 $X2=0.486
+ $Y2=0.036
r50 11 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.036 $X2=0.567 $Y2=0.045
r51 11 19 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.5265 $Y2=0.036
r52 10 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r53 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.486 $Y2=0.2025
r54 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.2025 $X2=0.486 $Y2=0.2025
r55 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0675 $X2=0.486 $Y2=0.036
r56 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.0675 $X2=0.486 $Y2=0.0675
r57 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0675 $X2=0.486 $Y2=0.0675
.ends

.subckt PM_XOR2X2_ASAP7_75T_R%9 1 2 VSS
c0 1 VSS 0.00243711f $X=0.395 $Y=0.0675
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.361 $Y2=0.0675
.ends


* END of "./XOR2x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt XOR2x2_ASAP7_75t_R  VSS VDD B A Y
* 
* Y	Y
* A	A
* B	B
M0 noxref_7 N_3_M0_g N_6_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 VSS N_B_M1_g noxref_7 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 noxref_7 N_A_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_9_M3_d N_A_M3_g N_3_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M4 VSS N_B_M4_g N_9_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M5 N_Y_M5_d N_6_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M6 N_Y_M6_d N_6_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M7 VDD N_3_M7_g N_6_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M8 noxref_10 N_B_M8_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M9 N_6_M9_d N_A_M9_g noxref_10 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M10 N_3_M10_d N_A_M10_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341
+ $Y=0.189
M11 VDD N_B_M11_g N_3_M11_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.395
+ $Y=0.189
M12 N_Y_M12_d N_6_M12_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M13 N_Y_M13_d N_6_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
*
* 
* .include "XOR2x2_ASAP7_75t_R.pex.sp.XOR2X2_ASAP7_75T_R.pxi"
* BEGIN of "./XOR2x2_ASAP7_75t_R.pex.sp.XOR2X2_ASAP7_75T_R.pxi"
* File: XOR2x2_ASAP7_75t_R.pex.sp.XOR2X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:08:17 2017
* 
x_PM_XOR2X2_ASAP7_75T_R%3 N_3_M0_g N_3_c_3_p N_3_M7_g N_3_M3_s N_3_c_8_p
+ N_3_M11_s N_3_M10_d N_3_c_31_p N_3_c_5_p N_3_c_26_p N_3_c_32_p N_3_c_2_p
+ N_3_c_7_p N_3_c_34_p N_3_c_6_p N_3_c_23_p N_3_c_22_p N_3_c_19_p N_3_c_15_p VSS
+ PM_XOR2X2_ASAP7_75T_R%3
x_PM_XOR2X2_ASAP7_75T_R%B N_B_M1_g N_B_c_39_n N_B_M8_g N_B_M4_g N_B_c_54_p
+ N_B_M11_g N_B_c_40_n N_B_c_41_n N_B_c_42_n N_B_c_66_p N_B_c_43_n N_B_c_44_n
+ N_B_c_57_p N_B_c_80_p N_B_c_75_p N_B_c_45_n N_B_c_46_n N_B_c_48_n N_B_c_52_p
+ N_B_c_59_p N_B_c_60_p N_B_c_71_p B VSS PM_XOR2X2_ASAP7_75T_R%B
x_PM_XOR2X2_ASAP7_75T_R%A N_A_M2_g N_A_M9_g N_A_M3_g N_A_c_85_n N_A_M10_g A
+ N_A_c_92_n N_A_c_94_n VSS PM_XOR2X2_ASAP7_75T_R%A
x_PM_XOR2X2_ASAP7_75T_R%6 N_6_M5_g N_6_M12_g N_6_M6_g N_6_c_126_n N_6_M13_g
+ N_6_M0_s N_6_M7_s N_6_c_115_n N_6_M9_d N_6_c_116_n N_6_c_127_n N_6_c_118_n
+ N_6_c_152_p N_6_c_119_n N_6_c_129_n N_6_c_143_p N_6_c_122_n N_6_c_144_p
+ N_6_c_145_p N_6_c_132_n N_6_c_123_n N_6_c_139_p N_6_c_137_p VSS
+ PM_XOR2X2_ASAP7_75T_R%6
x_PM_XOR2X2_ASAP7_75T_R%Y N_Y_M6_d N_Y_M5_d N_Y_M13_d N_Y_M12_d N_Y_c_164_n
+ N_Y_c_160_n N_Y_c_171_n N_Y_c_172_n N_Y_c_174_n N_Y_c_176_n Y N_Y_c_161_n
+ N_Y_c_179_n VSS PM_XOR2X2_ASAP7_75T_R%Y
x_PM_XOR2X2_ASAP7_75T_R%9 N_9_M4_s N_9_M3_d VSS PM_XOR2X2_ASAP7_75T_R%9
cc_1 N_3_M0_g N_B_M1_g 0.00323392f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_3_c_2_p N_B_M1_g 2.98356e-19 $X=0.144 $Y=0.198 $X2=0.135 $Y2=0.0675
cc_3 N_3_c_3_p N_B_c_39_n 9.46013e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_3_c_2_p N_B_c_40_n 7.96353e-19 $X=0.144 $Y=0.198 $X2=0.135 $Y2=0.135
cc_5 N_3_c_5_p N_B_c_41_n 0.00118958f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.128
cc_6 N_3_c_6_p N_B_c_42_n 7.27089e-19 $X=0.311 $Y=0.09 $X2=0.261 $Y2=0.078
cc_7 N_3_c_7_p N_B_c_43_n 0.00164688f $X=0.279 $Y=0.198 $X2=0.23 $Y2=0.078
cc_8 N_3_c_8_p N_B_c_44_n 4.55331e-19 $X=0.326 $Y=0.0675 $X2=0.27 $Y2=0.063
cc_9 N_3_c_8_p N_B_c_45_n 0.00117999f $X=0.326 $Y=0.0675 $X2=0.302 $Y2=0.036
cc_10 N_3_c_8_p N_B_c_46_n 0.0012608f $X=0.326 $Y=0.0675 $X2=0.32 $Y2=0.036
cc_11 N_3_c_6_p N_B_c_46_n 8.67348e-19 $X=0.311 $Y=0.09 $X2=0.32 $Y2=0.036
cc_12 N_3_c_8_p N_B_c_48_n 0.00195414f $X=0.326 $Y=0.0675 $X2=0.342 $Y2=0.036
cc_13 N_3_M0_g N_A_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_14 N_3_c_7_p N_A_M2_g 4.07897e-19 $X=0.279 $Y=0.198 $X2=0.135 $Y2=0.0675
cc_15 N_3_c_15_p N_A_M3_g 2.81878e-19 $X=0.36 $Y=0.198 $X2=0.405 $Y2=0.0675
cc_16 N_3_c_8_p N_A_c_85_n 0.00268514f $X=0.326 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_17 N_3_c_7_p N_A_c_85_n 0.00128776f $X=0.279 $Y=0.198 $X2=0.405 $Y2=0.135
cc_18 N_3_c_6_p N_A_c_85_n 0.00237361f $X=0.311 $Y=0.09 $X2=0.405 $Y2=0.135
cc_19 N_3_c_19_p N_A_c_85_n 5.46915e-19 $X=0.342 $Y=0.198 $X2=0.405 $Y2=0.135
cc_20 N_3_c_8_p A 0.00117729f $X=0.326 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_21 N_3_c_6_p A 0.0030137f $X=0.311 $Y=0.09 $X2=0.135 $Y2=0.135
cc_22 N_3_c_22_p A 2.72962e-19 $X=0.378 $Y=0.198 $X2=0.135 $Y2=0.135
cc_23 N_3_c_23_p N_A_c_92_n 0.00150685f $X=0.311 $Y=0.163 $X2=0.135 $Y2=0.121
cc_24 N_3_c_15_p N_A_c_92_n 0.00119465f $X=0.36 $Y=0.198 $X2=0.135 $Y2=0.121
cc_25 N_3_c_6_p N_A_c_94_n 0.00150685f $X=0.311 $Y=0.09 $X2=0.261 $Y2=0.078
cc_26 N_3_c_26_p N_6_c_115_n 0.00136014f $X=0.081 $Y=0.1695 $X2=0.144 $Y2=0.078
cc_27 N_3_c_7_p N_6_c_116_n 0.0031568f $X=0.279 $Y=0.198 $X2=0.27 $Y2=0.063
cc_28 N_3_c_23_p N_6_c_116_n 6.58653e-19 $X=0.311 $Y=0.163 $X2=0.27 $Y2=0.063
cc_29 N_3_c_5_p N_6_c_118_n 0.00344236f $X=0.081 $Y=0.135 $X2=0.342 $Y2=0.036
cc_30 N_3_M0_g N_6_c_119_n 2.34993e-19 $X=0.081 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_31 N_3_c_31_p N_6_c_119_n 0.00255062f $X=0.378 $Y=0.216 $X2=0.405 $Y2=0.135
cc_32 N_3_c_32_p N_6_c_119_n 0.0270759f $X=0.09 $Y=0.198 $X2=0.405 $Y2=0.135
cc_33 N_3_c_22_p N_6_c_122_n 9.4025e-19 $X=0.378 $Y=0.198 $X2=0 $Y2=0
cc_34 N_3_c_34_p N_6_c_123_n 2.07298e-19 $X=0.311 $Y=0.189 $X2=0 $Y2=0
cc_35 VSS N_3_c_8_p 0.00216384f $X=0.326 $Y=0.0675 $X2=0.135 $Y2=0.087
cc_36 VSS N_3_c_7_p 5.0983e-19 $X=0.279 $Y=0.198 $X2=0.135 $Y2=0.0675
cc_37 N_B_M1_g N_A_M2_g 0.00323392f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_38 N_B_c_43_n N_A_M2_g 4.15003e-19 $X=0.23 $Y=0.078 $X2=0.081 $Y2=0.0675
cc_39 N_B_M4_g N_A_M3_g 0.00344695f $X=0.405 $Y=0.0675 $X2=0.326 $Y2=0.0675
cc_40 N_B_c_52_p N_A_M3_g 2.38942e-19 $X=0.38 $Y=0.036 $X2=0.326 $Y2=0.0675
cc_41 N_B_c_39_n N_A_c_85_n 0.00106649f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_42 N_B_c_54_p N_A_c_85_n 8.77417e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_43 N_B_c_43_n N_A_c_85_n 0.00133346f $X=0.23 $Y=0.078 $X2=0 $Y2=0
cc_44 N_B_c_48_n N_A_c_85_n 2.02767e-19 $X=0.342 $Y=0.036 $X2=0 $Y2=0
cc_45 N_B_c_57_p A 3.38087e-19 $X=0.27 $Y=0.066 $X2=0.081 $Y2=0.189
cc_46 N_B_c_52_p A 0.00408388f $X=0.38 $Y=0.036 $X2=0.081 $Y2=0.189
cc_47 N_B_c_59_p A 6.32476e-19 $X=0.431 $Y=0.081 $X2=0.081 $Y2=0.189
cc_48 N_B_c_60_p A 0.00111817f $X=0.431 $Y=0.119 $X2=0.081 $Y2=0.189
cc_49 B N_A_c_92_n 5.60486e-19 $X=0.429 $Y=0.135 $X2=0.081 $Y2=0.135
cc_50 B N_A_c_94_n 8.81039e-19 $X=0.429 $Y=0.135 $X2=0.081 $Y2=0.15
cc_51 N_B_M4_g N_6_M5_g 0.00284417f $X=0.405 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_52 N_B_M4_g N_6_M6_g 2.31381e-19 $X=0.405 $Y=0.0675 $X2=0.326 $Y2=0.0675
cc_53 N_B_c_54_p N_6_c_126_n 9.54501e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_54 N_B_c_66_p N_6_c_127_n 5.62087e-19 $X=0.144 $Y=0.078 $X2=0.311 $Y2=0.09
cc_55 N_B_M1_g N_6_c_119_n 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_56 N_B_M4_g N_6_c_129_n 4.28653e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_57 B N_6_c_129_n 5.57996e-19 $X=0.429 $Y=0.135 $X2=0 $Y2=0
cc_58 B N_6_c_122_n 0.00101601f $X=0.429 $Y=0.135 $X2=0 $Y2=0
cc_59 N_B_c_71_p N_6_c_132_n 0.00200427f $X=0.431 $Y=0.1225 $X2=0 $Y2=0
cc_60 VSS N_B_c_43_n 3.32448e-19 $X=0.23 $Y=0.078 $X2=0.341 $Y2=0.0675
cc_61 VSS N_B_c_66_p 0.00137624f $X=0.144 $Y=0.078 $X2=0 $Y2=0
cc_62 VSS N_B_c_43_n 0.00337967f $X=0.23 $Y=0.078 $X2=0.378 $Y2=0.216
cc_63 VSS N_B_c_75_p 0.00123078f $X=0.279 $Y=0.036 $X2=0.378 $Y2=0.216
cc_64 VSS N_B_c_43_n 0.00222818f $X=0.23 $Y=0.078 $X2=0 $Y2=0
cc_65 VSS N_B_c_44_n 8.24756e-19 $X=0.27 $Y=0.063 $X2=0 $Y2=0
cc_66 VSS N_B_M1_g 2.60742e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.189
cc_67 VSS N_B_c_66_p 0.00337967f $X=0.144 $Y=0.078 $X2=0.081 $Y2=0.189
cc_68 N_B_c_80_p N_Y_c_160_n 0.00108419f $X=0.422 $Y=0.036 $X2=0 $Y2=0
cc_69 N_B_c_59_p N_Y_c_161_n 4.77035e-19 $X=0.431 $Y=0.081 $X2=0.279 $Y2=0.198
cc_70 N_A_M3_g N_6_M5_g 2.31381e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_71 N_A_c_85_n N_6_c_116_n 6.8292e-19 $X=0.351 $Y=0.135 $X2=0.144 $Y2=0.198
cc_72 N_A_M2_g N_6_c_119_n 2.65491e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_73 N_A_M3_g N_6_c_119_n 2.38942e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_74 VSS N_A_M2_g 2.90722e-19 $X=0.189 $Y=0.0675 $X2=0.378 $Y2=0.216
cc_75 VSS N_A_c_85_n 6.8292e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_76 VSS N_6_c_137_p 0.00391186f $X=0.054 $Y=0.036 $X2=0 $Y2=0
cc_77 VSS N_6_c_116_n 0.00169333f $X=0.214 $Y=0.2025 $X2=0 $Y2=0
cc_78 VSS N_6_c_139_p 6.5272e-19 $X=0.054 $Y=0.036 $X2=0.378 $Y2=0.216
cc_79 N_6_c_126_n N_Y_M6_d 3.80663e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_80 N_6_c_126_n N_Y_M13_d 3.80455e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_81 N_6_c_126_n N_Y_c_164_n 8.00061e-19 $X=0.513 $Y=0.135 $X2=0.326 $Y2=0.0675
cc_82 N_6_c_143_p N_Y_c_164_n 0.00130196f $X=0.477 $Y=0.198 $X2=0.326 $Y2=0.0675
cc_83 N_6_c_144_p N_Y_c_164_n 3.88373e-19 $X=0.4745 $Y=0.198 $X2=0.326
+ $Y2=0.0675
cc_84 N_6_c_145_p N_Y_c_164_n 7.24049e-19 $X=0.486 $Y=0.189 $X2=0.326 $Y2=0.0675
cc_85 N_6_c_132_n N_Y_c_164_n 5.3153e-19 $X=0.486 $Y=0.135 $X2=0.326 $Y2=0.0675
cc_86 N_6_c_123_n N_Y_c_164_n 7.53011e-19 $X=0.486 $Y=0.176 $X2=0.326 $Y2=0.0675
cc_87 N_6_c_132_n N_Y_c_160_n 3.89018e-19 $X=0.486 $Y=0.135 $X2=0 $Y2=0
cc_88 N_6_c_126_n N_Y_c_171_n 5.9618e-19 $X=0.513 $Y=0.135 $X2=0.395 $Y2=0.216
cc_89 N_6_M6_g N_Y_c_172_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.081 $Y2=0.189
cc_90 N_6_c_126_n N_Y_c_172_n 3.25494e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.189
cc_91 N_6_c_152_p N_Y_c_174_n 9.63474e-19 $X=0.423 $Y=0.234 $X2=0.081 $Y2=0.1695
cc_92 N_6_c_144_p N_Y_c_174_n 0.00176732f $X=0.4745 $Y=0.198 $X2=0.081
+ $Y2=0.1695
cc_93 N_6_M6_g N_Y_c_176_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.302 $Y2=0.198
cc_94 N_6_c_126_n N_Y_c_176_n 3.25494e-19 $X=0.513 $Y=0.135 $X2=0.302 $Y2=0.198
cc_95 N_6_c_145_p Y 9.12629e-19 $X=0.486 $Y=0.189 $X2=0.144 $Y2=0.198
cc_96 N_6_c_126_n N_Y_c_179_n 3.78282e-19 $X=0.513 $Y=0.135 $X2=0.311 $Y2=0.189
cc_97 N_6_c_132_n N_Y_c_179_n 9.12629e-19 $X=0.486 $Y=0.135 $X2=0.311 $Y2=0.189
cc_98 VSS N_6_c_119_n 3.33359e-19 $X=0.392 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./XOR2x2_ASAP7_75t_R.pex.sp.XOR2X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: XOR2xp5_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:08:40 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "XOR2xp5_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./XOR2xp5_ASAP7_75t_R.pex.sp.pex"
* File: XOR2xp5_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:08:40 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_XOR2XP5_ASAP7_75T_R%A 2 5 7 10 13 15 25 26 29 33 38 39 40 42 44 46 49
+ 53 54 VSS
c37 54 VSS 0.00752343f $X=0.018 $Y=0.135
c38 53 VSS 6.31991e-19 $X=0.351 $Y=0.169
c39 49 VSS 4.77226e-19 $X=0.351 $Y=0.135
c40 47 VSS 9.00374e-19 $X=0.351 $Y=0.189
c41 46 VSS 2.41739e-19 $X=0.299 $Y=0.198
c42 45 VSS 0.00174705f $X=0.256 $Y=0.198
c43 44 VSS 1.80165e-19 $X=0.225 $Y=0.198
c44 43 VSS 0.00292169f $X=0.342 $Y=0.198
c45 42 VSS 6.38596e-24 $X=0.216 $Y=0.225
c46 40 VSS 0.00133719f $X=0.18 $Y=0.234
c47 39 VSS 0.00181942f $X=0.162 $Y=0.234
c48 38 VSS 0.00321912f $X=0.144 $Y=0.234
c49 37 VSS 0.00131186f $X=0.106 $Y=0.234
c50 36 VSS 0.00145201f $X=0.094 $Y=0.234
c51 35 VSS 0.00785083f $X=0.078 $Y=0.234
c52 34 VSS 0.0032309f $X=0.027 $Y=0.234
c53 33 VSS 0.00486444f $X=0.207 $Y=0.234
c54 29 VSS 0.00203697f $X=0.06 $Y=0.134
c55 26 VSS 8.69458e-19 $X=0.018 $Y=0.207
c56 25 VSS 0.00218042f $X=0.018 $Y=0.189
c57 24 VSS 6.58554e-19 $X=0.018 $Y=0.225
c58 13 VSS 0.0014523f $X=0.351 $Y=0.135
c59 10 VSS 0.0618866f $X=0.351 $Y=0.0675
c60 5 VSS 0.00581295f $X=0.081 $Y=0.135
c61 2 VSS 0.0638905f $X=0.081 $Y=0.054
r62 52 53 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.149 $X2=0.351 $Y2=0.169
r63 49 52 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.149
r64 47 53 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.189 $X2=0.351 $Y2=0.169
r65 45 46 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.198 $X2=0.299 $Y2=0.198
r66 44 45 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.198 $X2=0.256 $Y2=0.198
r67 43 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.198 $X2=0.351 $Y2=0.189
r68 43 46 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.299 $Y2=0.198
r69 41 44 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.207 $X2=0.225 $Y2=0.198
r70 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.207 $X2=0.216 $Y2=0.225
r71 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.18 $Y2=0.234
r72 38 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.162 $Y2=0.234
r73 37 38 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.106
+ $Y=0.234 $X2=0.144 $Y2=0.234
r74 36 37 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.234 $X2=0.106 $Y2=0.234
r75 35 36 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.234 $X2=0.094 $Y2=0.234
r76 34 35 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.078 $Y2=0.234
r77 33 42 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.207 $Y=0.234 $X2=0.216 $Y2=0.225
r78 33 40 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.234 $X2=0.18 $Y2=0.234
r79 29 31 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r80 27 54 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r81 27 29 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.06 $Y2=0.135
r82 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.207
r83 24 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.225 $X2=0.027 $Y2=0.234
r84 24 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.225 $X2=0.018 $Y2=0.207
r85 23 54 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r86 23 25 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.189
r87 13 49 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r88 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r89 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r90 5 31 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r91 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r92 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.054 $X2=0.081 $Y2=0.135
.ends

.subckt PM_XOR2XP5_ASAP7_75T_R%B 2 7 10 13 15 24 VSS
c33 24 VSS 0.00327325f $X=0.136 $Y=0.135
c34 13 VSS 0.0170801f $X=0.297 $Y=0.135
c35 10 VSS 0.0656969f $X=0.297 $Y=0.0675
c36 2 VSS 0.0637809f $X=0.135 $Y=0.054
r37 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r38 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r39 5 13 202.5 $w=1.6e-08 $l=1.62e-07 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.297 $Y2=0.135
r40 5 24 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r41 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r42 2 5 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.054 $X2=0.135 $Y2=0.135
.ends

.subckt PM_XOR2XP5_ASAP7_75T_R%5 2 5 7 9 10 13 14 19 26 27 29 32 33 34 35 38 40
+ 41 42 43 51 53 VSS
c40 53 VSS 0.00205152f $X=0.171 $Y=0.072
c41 51 VSS 1.15487e-19 $X=0.405 $Y=0.1275
c42 50 VSS 0.00161525f $X=0.405 $Y=0.12
c43 48 VSS 2.98192e-19 $X=0.405 $Y=0.135
c44 45 VSS 1.56568e-19 $X=0.3915 $Y=0.072
c45 44 VSS 0.00218422f $X=0.387 $Y=0.072
c46 43 VSS 8.46035e-21 $X=0.36 $Y=0.072
c47 42 VSS 9.56695e-19 $X=0.342 $Y=0.072
c48 41 VSS 0.00278191f $X=0.256 $Y=0.072
c49 40 VSS 0.00149783f $X=0.207 $Y=0.072
c50 38 VSS 7.89418e-20 $X=0.396 $Y=0.072
c51 35 VSS 5.82771e-19 $X=0.171 $Y=0.15
c52 34 VSS 9.593e-19 $X=0.171 $Y=0.12
c53 33 VSS 0.0143473f $X=0.171 $Y=0.18
c54 32 VSS 9.04725e-19 $X=0.171 $Y=0.18
c55 29 VSS 9.37882e-19 $X=0.171 $Y=0.063
c56 27 VSS 0.00150698f $X=0.153 $Y=0.036
c57 26 VSS 0.00287092f $X=0.144 $Y=0.036
c58 21 VSS 0.00259308f $X=0.108 $Y=0.036
c59 19 VSS 0.00458651f $X=0.162 $Y=0.036
c60 17 VSS 4.79286e-19 $X=0.16 $Y=0.2025
c61 13 VSS 0.00800631f $X=0.108 $Y=0.054
c62 9 VSS 6.05457e-19 $X=0.125 $Y=0.054
c63 5 VSS 0.00172734f $X=0.405 $Y=0.135
c64 2 VSS 0.0664387f $X=0.405 $Y=0.0675
r65 50 51 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.12 $X2=0.405 $Y2=0.1275
r66 48 51 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.1275
r67 46 50 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.081 $X2=0.405 $Y2=0.12
r68 44 45 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.387
+ $Y=0.072 $X2=0.3915 $Y2=0.072
r69 43 44 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.072 $X2=0.387 $Y2=0.072
r70 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.072 $X2=0.36 $Y2=0.072
r71 41 42 5.83951 $w=1.8e-08 $l=8.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.072 $X2=0.342 $Y2=0.072
r72 40 41 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.072 $X2=0.256 $Y2=0.072
r73 39 53 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.072 $X2=0.171 $Y2=0.072
r74 39 40 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.072 $X2=0.207 $Y2=0.072
r75 38 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.072 $X2=0.405 $Y2=0.081
r76 38 45 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.072 $X2=0.3915 $Y2=0.072
r77 34 35 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.12 $X2=0.171 $Y2=0.15
r78 32 35 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.18 $X2=0.171 $Y2=0.15
r79 32 33 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.171 $Y=0.18 $X2=0.171
+ $Y2=0.18
r80 30 53 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.081 $X2=0.171 $Y2=0.072
r81 30 34 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.081 $X2=0.171 $Y2=0.12
r82 29 53 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.063 $X2=0.171 $Y2=0.072
r83 28 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.045 $X2=0.171 $Y2=0.063
r84 26 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.153 $Y2=0.036
r85 21 26 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.144 $Y2=0.036
r86 19 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.036 $X2=0.171 $Y2=0.045
r87 19 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.153 $Y2=0.036
r88 17 33 9.51166 $w=4.9e-08 $l=2.25e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.1745 $Y=0.2025 $X2=0.1745 $Y2=0.18
r89 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.2025 $X2=0.16 $Y2=0.2025
r90 13 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r91 10 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.054 $X2=0.108 $Y2=0.054
r92 9 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.054 $X2=0.108 $Y2=0.054
r93 5 48 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r94 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r95 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_XOR2XP5_ASAP7_75T_R%Y 1 6 11 14 19 23 24 29 31 33 39 VSS
c18 39 VSS 0.00328191f $X=0.45 $Y=0.234
c19 38 VSS 0.00277971f $X=0.459 $Y=0.234
c20 33 VSS 0.00258114f $X=0.459 $Y=0.207
c21 31 VSS 0.00142966f $X=0.459 $Y=0.099
c22 30 VSS 5.7946e-19 $X=0.459 $Y=0.063
c23 29 VSS 0.00223776f $X=0.457 $Y=0.135
c24 27 VSS 0.00102822f $X=0.459 $Y=0.225
c25 25 VSS 8.76814e-19 $X=0.423 $Y=0.036
c26 24 VSS 0.0161022f $X=0.414 $Y=0.036
c27 23 VSS 0.00677526f $X=0.432 $Y=0.036
c28 19 VSS 0.00505246f $X=0.27 $Y=0.036
c29 16 VSS 0.00607607f $X=0.45 $Y=0.036
c30 14 VSS 0.00327032f $X=0.43 $Y=0.2025
c31 9 VSS 2.69461e-19 $X=0.43 $Y=0.0675
c32 1 VSS 4.39464e-19 $X=0.287 $Y=0.0675
r33 39 40 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.4545 $Y2=0.234
r34 38 40 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.234 $X2=0.4545 $Y2=0.234
r35 35 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.45 $Y2=0.234
r36 32 33 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.149 $X2=0.459 $Y2=0.207
r37 30 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.063 $X2=0.459 $Y2=0.099
r38 29 32 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.149
r39 29 31 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.099
r40 27 38 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.234
r41 27 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.207
r42 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.063
r43 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.423 $Y2=0.036
r44 22 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.423 $Y2=0.036
r45 22 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r46 18 24 9.77778 $w=1.8e-08 $l=1.44e-07 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.414 $Y2=0.036
r47 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r48 16 26 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r49 16 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.432 $Y2=0.036
r50 14 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r51 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.43 $Y2=0.2025
r52 9 23 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r53 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.43 $Y2=0.0675
r54 4 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r55 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.272 $Y2=0.0675
.ends

.subckt PM_XOR2XP5_ASAP7_75T_R%9 1 2 VSS
c1 1 VSS 0.00224058f $X=0.125 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.091 $Y2=0.2025
.ends


* END of "./XOR2xp5_ASAP7_75t_R.pex.sp.pex"
* 
.subckt XOR2xp5_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 N_5_M0_d N_A_M0_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.027
M1 VSS N_B_M1_g N_5_M1_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.027
M2 noxref_8 N_B_M2_g N_Y_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M3 VSS N_A_M3_g noxref_8 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M4 N_Y_M4_d N_5_M4_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M5 N_9_M5_d N_A_M5_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M6 N_5_M6_d N_B_M6_g N_9_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M7 VDD N_B_M7_g noxref_6 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.162
M8 noxref_6 N_A_M8_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.162
M9 N_Y_M9_d N_5_M9_g noxref_6 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
*
* 
* .include "XOR2xp5_ASAP7_75t_R.pex.sp.XOR2XP5_ASAP7_75T_R.pxi"
* BEGIN of "./XOR2xp5_ASAP7_75t_R.pex.sp.XOR2XP5_ASAP7_75T_R.pxi"
* File: XOR2xp5_ASAP7_75t_R.pex.sp.XOR2XP5_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:08:40 2017
* 
x_PM_XOR2XP5_ASAP7_75T_R%A N_A_M0_g N_A_c_5_p N_A_M5_g N_A_M3_g N_A_c_6_p
+ N_A_M8_g N_A_c_9_p N_A_c_10_p A N_A_c_7_p N_A_c_2_p N_A_c_21_p N_A_c_18_p
+ N_A_c_30_p N_A_c_8_p N_A_c_4_p N_A_c_27_p N_A_c_32_p N_A_c_14_p VSS
+ PM_XOR2XP5_ASAP7_75T_R%A
x_PM_XOR2XP5_ASAP7_75T_R%B N_B_M1_g N_B_M6_g N_B_M2_g N_B_c_42_n N_B_M7_g B VSS
+ PM_XOR2XP5_ASAP7_75T_R%B
x_PM_XOR2XP5_ASAP7_75T_R%5 N_5_M4_g N_5_c_72_n N_5_M9_g N_5_M1_s N_5_M0_d
+ N_5_c_86_n N_5_M6_d N_5_c_106_p N_5_c_87_n N_5_c_89_n N_5_c_73_n N_5_c_74_n
+ N_5_c_76_n N_5_c_93_n N_5_c_94_n N_5_c_104_p N_5_c_96_n N_5_c_80_n N_5_c_81_n
+ N_5_c_82_n N_5_c_84_n N_5_c_98_n VSS PM_XOR2XP5_ASAP7_75T_R%5
x_PM_XOR2XP5_ASAP7_75T_R%Y N_Y_M2_s N_Y_M4_d N_Y_M9_d N_Y_c_125_n N_Y_c_113_n
+ N_Y_c_119_n N_Y_c_111_n Y N_Y_c_124_n N_Y_c_112_n N_Y_c_127_n VSS
+ PM_XOR2XP5_ASAP7_75T_R%Y
x_PM_XOR2XP5_ASAP7_75T_R%9 N_9_M6_s N_9_M5_d VSS PM_XOR2XP5_ASAP7_75T_R%9
cc_1 N_A_M0_g N_B_M1_g 0.00344695f $X=0.081 $Y=0.054 $X2=0.135 $Y2=0.054
cc_2 N_A_c_2_p N_B_M1_g 2.38942e-19 $X=0.144 $Y=0.234 $X2=0.135 $Y2=0.054
cc_3 N_A_M3_g N_B_M2_g 0.00323392f $X=0.351 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_4 N_A_c_4_p N_B_M2_g 2.45429e-19 $X=0.299 $Y=0.198 $X2=0.297 $Y2=0.0675
cc_5 N_A_c_5_p N_B_c_42_n 8.12544e-19 $X=0.081 $Y=0.135 $X2=0.297 $Y2=0.135
cc_6 N_A_c_6_p N_B_c_42_n 0.00106649f $X=0.351 $Y=0.135 $X2=0.297 $Y2=0.135
cc_7 N_A_c_7_p N_B_c_42_n 3.32907e-19 $X=0.207 $Y=0.234 $X2=0.297 $Y2=0.135
cc_8 N_A_c_8_p N_B_c_42_n 0.00124812f $X=0.225 $Y=0.198 $X2=0.297 $Y2=0.135
cc_9 N_A_c_9_p B 2.55557e-19 $X=0.018 $Y=0.189 $X2=0.136 $Y2=0.135
cc_10 N_A_c_10_p B 2.38976e-19 $X=0.018 $Y=0.207 $X2=0.136 $Y2=0.135
cc_11 A B 4.29558e-19 $X=0.06 $Y=0.134 $X2=0.136 $Y2=0.135
cc_12 N_A_c_2_p B 0.00409303f $X=0.144 $Y=0.234 $X2=0.136 $Y2=0.135
cc_13 N_A_c_8_p B 3.31105e-19 $X=0.225 $Y=0.198 $X2=0.136 $Y2=0.135
cc_14 N_A_c_14_p B 8.14212e-19 $X=0.018 $Y=0.135 $X2=0.136 $Y2=0.135
cc_15 N_A_M3_g N_5_M4_g 0.00323392f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.054
cc_16 N_A_c_6_p N_5_c_72_n 9.46013e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_17 N_A_c_14_p N_5_c_73_n 2.72061e-19 $X=0.018 $Y=0.135 $X2=0 $Y2=0
cc_18 N_A_c_18_p N_5_c_74_n 8.69266e-19 $X=0.18 $Y=0.234 $X2=0.135 $Y2=0.135
cc_19 N_A_c_8_p N_5_c_74_n 3.18815e-19 $X=0.225 $Y=0.198 $X2=0.135 $Y2=0.135
cc_20 N_A_c_7_p N_5_c_76_n 0.00142006f $X=0.207 $Y=0.234 $X2=0 $Y2=0
cc_21 N_A_c_21_p N_5_c_76_n 0.00161143f $X=0.162 $Y=0.234 $X2=0 $Y2=0
cc_22 N_A_c_18_p N_5_c_76_n 0.00130888f $X=0.18 $Y=0.234 $X2=0 $Y2=0
cc_23 N_A_c_8_p N_5_c_76_n 7.82924e-19 $X=0.225 $Y=0.198 $X2=0 $Y2=0
cc_24 N_A_c_8_p N_5_c_80_n 7.71444e-19 $X=0.225 $Y=0.198 $X2=0 $Y2=0
cc_25 N_A_c_4_p N_5_c_81_n 7.71444e-19 $X=0.299 $Y=0.198 $X2=0 $Y2=0
cc_26 N_A_M3_g N_5_c_82_n 3.0688e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_A_c_27_p N_5_c_82_n 8.07817e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_28 N_A_c_27_p N_5_c_84_n 0.00118961f $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_29 VSS N_A_c_4_p 3.29233e-19 $X=0.299 $Y=0.198 $X2=0.135 $Y2=0.054
cc_30 VSS N_A_c_30_p 6.7861e-19 $X=0.216 $Y=0.225 $X2=0.135 $Y2=0.135
cc_31 VSS N_A_c_4_p 0.00219077f $X=0.299 $Y=0.198 $X2=0.135 $Y2=0.135
cc_32 VSS N_A_c_32_p 0.00157748f $X=0.351 $Y=0.169 $X2=0.297 $Y2=0.0675
cc_33 VSS N_A_M3_g 2.34993e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_34 VSS N_A_c_7_p 0.00123555f $X=0.207 $Y=0.234 $X2=0 $Y2=0
cc_35 VSS N_A_c_4_p 0.00880208f $X=0.299 $Y=0.198 $X2=0 $Y2=0
cc_36 N_A_M3_g N_Y_c_111_n 2.38303e-19 $X=0.351 $Y=0.0675 $X2=0.136 $Y2=0.135
cc_37 N_A_c_32_p N_Y_c_112_n 6.04755e-19 $X=0.351 $Y=0.169 $X2=0 $Y2=0
cc_38 N_B_M2_g N_5_M4_g 2.34385e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.054
cc_39 B N_5_c_86_n 0.00184579f $X=0.136 $Y=0.135 $X2=0.351 $Y2=0.135
cc_40 N_B_M1_g N_5_c_87_n 2.35623e-19 $X=0.135 $Y=0.054 $X2=0.018 $Y2=0.207
cc_41 B N_5_c_87_n 0.00374777f $X=0.136 $Y=0.135 $X2=0.018 $Y2=0.207
cc_42 N_B_c_42_n N_5_c_89_n 2.91977e-19 $X=0.297 $Y=0.135 $X2=0.027 $Y2=0.135
cc_43 B N_5_c_74_n 0.0044259f $X=0.136 $Y=0.135 $X2=0 $Y2=0
cc_44 N_B_c_42_n N_5_c_76_n 0.00369057f $X=0.297 $Y=0.135 $X2=0.207 $Y2=0.234
cc_45 B N_5_c_76_n 5.02969e-19 $X=0.136 $Y=0.135 $X2=0.207 $Y2=0.234
cc_46 B N_5_c_93_n 0.00221295f $X=0.136 $Y=0.135 $X2=0.027 $Y2=0.234
cc_47 N_B_c_42_n N_5_c_94_n 0.00250832f $X=0.297 $Y=0.135 $X2=0.078 $Y2=0.234
cc_48 B N_5_c_94_n 0.00221295f $X=0.136 $Y=0.135 $X2=0.078 $Y2=0.234
cc_49 N_B_c_42_n N_5_c_96_n 0.00135939f $X=0.297 $Y=0.135 $X2=0.18 $Y2=0.234
cc_50 N_B_M2_g N_5_c_81_n 4.09048e-19 $X=0.297 $Y=0.0675 $X2=0.216 $Y2=0.225
cc_51 B N_5_c_98_n 0.00221295f $X=0.136 $Y=0.135 $X2=0.351 $Y2=0.169
cc_52 VSS N_B_c_42_n 6.8292e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_53 VSS N_B_M2_g 2.65491e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_54 N_B_c_42_n N_Y_c_113_n 6.8292e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_55 N_B_M2_g N_Y_c_111_n 2.65491e-19 $X=0.297 $Y=0.0675 $X2=0.018 $Y2=0.225
cc_56 B N_9_M6_s 2.00044e-19 $X=0.136 $Y=0.135 $X2=0.081 $Y2=0.054
cc_57 VSS N_5_c_76_n 0.00221794f $X=0.171 $Y=0.18 $X2=0.081 $Y2=0.135
cc_58 N_5_c_81_n N_Y_M2_s 3.29233e-19 $X=0.342 $Y=0.072 $X2=0.081 $Y2=0.054
cc_59 N_5_c_73_n N_Y_c_113_n 2.38811e-19 $X=0.171 $Y=0.063 $X2=0 $Y2=0
cc_60 N_5_c_93_n N_Y_c_113_n 5.58422e-19 $X=0.171 $Y=0.12 $X2=0 $Y2=0
cc_61 N_5_c_81_n N_Y_c_113_n 0.00284111f $X=0.342 $Y=0.072 $X2=0 $Y2=0
cc_62 N_5_c_104_p N_Y_c_119_n 0.00136624f $X=0.396 $Y=0.072 $X2=0.018 $Y2=0.144
cc_63 N_5_M4_g N_Y_c_111_n 2.34993e-19 $X=0.405 $Y=0.0675 $X2=0.018 $Y2=0.225
cc_64 N_5_c_106_p N_Y_c_111_n 5.49907e-19 $X=0.162 $Y=0.036 $X2=0.018 $Y2=0.225
cc_65 N_5_c_81_n N_Y_c_111_n 0.0133208f $X=0.342 $Y=0.072 $X2=0.018 $Y2=0.225
cc_66 N_5_c_84_n Y 0.00172057f $X=0.405 $Y=0.1275 $X2=0.06 $Y2=0.134
cc_67 N_5_c_104_p N_Y_c_124_n 0.00172057f $X=0.396 $Y=0.072 $X2=0.064 $Y2=0.135
cc_68 VSS N_5_c_81_n 5.15356e-19 $X=0.342 $Y=0.072 $X2=0.081 $Y2=0.054
cc_69 VSS N_Y_c_125_n 0.00395939f $X=0.378 $Y=0.2025 $X2=0.351 $Y2=0.2025
cc_70 VSS N_Y_c_113_n 0.00169333f $X=0.272 $Y=0.2025 $X2=0 $Y2=0
cc_71 VSS N_Y_c_127_n 6.5272e-19 $X=0.378 $Y=0.234 $X2=0.162 $Y2=0.234
cc_72 VSS N_Y_c_111_n 3.33359e-19 $X=0.414 $Y=0.036 $X2=0.081 $Y2=0.054

* END of "./XOR2xp5_ASAP7_75t_R.pex.sp.XOR2XP5_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: XNOR2x1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:06:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "XNOR2x1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./XNOR2x1_ASAP7_75t_R.pex.sp.pex"
* File: XNOR2x1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:06:48 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_XNOR2X1_ASAP7_75T_R%B 2 5 7 10 13 15 18 21 23 34 38 39 40 41 42 43 46
+ 51 52 53 55 58 59 60 62 65 71 72 83 92 VSS
c63 92 VSS 9.19488e-20 $X=0.513 $Y=0.128
c64 83 VSS 1.58347e-19 $X=0.513 $Y=0.135
c65 72 VSS 0.00258863f $X=0.513 $Y=0.081
c66 71 VSS 0.00559875f $X=0.513 $Y=0.081
c67 65 VSS 0.00770297f $X=0.018 $Y=0.135
c68 62 VSS 6.41874e-19 $X=0.351 $Y=0.135
c69 60 VSS 1.40425e-19 $X=0.323 $Y=0.135
c70 59 VSS 0.00137518f $X=0.314 $Y=0.121
c71 58 VSS 7.51698e-19 $X=0.314 $Y=0.095
c72 57 VSS 4.26488e-19 $X=0.314 $Y=0.126
c73 56 VSS 0.00161475f $X=0.314 $Y=0.085
c74 55 VSS 1.57364e-19 $X=0.2805 $Y=0.076
c75 54 VSS 0.00137179f $X=0.256 $Y=0.076
c76 53 VSS 3.79724e-19 $X=0.231 $Y=0.076
c77 52 VSS 1.68167e-19 $X=0.305 $Y=0.076
c78 51 VSS 2.80979e-20 $X=0.222 $Y=0.067
c79 46 VSS 0.00238557f $X=0.06 $Y=0.136
c80 43 VSS 0.00102062f $X=0.2025 $Y=0.036
c81 42 VSS 0.00132447f $X=0.192 $Y=0.036
c82 41 VSS 0.00269371f $X=0.174 $Y=0.036
c83 40 VSS 0.00142972f $X=0.144 $Y=0.036
c84 39 VSS 0.00192708f $X=0.126 $Y=0.036
c85 38 VSS 0.00156636f $X=0.107 $Y=0.036
c86 37 VSS 0.00122076f $X=0.092 $Y=0.036
c87 36 VSS 0.0075732f $X=0.078 $Y=0.036
c88 35 VSS 0.00323226f $X=0.027 $Y=0.036
c89 34 VSS 0.00322347f $X=0.213 $Y=0.036
c90 28 VSS 0.00210014f $X=0.018 $Y=0.121
c91 27 VSS 0.00169007f $X=0.018 $Y=0.082
c92 26 VSS 1.95142e-19 $X=0.018 $Y=0.126
c93 21 VSS 0.00101384f $X=0.513 $Y=0.135
c94 18 VSS 0.0608664f $X=0.513 $Y=0.0675
c95 13 VSS 0.00143642f $X=0.351 $Y=0.135
c96 10 VSS 0.0612409f $X=0.351 $Y=0.0675
c97 5 VSS 0.00625786f $X=0.081 $Y=0.135
c98 2 VSS 0.0638905f $X=0.081 $Y=0.0675
r99 91 92 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.121 $X2=0.513 $Y2=0.128
r100 83 92 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.128
r101 72 91 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.081 $X2=0.513 $Y2=0.121
r102 71 72 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.513 $Y=0.081 $X2=0.513
+ $Y2=0.081
r103 67 71 13.5123 $w=1.8e-08 $l=1.99e-07 $layer=M2 $thickness=3.6e-08 $X=0.314
+ $Y=0.081 $X2=0.513 $Y2=0.081
r104 67 68 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.314 $Y=0.081 $X2=0.314
+ $Y2=0.081
r105 60 62 1.90123 $w=1.8e-08 $l=2.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.323
+ $Y=0.135 $X2=0.351 $Y2=0.135
r106 58 59 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.314
+ $Y=0.095 $X2=0.314 $Y2=0.121
r107 57 60 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.314 $Y=0.126 $X2=0.323 $Y2=0.135
r108 57 59 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.314
+ $Y=0.126 $X2=0.314 $Y2=0.121
r109 56 68 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.314
+ $Y=0.085 $X2=0.314 $Y2=0.076
r110 56 58 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.314
+ $Y=0.085 $X2=0.314 $Y2=0.095
r111 54 55 1.66358 $w=1.8e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.076 $X2=0.2805 $Y2=0.076
r112 53 54 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.231
+ $Y=0.076 $X2=0.256 $Y2=0.076
r113 52 68 0.341445 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.305
+ $Y=0.076 $X2=0.314 $Y2=0.076
r114 52 55 1.66358 $w=1.8e-08 $l=2.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.305
+ $Y=0.076 $X2=0.2805 $Y2=0.076
r115 51 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.222 $Y=0.067 $X2=0.231 $Y2=0.076
r116 50 51 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.222
+ $Y=0.045 $X2=0.222 $Y2=0.067
r117 46 48 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r118 44 65 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r119 44 46 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.06 $Y2=0.135
r120 42 43 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.192
+ $Y=0.036 $X2=0.2025 $Y2=0.036
r121 41 42 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.174
+ $Y=0.036 $X2=0.192 $Y2=0.036
r122 40 41 2.03704 $w=1.8e-08 $l=3e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.174 $Y2=0.036
r123 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.144 $Y2=0.036
r124 38 39 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.107
+ $Y=0.036 $X2=0.126 $Y2=0.036
r125 37 38 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.092
+ $Y=0.036 $X2=0.107 $Y2=0.036
r126 36 37 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.036 $X2=0.092 $Y2=0.036
r127 35 36 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.078 $Y2=0.036
r128 34 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.213 $Y=0.036 $X2=0.222 $Y2=0.045
r129 34 43 0.712963 $w=1.8e-08 $l=1.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.213
+ $Y=0.036 $X2=0.2025 $Y2=0.036
r130 27 28 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.082 $X2=0.018 $Y2=0.121
r131 26 65 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.135
r132 26 28 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.121
r133 25 35 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r134 25 27 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.082
r135 21 83 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r136 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r137 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r138 13 62 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r139 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.135 $X2=0.351 $Y2=0.2025
r140 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.351 $Y=0.0675 $X2=0.351 $Y2=0.135
r141 5 48 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r142 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r143 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_XNOR2X1_ASAP7_75T_R%A 2 7 10 13 15 18 21 23 27 33 36 40 43 46 48 49
+ 50 51 VSS
c65 51 VSS 0.00555131f $X=0.527 $Y=0.189
c66 50 VSS 0.00750476f $X=0.298 $Y=0.189
c67 49 VSS 9.03934e-19 $X=0.567 $Y=0.189
c68 48 VSS 0.00230547f $X=0.567 $Y=0.189
c69 43 VSS 0.00192743f $X=0.135 $Y=0.189
c70 40 VSS 3.99651e-19 $X=0.567 $Y=0.1705
c71 36 VSS 2.08027e-19 $X=0.567 $Y=0.135
c72 33 VSS 3.21653e-19 $X=0.135 $Y=0.1665
c73 27 VSS 2.96695e-19 $X=0.135 $Y=0.135
c74 21 VSS 0.00214256f $X=0.567 $Y=0.135
c75 18 VSS 0.0661499f $X=0.567 $Y=0.0675
c76 13 VSS 0.0184971f $X=0.297 $Y=0.135
c77 10 VSS 0.0656751f $X=0.297 $Y=0.0675
c78 2 VSS 0.0639533f $X=0.135 $Y=0.0675
r79 50 51 15.5494 $w=1.8e-08 $l=2.29e-07 $layer=M2 $thickness=3.6e-08 $X=0.298
+ $Y=0.189 $X2=0.527 $Y2=0.189
r80 48 51 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.567
+ $Y=0.189 $X2=0.527 $Y2=0.189
r81 48 49 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.567 $Y=0.189 $X2=0.567
+ $Y2=0.189
r82 46 50 5.6358 $w=1.8e-08 $l=8.3e-08 $layer=M2 $thickness=3.6e-08 $X=0.215
+ $Y=0.189 $X2=0.298 $Y2=0.189
r83 42 46 5.4321 $w=1.8e-08 $l=8e-08 $layer=M2 $thickness=3.6e-08 $X=0.135
+ $Y=0.189 $X2=0.215 $Y2=0.189
r84 42 43 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.135 $Y=0.189 $X2=0.135
+ $Y2=0.189
r85 40 49 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.1705 $X2=0.567 $Y2=0.189
r86 39 40 1.25617 $w=1.8e-08 $l=1.85e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.152 $X2=0.567 $Y2=0.1705
r87 36 39 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.152
r88 33 43 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.1665 $X2=0.135 $Y2=0.189
r89 32 33 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.144 $X2=0.135 $Y2=0.1665
r90 27 32 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.144
r91 21 36 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r92 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r93 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r94 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r95 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r96 5 13 202.5 $w=1.6e-08 $l=1.62e-07 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.297 $Y2=0.135
r97 5 27 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r98 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r99 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_XNOR2X1_ASAP7_75T_R%5 2 7 10 13 15 17 20 22 23 26 27 34 35 36 38 44
+ 46 47 49 50 51 52 53 55 61 62 VSS
c63 62 VSS 0.0012649f $X=0.1835 $Y=0.198
c64 61 VSS 4.92178e-19 $X=0.405 $Y=0.1665
c65 55 VSS 3.22958e-19 $X=0.405 $Y=0.135
c66 53 VSS 9.46817e-19 $X=0.405 $Y=0.189
c67 52 VSS 1.01588e-19 $X=0.365 $Y=0.198
c68 51 VSS 3.21516e-19 $X=0.305 $Y=0.198
c69 50 VSS 0.00264353f $X=0.256 $Y=0.198
c70 49 VSS 0.00102041f $X=0.213 $Y=0.198
c71 47 VSS 0.00225686f $X=0.396 $Y=0.198
c72 46 VSS 6.74689e-19 $X=0.1835 $Y=0.225
c73 44 VSS 3.45913e-19 $X=0.183 $Y=0.144
c74 38 VSS 0.0018536f $X=0.183 $Y=0.096
c75 36 VSS 0.0018106f $X=0.183 $Y=0.189
c76 35 VSS 0.0024907f $X=0.159 $Y=0.234
c77 34 VSS 0.00286142f $X=0.144 $Y=0.234
c78 29 VSS 0.0027761f $X=0.108 $Y=0.234
c79 27 VSS 0.00524826f $X=0.174 $Y=0.234
c80 26 VSS 0.0102544f $X=0.108 $Y=0.2025
c81 22 VSS 5.72255e-19 $X=0.125 $Y=0.2025
c82 20 VSS 0.0136365f $X=0.16 $Y=0.0675
c83 13 VSS 0.00334187f $X=0.459 $Y=0.135
c84 10 VSS 0.0625141f $X=0.459 $Y=0.0675
c85 2 VSS 0.0619268f $X=0.405 $Y=0.0675
r86 60 61 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.144 $X2=0.405 $Y2=0.1665
r87 55 60 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.144
r88 53 61 1.52778 $w=1.8e-08 $l=2.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.1665
r89 51 52 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.305
+ $Y=0.198 $X2=0.365 $Y2=0.198
r90 50 51 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.198 $X2=0.305 $Y2=0.198
r91 49 50 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.213
+ $Y=0.198 $X2=0.256 $Y2=0.198
r92 48 62 0.144403 $w=3.7e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.193
+ $Y=0.198 $X2=0.1835 $Y2=0.198
r93 48 49 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.193
+ $Y=0.198 $X2=0.213 $Y2=0.198
r94 47 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.198 $X2=0.405 $Y2=0.189
r95 47 52 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.365 $Y2=0.198
r96 45 62 0.505846 $w=1.9e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.1835
+ $Y=0.207 $X2=0.1835 $Y2=0.198
r97 45 46 1.14327 $w=1.9e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.1835
+ $Y=0.207 $X2=0.1835 $Y2=0.225
r98 43 44 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.183
+ $Y=0.121 $X2=0.183 $Y2=0.144
r99 38 43 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.183
+ $Y=0.096 $X2=0.183 $Y2=0.121
r100 36 62 0.505846 $w=1.9e-08 $l=9.24662e-09 $layer=M1 $thickness=3.6e-08
+ $X=0.183 $Y=0.189 $X2=0.1835 $Y2=0.198
r101 36 44 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.183
+ $Y=0.189 $X2=0.183 $Y2=0.144
r102 34 35 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.159 $Y2=0.234
r103 29 34 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.144 $Y2=0.234
r104 27 46 0.68354 $w=1.9e-08 $l=1.32571e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.174 $Y=0.234 $X2=0.1835 $Y2=0.225
r105 27 35 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.174
+ $Y=0.234 $X2=0.159 $Y2=0.234
r106 26 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234
+ $X2=0.108 $Y2=0.234
r107 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r108 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r109 20 38 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.183 $Y=0.096
+ $X2=0.183 $Y2=0.096
r110 17 20 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.16 $Y2=0.0675
r111 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r112 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r113 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r114 5 55 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r115 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r116 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_XNOR2X1_ASAP7_75T_R%Y 1 2 5 6 9 11 12 15 16 19 29 30 34 35 36 38 43
+ 44 46 53 54 VSS
c51 57 VSS 0.00176645f $X=0.459 $Y=0.234
c52 54 VSS 4.50279e-19 $X=0.45 $Y=0.086
c53 53 VSS 2.6023e-19 $X=0.459 $Y=0.086
c54 46 VSS 0.00425279f $X=0.576 $Y=0.234
c55 45 VSS 4.0861e-19 $X=0.526 $Y=0.234
c56 44 VSS 0.00147038f $X=0.522 $Y=0.234
c57 43 VSS 0.0062512f $X=0.504 $Y=0.234
c58 41 VSS 0.00513487f $X=0.594 $Y=0.234
c59 38 VSS 6.8211e-19 $X=0.459 $Y=0.207
c60 36 VSS 1.37072e-19 $X=0.459 $Y=0.152
c61 35 VSS 4.74957e-19 $X=0.459 $Y=0.121
c62 34 VSS 0.00108231f $X=0.457 $Y=0.178
c63 32 VSS 8.65169e-19 $X=0.459 $Y=0.225
c64 30 VSS 5.32692e-19 $X=0.418 $Y=0.234
c65 29 VSS 0.016166f $X=0.414 $Y=0.234
c66 21 VSS 0.00269031f $X=0.45 $Y=0.234
c67 19 VSS 0.00386033f $X=0.592 $Y=0.2025
c68 15 VSS 0.011938f $X=0.432 $Y=0.2025
c69 11 VSS 5.25448e-19 $X=0.449 $Y=0.2025
c70 9 VSS 0.00600583f $X=0.272 $Y=0.2025
c71 6 VSS 4.39464e-19 $X=0.287 $Y=0.2025
c72 5 VSS 0.00327881f $X=0.432 $Y=0.0675
c73 1 VSS 5.83596e-19 $X=0.449 $Y=0.0675
r74 54 55 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.086 $X2=0.4545 $Y2=0.086
r75 53 55 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.086 $X2=0.4545 $Y2=0.086
r76 50 54 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.086 $X2=0.45 $Y2=0.086
r77 45 46 3.39506 $w=1.8e-08 $l=5e-08 $layer=M1 $thickness=3.6e-08 $X=0.526
+ $Y=0.234 $X2=0.576 $Y2=0.234
r78 44 45 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.522
+ $Y=0.234 $X2=0.526 $Y2=0.234
r79 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.504
+ $Y=0.234 $X2=0.522 $Y2=0.234
r80 41 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.594
+ $Y=0.234 $X2=0.576 $Y2=0.234
r81 39 57 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.459 $Y2=0.234
r82 39 43 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.504 $Y2=0.234
r83 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.189 $X2=0.459 $Y2=0.207
r84 35 36 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.121 $X2=0.459 $Y2=0.152
r85 34 37 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.178 $X2=0.459 $Y2=0.189
r86 34 36 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.178 $X2=0.459 $Y2=0.152
r87 32 57 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.234
r88 32 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.207
r89 31 53 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.095 $X2=0.459 $Y2=0.086
r90 31 35 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.095 $X2=0.459 $Y2=0.121
r91 29 30 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.418 $Y2=0.234
r92 27 30 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.418 $Y2=0.234
r93 23 29 9.77778 $w=1.8e-08 $l=1.44e-07 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.414 $Y2=0.234
r94 21 57 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.459 $Y2=0.234
r95 21 27 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.432 $Y2=0.234
r96 19 41 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.594 $Y=0.234 $X2=0.594
+ $Y2=0.234
r97 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.577 $Y=0.2025 $X2=0.592 $Y2=0.2025
r98 15 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r99 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.432 $Y2=0.2025
r100 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.2025 $X2=0.432 $Y2=0.2025
r101 9 23 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r102 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.272 $Y2=0.2025
r103 5 50 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.086 $X2=0.432
+ $Y2=0.086
r104 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.0675 $X2=0.432 $Y2=0.0675
r105 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.449 $Y=0.0675 $X2=0.432 $Y2=0.0675
.ends

.subckt PM_XNOR2X1_ASAP7_75T_R%8 1 2 VSS
c2 1 VSS 0.00180539f $X=0.125 $Y=0.0675
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends


* END of "./XNOR2x1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt XNOR2x1_ASAP7_75t_R  VSS VDD B A Y
* 
* Y	Y
* A	A
* B	B
M0 N_8_M0_d N_B_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_5_M1_d N_A_M1_g N_8_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_A_M2_g noxref_6 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M3 noxref_6 N_B_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M4 N_Y_M4_d N_5_M4_g noxref_6 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 N_Y_M5_d N_5_M5_g noxref_6 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M6 noxref_6 N_B_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M7 VSS N_A_M7_g noxref_6 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557 $Y=0.027
M8 N_5_M8_d N_B_M8_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M9 VDD N_A_M9_g N_5_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M10 N_Y_M10_d N_A_M10_g noxref_9 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M11 noxref_9 N_B_M11_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M12 N_Y_M12_d N_5_M12_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M13 N_Y_M13_d N_5_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M14 noxref_10 N_B_M14_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
M15 N_Y_M15_d N_A_M15_g noxref_10 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
*
* 
* .include "XNOR2x1_ASAP7_75t_R.pex.sp.XNOR2X1_ASAP7_75T_R.pxi"
* BEGIN of "./XNOR2x1_ASAP7_75t_R.pex.sp.XNOR2X1_ASAP7_75T_R.pxi"
* File: XNOR2x1_ASAP7_75t_R.pex.sp.XNOR2X1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:06:48 2017
* 
x_PM_XNOR2X1_ASAP7_75T_R%B N_B_M0_g N_B_c_6_p N_B_M8_g N_B_M3_g N_B_c_7_p
+ N_B_M11_g N_B_M6_g N_B_c_12_p N_B_M14_g N_B_c_43_p N_B_c_61_p N_B_c_62_p
+ N_B_c_2_p N_B_c_8_p N_B_c_28_p N_B_c_29_p B N_B_c_30_p N_B_c_4_p N_B_c_9_p
+ N_B_c_33_p N_B_c_41_p N_B_c_5_p N_B_c_10_p N_B_c_36_p N_B_c_15_p N_B_c_20_p
+ N_B_c_49_p N_B_c_57_p N_B_c_16_p VSS PM_XNOR2X1_ASAP7_75T_R%B
x_PM_XNOR2X1_ASAP7_75T_R%A N_A_M1_g N_A_M9_g N_A_M2_g N_A_c_69_n N_A_M10_g
+ N_A_M7_g N_A_c_75_n N_A_M15_g N_A_c_76_n N_A_c_78_n N_A_c_79_n N_A_c_116_p
+ N_A_c_89_p A N_A_c_117_p N_A_c_122_p N_A_c_80_n N_A_c_82_n VSS
+ PM_XNOR2X1_ASAP7_75T_R%A
x_PM_XNOR2X1_ASAP7_75T_R%5 N_5_M4_g N_5_M12_g N_5_M5_g N_5_c_133_n N_5_M13_g
+ N_5_M1_d N_5_c_135_n N_5_M9_s N_5_M8_d N_5_c_149_n N_5_c_183_p N_5_c_151_n
+ N_5_c_153_n N_5_c_155_n N_5_c_139_n N_5_c_157_n N_5_c_177_p N_5_c_159_n
+ N_5_c_160_n N_5_c_140_n N_5_c_141_n N_5_c_142_n N_5_c_166_n N_5_c_144_n
+ N_5_c_181_p N_5_c_167_n VSS PM_XNOR2X1_ASAP7_75T_R%5
x_PM_XNOR2X1_ASAP7_75T_R%Y N_Y_M5_d N_Y_M4_d N_Y_c_217_n N_Y_M10_d N_Y_c_201_n
+ N_Y_M13_d N_Y_M12_d N_Y_c_203_n N_Y_M15_d N_Y_c_204_n N_Y_c_192_n N_Y_c_207_n
+ Y N_Y_c_193_n N_Y_c_195_n N_Y_c_210_n N_Y_c_212_n N_Y_c_196_n N_Y_c_213_n
+ N_Y_c_198_n N_Y_c_200_n VSS PM_XNOR2X1_ASAP7_75T_R%Y
x_PM_XNOR2X1_ASAP7_75T_R%8 N_8_M1_s N_8_M0_d VSS PM_XNOR2X1_ASAP7_75T_R%8
cc_1 N_B_M0_g N_A_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_B_c_2_p N_A_M1_g 3.72893e-19 $X=0.144 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_3 N_B_M3_g N_A_M2_g 0.00323392f $X=0.351 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_4 N_B_c_4_p N_A_M2_g 3.987e-19 $X=0.305 $Y=0.076 $X2=0.297 $Y2=0.0675
cc_5 N_B_c_5_p N_A_M2_g 3.81992e-19 $X=0.314 $Y=0.121 $X2=0.297 $Y2=0.0675
cc_6 N_B_c_6_p N_A_c_69_n 8.12544e-19 $X=0.081 $Y=0.135 $X2=0.297 $Y2=0.135
cc_7 N_B_c_7_p N_A_c_69_n 0.00113906f $X=0.351 $Y=0.135 $X2=0.297 $Y2=0.135
cc_8 N_B_c_8_p N_A_c_69_n 2.65814e-19 $X=0.174 $Y=0.036 $X2=0.297 $Y2=0.135
cc_9 N_B_c_9_p N_A_c_69_n 0.0010895f $X=0.231 $Y=0.076 $X2=0.297 $Y2=0.135
cc_10 N_B_c_10_p N_A_c_69_n 0.00113991f $X=0.323 $Y=0.135 $X2=0.297 $Y2=0.135
cc_11 N_B_M6_g N_A_M7_g 0.00323392f $X=0.513 $Y=0.0675 $X2=0.567 $Y2=0.0675
cc_12 N_B_c_12_p N_A_c_75_n 9.33263e-19 $X=0.513 $Y=0.135 $X2=0.567 $Y2=0.135
cc_13 N_B_c_2_p N_A_c_76_n 3.94969e-19 $X=0.144 $Y=0.036 $X2=0.135 $Y2=0.135
cc_14 B N_A_c_76_n 4.29558e-19 $X=0.06 $Y=0.136 $X2=0.135 $Y2=0.135
cc_15 N_B_c_15_p N_A_c_78_n 4.74678e-19 $X=0.018 $Y=0.135 $X2=0.135 $Y2=0.1665
cc_16 N_B_c_16_p N_A_c_79_n 0.0012977f $X=0.513 $Y=0.128 $X2=0.567 $Y2=0.135
cc_17 N_B_c_8_p N_A_c_80_n 2.55398e-19 $X=0.174 $Y=0.036 $X2=0.298 $Y2=0.189
cc_18 N_B_c_9_p N_A_c_80_n 9.35543e-19 $X=0.231 $Y=0.076 $X2=0.298 $Y2=0.189
cc_19 N_B_c_10_p N_A_c_82_n 3.08473e-19 $X=0.323 $Y=0.135 $X2=0.527 $Y2=0.189
cc_20 N_B_c_20_p N_A_c_82_n 0.00480718f $X=0.513 $Y=0.081 $X2=0.527 $Y2=0.189
cc_21 N_B_M3_g N_5_M4_g 0.00323392f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_22 N_B_M6_g N_5_M4_g 2.69148e-19 $X=0.513 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_23 N_B_M3_g N_5_M5_g 2.69148e-19 $X=0.351 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_24 N_B_M6_g N_5_M5_g 0.00323392f $X=0.513 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_25 N_B_c_7_p N_5_c_133_n 0.00118234f $X=0.351 $Y=0.135 $X2=0.297 $Y2=0.135
cc_26 N_B_c_12_p N_5_c_133_n 9.33059e-19 $X=0.513 $Y=0.135 $X2=0.297 $Y2=0.135
cc_27 N_B_c_8_p N_5_c_135_n 0.00258171f $X=0.174 $Y=0.036 $X2=0.567 $Y2=0.135
cc_28 N_B_c_28_p N_5_c_135_n 0.00116706f $X=0.192 $Y=0.036 $X2=0.567 $Y2=0.135
cc_29 N_B_c_29_p N_5_c_135_n 8.50062e-19 $X=0.2025 $Y=0.036 $X2=0.567 $Y2=0.135
cc_30 N_B_c_30_p N_5_c_135_n 0.00100151f $X=0.222 $Y=0.067 $X2=0.567 $Y2=0.135
cc_31 N_B_c_28_p N_5_c_139_n 6.81694e-19 $X=0.192 $Y=0.036 $X2=0 $Y2=0
cc_32 N_B_c_9_p N_5_c_140_n 3.73122e-19 $X=0.231 $Y=0.076 $X2=0.298 $Y2=0.189
cc_33 N_B_c_33_p N_5_c_141_n 3.73122e-19 $X=0.2805 $Y=0.076 $X2=0.527 $Y2=0.189
cc_34 N_B_M3_g N_5_c_142_n 3.36975e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_35 N_B_c_10_p N_5_c_142_n 0.00215596f $X=0.323 $Y=0.135 $X2=0 $Y2=0
cc_36 N_B_c_36_p N_5_c_144_n 8.71544e-19 $X=0.351 $Y=0.135 $X2=0.297 $Y2=0.135
cc_37 VSS N_B_c_33_p 2.87556e-19 $X=0.2805 $Y=0.076 $X2=0.135 $Y2=0.0675
cc_38 VSS N_B_c_30_p 9.1988e-19 $X=0.222 $Y=0.067 $X2=0.567 $Y2=0.2025
cc_39 VSS N_B_c_4_p 4.50928e-19 $X=0.305 $Y=0.076 $X2=0.567 $Y2=0.2025
cc_40 VSS N_B_c_33_p 0.00191341f $X=0.2805 $Y=0.076 $X2=0.567 $Y2=0.2025
cc_41 VSS N_B_c_41_p 5.25032e-19 $X=0.314 $Y=0.095 $X2=0.567 $Y2=0.2025
cc_42 VSS N_B_c_20_p 3.98572e-19 $X=0.513 $Y=0.081 $X2=0.135 $Y2=0.135
cc_43 VSS N_B_c_43_p 0.00162699f $X=0.213 $Y=0.036 $X2=0.135 $Y2=0.135
cc_44 VSS N_B_c_33_p 0.00468689f $X=0.2805 $Y=0.076 $X2=0.135 $Y2=0.135
cc_45 VSS N_B_M3_g 4.26368e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_46 VSS N_B_c_36_p 4.87592e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_47 VSS N_B_c_20_p 0.00261669f $X=0.513 $Y=0.081 $X2=0 $Y2=0
cc_48 VSS N_B_c_20_p 2.66313e-19 $X=0.513 $Y=0.081 $X2=0.135 $Y2=0.144
cc_49 VSS N_B_c_49_p 0.0010042f $X=0.513 $Y=0.081 $X2=0.135 $Y2=0.144
cc_50 VSS N_B_M6_g 2.63086e-19 $X=0.513 $Y=0.0675 $X2=0.135 $Y2=0.189
cc_51 VSS N_B_c_49_p 0.00118811f $X=0.513 $Y=0.081 $X2=0.135 $Y2=0.189
cc_52 N_B_M3_g N_Y_c_192_n 2.63664e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_53 N_B_c_5_p N_Y_c_193_n 2.51979e-19 $X=0.314 $Y=0.121 $X2=0.567 $Y2=0.135
cc_54 N_B_c_49_p N_Y_c_193_n 0.0010248f $X=0.513 $Y=0.081 $X2=0.567 $Y2=0.135
cc_55 N_B_c_16_p N_Y_c_195_n 0.0010248f $X=0.513 $Y=0.128 $X2=0.567 $Y2=0.135
cc_56 N_B_M6_g N_Y_c_196_n 3.7388e-19 $X=0.513 $Y=0.0675 $X2=0 $Y2=0
cc_57 N_B_c_57_p N_Y_c_196_n 2.45728e-19 $X=0.513 $Y=0.135 $X2=0 $Y2=0
cc_58 N_B_c_20_p N_Y_c_198_n 6.12216e-19 $X=0.513 $Y=0.081 $X2=0.135 $Y2=0.135
cc_59 N_B_c_49_p N_Y_c_198_n 0.0010248f $X=0.513 $Y=0.081 $X2=0.135 $Y2=0.135
cc_60 N_B_c_20_p N_Y_c_200_n 6.55744e-19 $X=0.513 $Y=0.081 $X2=0 $Y2=0
cc_61 N_B_c_61_p N_8_M1_s 2.09605e-19 $X=0.107 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_62 N_B_c_62_p N_8_M1_s 2.34185e-19 $X=0.126 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_63 VSS N_B_c_10_p 5.39108e-19 $X=0.323 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_64 N_A_M2_g N_5_M4_g 2.34385e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_65 N_A_M7_g N_5_M5_g 2.34385e-19 $X=0.567 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_66 N_A_c_82_n N_5_c_133_n 2.36611e-19 $X=0.527 $Y=0.189 $X2=0.351 $Y2=0.135
cc_67 N_A_c_69_n N_5_c_135_n 0.00247099f $X=0.297 $Y=0.135 $X2=0.513 $Y2=0.135
cc_68 N_A_c_78_n N_5_c_149_n 8.20453e-19 $X=0.135 $Y=0.1665 $X2=0.018 $Y2=0.126
cc_69 N_A_c_89_p N_5_c_149_n 0.00122578f $X=0.135 $Y=0.189 $X2=0.018 $Y2=0.126
cc_70 N_A_M1_g N_5_c_151_n 2.34628e-19 $X=0.135 $Y=0.0675 $X2=0.213 $Y2=0.036
cc_71 N_A_c_89_p N_5_c_151_n 0.00382236f $X=0.135 $Y=0.189 $X2=0.213 $Y2=0.036
cc_72 N_A_c_69_n N_5_c_153_n 3.48111e-19 $X=0.297 $Y=0.135 $X2=0.027 $Y2=0.036
cc_73 N_A_c_80_n N_5_c_153_n 3.78066e-19 $X=0.298 $Y=0.189 $X2=0.027 $Y2=0.036
cc_74 N_A_c_76_n N_5_c_155_n 0.00148138f $X=0.135 $Y=0.135 $X2=0.078 $Y2=0.036
cc_75 N_A_c_80_n N_5_c_155_n 5.35839e-19 $X=0.298 $Y=0.189 $X2=0.078 $Y2=0.036
cc_76 N_A_c_69_n N_5_c_157_n 0.00210929f $X=0.297 $Y=0.135 $X2=0.027 $Y2=0.135
cc_77 N_A_c_76_n N_5_c_157_n 0.00148138f $X=0.135 $Y=0.135 $X2=0.027 $Y2=0.135
cc_78 N_A_c_82_n N_5_c_159_n 0.00133833f $X=0.527 $Y=0.189 $X2=0.064 $Y2=0.135
cc_79 N_A_c_69_n N_5_c_160_n 9.68215e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_80 N_A_c_80_n N_5_c_160_n 5.10242e-19 $X=0.298 $Y=0.189 $X2=0 $Y2=0
cc_81 N_A_c_80_n N_5_c_140_n 0.001214f $X=0.298 $Y=0.189 $X2=0.222 $Y2=0.045
cc_82 N_A_M2_g N_5_c_141_n 4.31042e-19 $X=0.297 $Y=0.0675 $X2=0.222 $Y2=0.067
cc_83 N_A_c_80_n N_5_c_141_n 0.00109315f $X=0.298 $Y=0.189 $X2=0.222 $Y2=0.067
cc_84 N_A_c_82_n N_5_c_142_n 0.00150184f $X=0.527 $Y=0.189 $X2=0.305 $Y2=0.076
cc_85 N_A_c_82_n N_5_c_166_n 7.13114e-19 $X=0.527 $Y=0.189 $X2=0.231 $Y2=0.076
cc_86 N_A_c_89_p N_5_c_167_n 0.00148138f $X=0.135 $Y=0.189 $X2=0.351 $Y2=0.135
cc_87 N_A_c_80_n N_5_c_167_n 3.03428e-19 $X=0.298 $Y=0.189 $X2=0.351 $Y2=0.135
cc_88 VSS N_A_c_69_n 6.8292e-19 $X=0.297 $Y=0.135 $X2=0.513 $Y2=0.2025
cc_89 VSS N_A_M2_g 2.82011e-19 $X=0.297 $Y=0.0675 $X2=0.018 $Y2=0.121
cc_90 VSS N_A_c_82_n 3.45043e-19 $X=0.527 $Y=0.189 $X2=0.2025 $Y2=0.036
cc_91 VSS N_A_M7_g 3.69259e-19 $X=0.567 $Y=0.0675 $X2=0.027 $Y2=0.135
cc_92 VSS N_A_c_79_n 3.92849e-19 $X=0.567 $Y=0.135 $X2=0.027 $Y2=0.135
cc_93 N_A_c_69_n N_Y_c_201_n 6.8292e-19 $X=0.297 $Y=0.135 $X2=0.351 $Y2=0.0675
cc_94 N_A_c_80_n N_Y_c_201_n 4.64672e-19 $X=0.298 $Y=0.189 $X2=0.351 $Y2=0.0675
cc_95 N_A_c_82_n N_Y_c_203_n 3.14976e-19 $X=0.527 $Y=0.189 $X2=0.351 $Y2=0.2025
cc_96 N_A_c_116_p N_Y_c_204_n 0.00126701f $X=0.567 $Y=0.1705 $X2=0 $Y2=0
cc_97 N_A_c_117_p N_Y_c_204_n 3.10247e-19 $X=0.567 $Y=0.189 $X2=0 $Y2=0
cc_98 N_A_M2_g N_Y_c_192_n 2.64369e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_99 N_A_c_82_n N_Y_c_207_n 4.77607e-19 $X=0.527 $Y=0.189 $X2=0 $Y2=0
cc_100 N_A_c_116_p Y 4.91816e-19 $X=0.567 $Y=0.1705 $X2=0.213 $Y2=0.036
cc_101 N_A_c_82_n Y 7.65288e-19 $X=0.527 $Y=0.189 $X2=0.213 $Y2=0.036
cc_102 N_A_c_122_p N_Y_c_210_n 4.01135e-19 $X=0.567 $Y=0.189 $X2=0.107 $Y2=0.036
cc_103 N_A_c_82_n N_Y_c_210_n 4.49897e-19 $X=0.527 $Y=0.189 $X2=0.107 $Y2=0.036
cc_104 N_A_c_82_n N_Y_c_212_n 9.16084e-19 $X=0.527 $Y=0.189 $X2=0.2025 $Y2=0.036
cc_105 N_A_M7_g N_Y_c_213_n 2.37298e-19 $X=0.567 $Y=0.0675 $X2=0.06 $Y2=0.136
cc_106 N_A_c_122_p N_Y_c_213_n 0.00520809f $X=0.567 $Y=0.189 $X2=0.06 $Y2=0.136
cc_107 N_A_c_82_n N_Y_c_200_n 2.40707e-19 $X=0.527 $Y=0.189 $X2=0.256 $Y2=0.076
cc_108 VSS N_A_c_122_p 3.03729e-19 $X=0.567 $Y=0.189 $X2=0.081 $Y2=0.0675
cc_109 VSS N_5_c_135_n 0.00251508f $X=0.16 $Y=0.0675 $X2=0.513 $Y2=0.2025
cc_110 VSS N_5_M4_g 3.77795e-19 $X=0.405 $Y=0.0675 $X2=0.213 $Y2=0.036
cc_111 VSS N_5_c_144_n 2.31252e-19 $X=0.405 $Y=0.135 $X2=0.213 $Y2=0.036
cc_112 VSS N_5_M5_g 2.86067e-19 $X=0.459 $Y=0.0675 $X2=0.078 $Y2=0.036
cc_113 N_5_c_133_n N_Y_M5_d 4.0989e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_114 N_5_c_133_n N_Y_c_217_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.135
cc_115 N_5_c_141_n N_Y_M10_d 3.26345e-19 $X=0.305 $Y=0.198 $X2=0.081 $Y2=0.2025
cc_116 N_5_c_155_n N_Y_c_201_n 3.69284e-19 $X=0.183 $Y=0.189 $X2=0.351
+ $Y2=0.0675
cc_117 N_5_c_177_p N_Y_c_201_n 3.59575e-19 $X=0.1835 $Y=0.225 $X2=0.351
+ $Y2=0.0675
cc_118 N_5_c_141_n N_Y_c_201_n 0.00279801f $X=0.305 $Y=0.198 $X2=0.351
+ $Y2=0.0675
cc_119 N_5_c_133_n N_Y_M13_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_120 N_5_c_133_n N_Y_c_203_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0.351
+ $Y2=0.2025
cc_121 N_5_c_181_p N_Y_c_203_n 0.00107102f $X=0.405 $Y=0.1665 $X2=0.351
+ $Y2=0.2025
cc_122 N_5_M4_g N_Y_c_192_n 2.34002e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_123 N_5_c_183_p N_Y_c_192_n 6.66585e-19 $X=0.174 $Y=0.234 $X2=0 $Y2=0
cc_124 N_5_c_141_n N_Y_c_192_n 0.0130846f $X=0.305 $Y=0.198 $X2=0 $Y2=0
cc_125 N_5_M5_g Y 3.07672e-19 $X=0.459 $Y=0.0675 $X2=0.213 $Y2=0.036
cc_126 N_5_c_144_n Y 0.0011985f $X=0.405 $Y=0.135 $X2=0.213 $Y2=0.036
cc_127 N_5_c_133_n N_Y_c_195_n 0.00230337f $X=0.459 $Y=0.135 $X2=0.078 $Y2=0.036
cc_128 N_5_c_144_n N_Y_c_195_n 0.0011985f $X=0.405 $Y=0.135 $X2=0.078 $Y2=0.036
cc_129 N_5_c_166_n N_Y_c_210_n 0.0011985f $X=0.405 $Y=0.189 $X2=0.107 $Y2=0.036
cc_130 N_5_c_133_n N_Y_c_200_n 4.91185e-19 $X=0.459 $Y=0.135 $X2=0.256 $Y2=0.076
cc_131 VSS N_5_c_142_n 4.42394e-19 $X=0.365 $Y=0.198 $X2=0.081 $Y2=0.0675
cc_132 VSS N_Y_c_217_n 0.0038608f $X=0.378 $Y=0.036 $X2=0.081 $Y2=0.135
cc_133 VSS N_Y_c_217_n 0.00387022f $X=0.486 $Y=0.036 $X2=0.081 $Y2=0.135
cc_134 VSS N_Y_c_217_n 0.00263673f $X=0.468 $Y=0.036 $X2=0.081 $Y2=0.135
cc_135 VSS N_Y_c_201_n 0.00169333f $X=0.27 $Y=0.036 $X2=0.351 $Y2=0.0675
cc_136 VSS N_Y_c_204_n 0.00107252f $X=0.594 $Y=0.036 $X2=0 $Y2=0
cc_137 VSS N_Y_c_198_n 6.21879e-19 $X=0.486 $Y=0.036 $X2=0.231 $Y2=0.076
cc_138 VSS N_Y_c_200_n 2.19246e-19 $X=0.378 $Y=0.036 $X2=0.256 $Y2=0.076
cc_139 VSS N_Y_c_200_n 0.00238589f $X=0.468 $Y=0.036 $X2=0.256 $Y2=0.076
cc_140 VSS N_Y_c_192_n 3.19084e-19 $X=0.414 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./XNOR2x1_ASAP7_75t_R.pex.sp.XNOR2X1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: XNOR2x2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:07:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "XNOR2x2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./XNOR2x2_ASAP7_75t_R.pex.sp.pex"
* File: XNOR2x2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:07:10 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_XNOR2X2_ASAP7_75T_R%3 2 5 7 9 10 13 14 24 27 30 31 34 35 36 37 42 44
+ 45 VSS
c36 49 VSS 0.00179571f $X=0.311 $Y=0.072
c37 45 VSS 7.99121e-21 $X=0.36 $Y=0.072
c38 44 VSS 0.00213751f $X=0.342 $Y=0.072
c39 42 VSS 6.88106e-19 $X=0.378 $Y=0.072
c40 37 VSS 7.70271e-19 $X=0.311 $Y=0.12
c41 36 VSS 7.6369e-19 $X=0.311 $Y=0.107
c42 35 VSS 0.014335f $X=0.311 $Y=0.18
c43 34 VSS 0.00135266f $X=0.311 $Y=0.18
c44 31 VSS 0.00208239f $X=0.279 $Y=0.072
c45 30 VSS 8.46035e-21 $X=0.144 $Y=0.072
c46 29 VSS 0.00220046f $X=0.126 $Y=0.072
c47 28 VSS 1.81812e-19 $X=0.099 $Y=0.072
c48 27 VSS 4.67334e-20 $X=0.09 $Y=0.072
c49 26 VSS 3.79585e-19 $X=0.302 $Y=0.072
c50 24 VSS 1.15487e-19 $X=0.081 $Y=0.1275
c51 23 VSS 0.00161525f $X=0.081 $Y=0.12
c52 21 VSS 2.98192e-19 $X=0.081 $Y=0.135
c53 14 VSS 4.79903e-19 $X=0.341 $Y=0.2025
c54 13 VSS 0.024763f $X=0.378 $Y=0.054
c55 9 VSS 5.52978e-19 $X=0.395 $Y=0.054
c56 5 VSS 0.00172734f $X=0.081 $Y=0.135
c57 2 VSS 0.0664387f $X=0.081 $Y=0.0675
r58 44 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.072 $X2=0.36 $Y2=0.072
r59 42 45 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.072 $X2=0.36 $Y2=0.072
r60 40 49 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.32
+ $Y=0.072 $X2=0.311 $Y2=0.072
r61 40 44 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.32
+ $Y=0.072 $X2=0.342 $Y2=0.072
r62 36 37 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.107 $X2=0.311 $Y2=0.12
r63 34 37 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.18 $X2=0.311 $Y2=0.12
r64 34 35 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.311 $Y=0.18 $X2=0.311
+ $Y2=0.18
r65 32 49 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.081 $X2=0.311 $Y2=0.072
r66 32 36 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.311
+ $Y=0.081 $X2=0.311 $Y2=0.107
r67 30 31 9.16667 $w=1.8e-08 $l=1.35e-07 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.072 $X2=0.279 $Y2=0.072
r68 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.072 $X2=0.144 $Y2=0.072
r69 28 29 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.099
+ $Y=0.072 $X2=0.126 $Y2=0.072
r70 27 28 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.099 $Y2=0.072
r71 26 49 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.302
+ $Y=0.072 $X2=0.311 $Y2=0.072
r72 26 31 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.302
+ $Y=0.072 $X2=0.279 $Y2=0.072
r73 23 24 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.12 $X2=0.081 $Y2=0.1275
r74 21 24 0.509259 $w=1.8e-08 $l=7.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1275
r75 19 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.081 $X2=0.09 $Y2=0.072
r76 19 23 2.64815 $w=1.8e-08 $l=3.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.081 $X2=0.081 $Y2=0.12
r77 17 35 9.51166 $w=4.9e-08 $l=2.25e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.3115 $Y=0.2025 $X2=0.3115 $Y2=0.18
r78 14 17 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.341 $Y=0.2025 $X2=0.326 $Y2=0.2025
r79 13 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.072 $X2=0.378
+ $Y2=0.072
r80 10 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.054 $X2=0.378 $Y2=0.054
r81 9 13 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.054 $X2=0.378 $Y2=0.054
r82 5 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r83 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r84 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_XNOR2X2_ASAP7_75T_R%A 2 5 7 10 13 15 19 23 24 25 26 30 32 33 34 35 36
+ 37 43 44 45 47 49 54 VSS
c47 55 VSS 4.47597e-19 $X=0.422 $Y=0.135
c48 54 VSS 3.7015e-19 $X=0.431 $Y=0.135
c49 49 VSS 3.89437e-19 $X=0.405 $Y=0.135
c50 47 VSS 0.00109749f $X=0.431 $Y=0.207
c51 45 VSS 2.19188e-19 $X=0.431 $Y=0.1595
c52 44 VSS 1.73467e-19 $X=0.431 $Y=0.151
c53 43 VSS 0.00227175f $X=0.435 $Y=0.168
c54 41 VSS 9.62667e-19 $X=0.431 $Y=0.225
c55 39 VSS 0.00128265f $X=0.4065 $Y=0.234
c56 38 VSS 0.00120569f $X=0.391 $Y=0.234
c57 37 VSS 0.00322944f $X=0.38 $Y=0.234
c58 36 VSS 0.00199133f $X=0.342 $Y=0.234
c59 35 VSS 0.00134741f $X=0.32 $Y=0.234
c60 34 VSS 0.00205247f $X=0.302 $Y=0.234
c61 33 VSS 0.00231441f $X=0.279 $Y=0.234
c62 32 VSS 0.00518267f $X=0.422 $Y=0.234
c63 31 VSS 3.48791e-20 $X=0.27 $Y=0.216
c64 30 VSS 9.67341e-21 $X=0.27 $Y=0.207
c65 29 VSS 3.29414e-20 $X=0.27 $Y=0.225
c66 27 VSS 8.52667e-19 $X=0.2455 $Y=0.192
c67 26 VSS 0.00320415f $X=0.23 $Y=0.192
c68 25 VSS 5.19699e-20 $X=0.144 $Y=0.192
c69 24 VSS 9.56956e-19 $X=0.261 $Y=0.192
c70 23 VSS 3.43945e-19 $X=0.135 $Y=0.166
c71 19 VSS 2.89281e-19 $X=0.135 $Y=0.135
c72 17 VSS 7.57456e-19 $X=0.135 $Y=0.183
c73 13 VSS 0.00159436f $X=0.405 $Y=0.135
c74 10 VSS 0.0595161f $X=0.405 $Y=0.054
c75 5 VSS 0.0014528f $X=0.135 $Y=0.135
c76 2 VSS 0.0618866f $X=0.135 $Y=0.0675
r77 55 56 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.422
+ $Y=0.135 $X2=0.423 $Y2=0.135
r78 54 56 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.135 $X2=0.423 $Y2=0.135
r79 49 55 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.422 $Y2=0.135
r80 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.189 $X2=0.431 $Y2=0.207
r81 44 45 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.151 $X2=0.431 $Y2=0.1595
r82 43 46 1.42593 $w=1.8e-08 $l=2.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.168 $X2=0.431 $Y2=0.189
r83 43 45 0.57716 $w=1.8e-08 $l=8.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.168 $X2=0.431 $Y2=0.1595
r84 41 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.225 $X2=0.431 $Y2=0.207
r85 40 54 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.144 $X2=0.431 $Y2=0.135
r86 40 44 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.431
+ $Y=0.144 $X2=0.431 $Y2=0.151
r87 38 39 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.391
+ $Y=0.234 $X2=0.4065 $Y2=0.234
r88 37 38 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.38
+ $Y=0.234 $X2=0.391 $Y2=0.234
r89 36 37 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.38 $Y2=0.234
r90 35 36 1.49383 $w=1.8e-08 $l=2.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.32
+ $Y=0.234 $X2=0.342 $Y2=0.234
r91 34 35 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.302
+ $Y=0.234 $X2=0.32 $Y2=0.234
r92 33 34 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.279
+ $Y=0.234 $X2=0.302 $Y2=0.234
r93 32 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.422 $Y=0.234 $X2=0.431 $Y2=0.225
r94 32 39 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.422
+ $Y=0.234 $X2=0.4065 $Y2=0.234
r95 30 31 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.207 $X2=0.27 $Y2=0.216
r96 29 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.27 $Y=0.225 $X2=0.279 $Y2=0.234
r97 29 31 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.225 $X2=0.27 $Y2=0.216
r98 28 30 0.407407 $w=1.8e-08 $l=6e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.201 $X2=0.27 $Y2=0.207
r99 26 27 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.192 $X2=0.2455 $Y2=0.192
r100 25 26 5.83951 $w=1.8e-08 $l=8.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.192 $X2=0.23 $Y2=0.192
r101 24 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.261 $Y=0.192 $X2=0.27 $Y2=0.201
r102 24 27 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.192 $X2=0.2455 $Y2=0.192
r103 22 23 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.149 $X2=0.135 $Y2=0.166
r104 19 22 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.149
r105 17 25 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.135 $Y=0.183 $X2=0.144 $Y2=0.192
r106 17 23 1.15432 $w=1.8e-08 $l=1.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.183 $X2=0.135 $Y2=0.166
r107 13 49 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r108 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r109 10 13 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.054 $X2=0.405 $Y2=0.135
r110 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r111 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r112 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_XNOR2X2_ASAP7_75T_R%B 2 7 10 13 15 19 VSS
c33 19 VSS 0.00174301f $X=0.35 $Y=0.135
c34 13 VSS 0.0161697f $X=0.351 $Y=0.135
c35 10 VSS 0.0634112f $X=0.351 $Y=0.054
c36 2 VSS 0.0655384f $X=0.189 $Y=0.0675
r37 13 19 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r38 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r39 10 13 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.054 $X2=0.351 $Y2=0.135
r40 5 13 202.5 $w=1.6e-08 $l=1.62e-07 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.351 $Y2=0.135
r41 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r42 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_XNOR2X2_ASAP7_75T_R%6 2 7 10 13 15 17 22 25 27 30 35 36 38 42 45 48
+ 49 52 53 55 58 60 61 66 VSS
c46 69 VSS 9.17717e-19 $X=0.045 $Y=0.234
c47 68 VSS 0.00328948f $X=0.036 $Y=0.234
c48 66 VSS 0.0023031f $X=0.054 $Y=0.234
c49 61 VSS 6.14257e-19 $X=0.486 $Y=0.126
c50 60 VSS 7.00628e-19 $X=0.486 $Y=0.107
c51 58 VSS 6.14726e-19 $X=0.486 $Y=0.135
c52 55 VSS 5.06567e-20 $X=0.4745 $Y=0.072
c53 54 VSS 0.00185179f $X=0.472 $Y=0.072
c54 53 VSS 0.00120419f $X=0.441 $Y=0.072
c55 52 VSS 1.3551e-19 $X=0.477 $Y=0.072
c56 51 VSS 6.41935e-19 $X=0.432 $Y=0.063
c57 49 VSS 0.00134702f $X=0.4075 $Y=0.036
c58 48 VSS 0.0323459f $X=0.392 $Y=0.036
c59 47 VSS 8.76814e-19 $X=0.072 $Y=0.036
c60 46 VSS 0.00270525f $X=0.063 $Y=0.036
c61 45 VSS 0.00505797f $X=0.216 $Y=0.036
c62 42 VSS 0.00677526f $X=0.054 $Y=0.036
c63 39 VSS 0.00341041f $X=0.036 $Y=0.036
c64 38 VSS 0.00511688f $X=0.423 $Y=0.036
c65 37 VSS 3.97344e-19 $X=0.027 $Y=0.213
c66 36 VSS 0.0023522f $X=0.027 $Y=0.201
c67 35 VSS 0.00368965f $X=0.027 $Y=0.149
c68 34 VSS 5.7946e-19 $X=0.027 $Y=0.063
c69 33 VSS 3.80788e-19 $X=0.027 $Y=0.225
c70 30 VSS 0.002959f $X=0.056 $Y=0.2025
c71 27 VSS 3.25039e-19 $X=0.071 $Y=0.2025
c72 25 VSS 4.39464e-19 $X=0.214 $Y=0.0675
c73 17 VSS 2.69461e-19 $X=0.071 $Y=0.0675
c74 13 VSS 0.00427632f $X=0.513 $Y=0.135
c75 10 VSS 0.0639847f $X=0.513 $Y=0.0675
c76 2 VSS 0.0613093f $X=0.459 $Y=0.0675
r77 68 69 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.045 $Y2=0.234
r78 66 69 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.045 $Y2=0.234
r79 63 68 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.036 $Y2=0.234
r80 60 61 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.107 $X2=0.486 $Y2=0.126
r81 58 61 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.135 $X2=0.486 $Y2=0.126
r82 58 59 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.486 $Y=0.135 $X2=0.486
+ $Y2=0.135
r83 56 60 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.081 $X2=0.486 $Y2=0.107
r84 54 55 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.472
+ $Y=0.072 $X2=0.4745 $Y2=0.072
r85 53 54 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.441
+ $Y=0.072 $X2=0.472 $Y2=0.072
r86 52 56 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.477 $Y=0.072 $X2=0.486 $Y2=0.081
r87 52 55 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.477
+ $Y=0.072 $X2=0.4745 $Y2=0.072
r88 51 53 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.432 $Y=0.063 $X2=0.441 $Y2=0.072
r89 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.045 $X2=0.432 $Y2=0.063
r90 48 49 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.392
+ $Y=0.036 $X2=0.4075 $Y2=0.036
r91 46 47 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.036 $X2=0.072 $Y2=0.036
r92 44 48 11.9506 $w=1.8e-08 $l=1.76e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.392 $Y2=0.036
r93 44 47 9.77778 $w=1.8e-08 $l=1.44e-07 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.036 $X2=0.072 $Y2=0.036
r94 44 45 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.036 $X2=0.216
+ $Y2=0.036
r95 41 46 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.063 $Y2=0.036
r96 41 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r97 39 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.054 $Y2=0.036
r98 38 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.423 $Y=0.036 $X2=0.432 $Y2=0.045
r99 38 49 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.423
+ $Y=0.036 $X2=0.4075 $Y2=0.036
r100 36 37 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.201 $X2=0.027 $Y2=0.213
r101 35 36 3.53086 $w=1.8e-08 $l=5.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.149 $X2=0.027 $Y2=0.201
r102 34 35 5.83951 $w=1.8e-08 $l=8.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.063 $X2=0.027 $Y2=0.149
r103 33 63 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.234
r104 33 37 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.213
r105 32 39 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.045 $X2=0.036 $Y2=0.036
r106 32 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.063
r107 30 66 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234
+ $X2=0.054 $Y2=0.234
r108 27 30 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2025 $X2=0.056 $Y2=0.2025
r109 25 45 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.216 $Y=0.0675 $X2=0.216 $Y2=0.036
r110 22 25 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.214 $Y2=0.0675
r111 20 42 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08
+ $X=0.054 $Y=0.0675 $X2=0.054 $Y2=0.036
r112 17 20 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0675 $X2=0.056 $Y2=0.0675
r113 13 59 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.513
+ $Y=0.135 $X2=0.486 $Y2=0.135
r114 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.135 $X2=0.513 $Y2=0.2025
r115 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.513 $Y=0.0675 $X2=0.513 $Y2=0.135
r116 5 59 24.5455 $w=2.2e-08 $l=2.7e-08 $layer=LIG $thickness=5e-08 $X=0.459
+ $Y=0.135 $X2=0.486 $Y2=0.135
r117 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r118 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
.ends

.subckt PM_XNOR2X2_ASAP7_75T_R%Y 1 2 6 7 10 14 16 17 20 26 28 30 32 34 VSS
c21 34 VSS 0.00219831f $X=0.567 $Y=0.188
c22 32 VSS 0.00213894f $X=0.567 $Y=0.10525
c23 31 VSS 8.85605e-19 $X=0.567 $Y=0.063
c24 30 VSS 0.00213572f $X=0.567 $Y=0.1475
c25 28 VSS 0.00190935f $X=0.567 $Y=0.225
c26 26 VSS 0.00278214f $X=0.5265 $Y=0.234
c27 25 VSS 0.00107061f $X=0.495 $Y=0.234
c28 20 VSS 0.00154248f $X=0.486 $Y=0.234
c29 18 VSS 0.00875248f $X=0.558 $Y=0.234
c30 17 VSS 0.00278214f $X=0.5265 $Y=0.036
c31 16 VSS 0.00252716f $X=0.495 $Y=0.036
c32 14 VSS 0.0108098f $X=0.486 $Y=0.036
c33 11 VSS 0.00875248f $X=0.558 $Y=0.036
c34 10 VSS 0.00915654f $X=0.486 $Y=0.2025
c35 6 VSS 5.72268e-19 $X=0.503 $Y=0.2025
c36 1 VSS 6.04166e-19 $X=0.503 $Y=0.0675
r37 33 34 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.151 $X2=0.567 $Y2=0.188
r38 31 32 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.063 $X2=0.567 $Y2=0.10525
r39 30 33 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.1475 $X2=0.567 $Y2=0.151
r40 30 32 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.1475 $X2=0.567 $Y2=0.10525
r41 28 34 2.51235 $w=1.8e-08 $l=3.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.225 $X2=0.567 $Y2=0.188
r42 27 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.567
+ $Y=0.045 $X2=0.567 $Y2=0.063
r43 25 26 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.234 $X2=0.5265 $Y2=0.234
r44 20 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.234 $X2=0.495 $Y2=0.234
r45 18 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.234 $X2=0.567 $Y2=0.225
r46 18 26 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.5265 $Y2=0.234
r47 16 17 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.495
+ $Y=0.036 $X2=0.5265 $Y2=0.036
r48 13 16 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.495 $Y2=0.036
r49 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036 $X2=0.486
+ $Y2=0.036
r50 11 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.558 $Y=0.036 $X2=0.567 $Y2=0.045
r51 11 17 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.5265 $Y2=0.036
r52 10 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r53 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.486 $Y2=0.2025
r54 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.2025 $X2=0.486 $Y2=0.2025
r55 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0675 $X2=0.486 $Y2=0.036
r56 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.0675 $X2=0.486 $Y2=0.0675
r57 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.503
+ $Y=0.0675 $X2=0.486 $Y2=0.0675
.ends

.subckt PM_XNOR2X2_ASAP7_75T_R%10 1 2 VSS
c0 1 VSS 0.00243838f $X=0.395 $Y=0.2025
r1 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.2025 $X2=0.361 $Y2=0.2025
.ends


* END of "./XNOR2x2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt XNOR2x2_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 VSS N_3_M0_g N_6_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 noxref_9 N_A_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_6_M2_d N_B_M2_g noxref_9 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_3_M3_d N_B_M3_g VSS VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.341 $Y=0.027
M4 VSS N_A_M4_g N_3_M4_s VSS NMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.395 $Y=0.027
M5 N_Y_M5_d N_6_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M6 N_Y_M6_d N_6_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503 $Y=0.027
M7 noxref_7 N_3_M7_g N_6_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M8 VDD N_A_M8_g noxref_7 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M9 noxref_7 N_B_M9_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.162
M10 N_10_M10_d N_B_M10_g N_3_M10_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.341 $Y=0.162
M11 VDD N_A_M11_g N_10_M11_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M12 N_Y_M12_d N_6_M12_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
M13 N_Y_M13_d N_6_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.162
*
* 
* .include "XNOR2x2_ASAP7_75t_R.pex.sp.XNOR2X2_ASAP7_75T_R.pxi"
* BEGIN of "./XNOR2x2_ASAP7_75t_R.pex.sp.XNOR2X2_ASAP7_75T_R.pxi"
* File: XNOR2x2_ASAP7_75t_R.pex.sp.XNOR2X2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:07:10 2017
* 
x_PM_XNOR2X2_ASAP7_75T_R%3 N_3_M0_g N_3_c_3_p N_3_M7_g N_3_M4_s N_3_M3_d
+ N_3_c_32_p N_3_M10_s N_3_c_4_p N_3_c_27_p N_3_c_2_p N_3_c_9_p N_3_c_6_p
+ N_3_c_8_p N_3_c_30_p N_3_c_23_p N_3_c_24_p N_3_c_20_p N_3_c_16_p VSS
+ PM_XNOR2X2_ASAP7_75T_R%3
x_PM_XNOR2X2_ASAP7_75T_R%A N_A_M1_g N_A_c_39_n N_A_M8_g N_A_M4_g N_A_c_55_p
+ N_A_M11_g N_A_c_40_n N_A_c_67_p N_A_c_43_n N_A_c_80_p N_A_c_45_n N_A_c_76_p
+ N_A_c_81_p N_A_c_78_p N_A_c_46_n N_A_c_47_n N_A_c_49_n N_A_c_53_p A N_A_c_60_p
+ N_A_c_61_p N_A_c_62_p N_A_c_63_p N_A_c_72_p VSS PM_XNOR2X2_ASAP7_75T_R%A
x_PM_XNOR2X2_ASAP7_75T_R%B N_B_M2_g N_B_M9_g N_B_M3_g N_B_c_87_n N_B_M10_g B VSS
+ PM_XNOR2X2_ASAP7_75T_R%B
x_PM_XNOR2X2_ASAP7_75T_R%6 N_6_M5_g N_6_M12_g N_6_M6_g N_6_c_128_n N_6_M13_g
+ N_6_M0_s N_6_M2_d N_6_c_117_n N_6_M7_s N_6_c_141_p N_6_c_118_n N_6_c_129_n
+ N_6_c_130_n N_6_c_119_n N_6_c_120_n N_6_c_122_n N_6_c_132_n N_6_c_148_p
+ N_6_c_125_n N_6_c_149_p N_6_c_135_n N_6_c_150_p N_6_c_140_n N_6_c_143_p VSS
+ PM_XNOR2X2_ASAP7_75T_R%6
x_PM_XNOR2X2_ASAP7_75T_R%Y N_Y_M6_d N_Y_M5_d N_Y_M13_d N_Y_M12_d N_Y_c_168_n
+ N_Y_c_169_n N_Y_c_174_n N_Y_c_176_n N_Y_c_163_n N_Y_c_179_n N_Y_c_164_n Y
+ N_Y_c_183_n N_Y_c_165_n VSS PM_XNOR2X2_ASAP7_75T_R%Y
x_PM_XNOR2X2_ASAP7_75T_R%10 N_10_M11_s N_10_M10_d VSS PM_XNOR2X2_ASAP7_75T_R%10
cc_1 N_3_M0_g N_A_M1_g 0.00323392f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_3_c_2_p N_A_M1_g 2.98356e-19 $X=0.144 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_3 N_3_c_3_p N_A_c_39_n 9.46013e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_4 N_3_c_4_p N_A_c_40_n 0.00118961f $X=0.081 $Y=0.1275 $X2=0.135 $Y2=0.135
cc_5 N_3_c_2_p N_A_c_40_n 7.96353e-19 $X=0.144 $Y=0.072 $X2=0.135 $Y2=0.135
cc_6 N_3_c_6_p N_A_c_40_n 2.88965e-19 $X=0.311 $Y=0.18 $X2=0.135 $Y2=0.135
cc_7 N_3_c_6_p N_A_c_43_n 7.35029e-19 $X=0.311 $Y=0.18 $X2=0.261 $Y2=0.192
cc_8 N_3_c_8_p N_A_c_43_n 4.85208e-19 $X=0.311 $Y=0.18 $X2=0.261 $Y2=0.192
cc_9 N_3_c_9_p N_A_c_45_n 0.00164688f $X=0.279 $Y=0.072 $X2=0.23 $Y2=0.192
cc_10 N_3_c_8_p N_A_c_46_n 0.00117999f $X=0.311 $Y=0.18 $X2=0.302 $Y2=0.234
cc_11 N_3_c_6_p N_A_c_47_n 8.67348e-19 $X=0.311 $Y=0.18 $X2=0.32 $Y2=0.234
cc_12 N_3_c_8_p N_A_c_47_n 0.0012608f $X=0.311 $Y=0.18 $X2=0.32 $Y2=0.234
cc_13 N_3_c_8_p N_A_c_49_n 0.00195414f $X=0.311 $Y=0.18 $X2=0.342 $Y2=0.234
cc_14 N_3_M0_g N_B_M2_g 2.34385e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_15 N_3_c_9_p N_B_M2_g 4.07897e-19 $X=0.279 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_16 N_3_c_16_p N_B_M3_g 2.81878e-19 $X=0.36 $Y=0.072 $X2=0.405 $Y2=0.054
cc_17 N_3_c_9_p N_B_c_87_n 0.00128776f $X=0.279 $Y=0.072 $X2=0.405 $Y2=0.135
cc_18 N_3_c_6_p N_B_c_87_n 0.00237361f $X=0.311 $Y=0.18 $X2=0.405 $Y2=0.135
cc_19 N_3_c_8_p N_B_c_87_n 0.00268514f $X=0.311 $Y=0.18 $X2=0.405 $Y2=0.135
cc_20 N_3_c_20_p N_B_c_87_n 5.46915e-19 $X=0.342 $Y=0.072 $X2=0.405 $Y2=0.135
cc_21 N_3_c_6_p B 0.00402878f $X=0.311 $Y=0.18 $X2=0.135 $Y2=0.135
cc_22 N_3_c_8_p B 0.00117504f $X=0.311 $Y=0.18 $X2=0.135 $Y2=0.135
cc_23 N_3_c_23_p B 0.00201439f $X=0.311 $Y=0.12 $X2=0.135 $Y2=0.135
cc_24 N_3_c_24_p B 2.72962e-19 $X=0.378 $Y=0.072 $X2=0.135 $Y2=0.135
cc_25 N_3_c_16_p B 0.00119465f $X=0.36 $Y=0.072 $X2=0.135 $Y2=0.135
cc_26 N_3_c_9_p N_6_c_117_n 3.28501e-19 $X=0.279 $Y=0.072 $X2=0.144 $Y2=0.192
cc_27 N_3_c_27_p N_6_c_118_n 0.00345167f $X=0.09 $Y=0.072 $X2=0.32 $Y2=0.234
cc_28 N_3_c_27_p N_6_c_119_n 0.00136685f $X=0.09 $Y=0.072 $X2=0.431 $Y2=0.168
cc_29 N_3_c_9_p N_6_c_120_n 0.0028283f $X=0.279 $Y=0.072 $X2=0.431 $Y2=0.1595
cc_30 N_3_c_30_p N_6_c_120_n 6.58653e-19 $X=0.311 $Y=0.107 $X2=0.431 $Y2=0.1595
cc_31 N_3_M0_g N_6_c_122_n 2.34993e-19 $X=0.081 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_32 N_3_c_32_p N_6_c_122_n 0.00255062f $X=0.378 $Y=0.054 $X2=0.405 $Y2=0.135
cc_33 N_3_c_27_p N_6_c_122_n 0.0270759f $X=0.09 $Y=0.072 $X2=0.405 $Y2=0.135
cc_34 N_3_c_24_p N_6_c_125_n 9.4025e-19 $X=0.378 $Y=0.072 $X2=0 $Y2=0
cc_35 VSS N_3_c_8_p 0.00216384f $X=0.311 $Y=0.18 $X2=0.405 $Y2=0.054
cc_36 VSS N_3_c_9_p 5.0983e-19 $X=0.279 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_37 N_A_M1_g N_B_M2_g 0.00323392f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_38 N_A_c_45_n N_B_M2_g 4.15003e-19 $X=0.23 $Y=0.192 $X2=0.081 $Y2=0.0675
cc_39 N_A_M4_g N_B_M3_g 0.00344695f $X=0.405 $Y=0.054 $X2=0.361 $Y2=0.054
cc_40 N_A_c_53_p N_B_M3_g 2.38942e-19 $X=0.38 $Y=0.234 $X2=0.361 $Y2=0.054
cc_41 N_A_c_39_n N_B_c_87_n 0.00106649f $X=0.135 $Y=0.135 $X2=0.378 $Y2=0.054
cc_42 N_A_c_55_p N_B_c_87_n 8.77417e-19 $X=0.405 $Y=0.135 $X2=0.378 $Y2=0.054
cc_43 N_A_c_45_n N_B_c_87_n 0.00133346f $X=0.23 $Y=0.192 $X2=0.378 $Y2=0.054
cc_44 N_A_c_49_n N_B_c_87_n 2.02767e-19 $X=0.342 $Y=0.234 $X2=0.378 $Y2=0.054
cc_45 N_A_c_43_n B 3.36274e-19 $X=0.261 $Y=0.192 $X2=0.081 $Y2=0.081
cc_46 N_A_c_53_p B 0.00408388f $X=0.38 $Y=0.234 $X2=0.081 $Y2=0.081
cc_47 N_A_c_60_p B 5.60314e-19 $X=0.431 $Y=0.151 $X2=0.081 $Y2=0.081
cc_48 N_A_c_61_p B 5.60314e-19 $X=0.431 $Y=0.1595 $X2=0.081 $Y2=0.081
cc_49 N_A_c_62_p B 6.37279e-19 $X=0.431 $Y=0.207 $X2=0.081 $Y2=0.081
cc_50 N_A_c_63_p B 8.81039e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.081
cc_51 N_A_M4_g N_6_M5_g 0.00284417f $X=0.405 $Y=0.054 $X2=0.081 $Y2=0.0675
cc_52 N_A_M4_g N_6_M6_g 2.31381e-19 $X=0.405 $Y=0.054 $X2=0.361 $Y2=0.054
cc_53 N_A_c_55_p N_6_c_128_n 0.00102897f $X=0.405 $Y=0.135 $X2=0.378 $Y2=0.054
cc_54 N_A_c_67_p N_6_c_129_n 5.60011e-19 $X=0.135 $Y=0.166 $X2=0.311 $Y2=0.107
cc_55 N_A_c_63_p N_6_c_130_n 3.07195e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_56 N_A_M1_g N_6_c_122_n 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_57 N_A_M4_g N_6_c_132_n 2.67908e-19 $X=0.405 $Y=0.054 $X2=0.311 $Y2=0.072
cc_58 N_A_c_63_p N_6_c_132_n 3.07195e-19 $X=0.405 $Y=0.135 $X2=0.311 $Y2=0.072
cc_59 N_A_c_72_p N_6_c_125_n 7.6078e-19 $X=0.431 $Y=0.135 $X2=0.3115 $Y2=0.18
cc_60 N_A_c_72_p N_6_c_135_n 0.00112769f $X=0.431 $Y=0.135 $X2=0 $Y2=0
cc_61 VSS N_A_c_67_p 0.00136835f $X=0.135 $Y=0.166 $X2=0.081 $Y2=0.135
cc_62 VSS N_A_c_45_n 0.00256063f $X=0.23 $Y=0.192 $X2=0.395 $Y2=0.054
cc_63 VSS N_A_c_76_p 8.24756e-19 $X=0.27 $Y=0.207 $X2=0.395 $Y2=0.054
cc_64 VSS N_A_c_45_n 0.00337967f $X=0.23 $Y=0.192 $X2=0 $Y2=0
cc_65 VSS N_A_c_78_p 0.00123078f $X=0.279 $Y=0.234 $X2=0 $Y2=0
cc_66 VSS N_A_M1_g 2.60742e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.081
cc_67 VSS N_A_c_80_p 0.00337967f $X=0.144 $Y=0.192 $X2=0.081 $Y2=0.081
cc_68 N_A_c_81_p N_Y_c_163_n 0.00108419f $X=0.422 $Y=0.234 $X2=0.081 $Y2=0.135
cc_69 N_A_c_61_p N_Y_c_164_n 2.15083e-19 $X=0.431 $Y=0.1595 $X2=0.099 $Y2=0.072
cc_70 N_A_c_72_p N_Y_c_165_n 2.15083e-19 $X=0.431 $Y=0.135 $X2=0.311 $Y2=0.18
cc_71 N_B_M3_g N_6_M5_g 2.31381e-19 $X=0.351 $Y=0.054 $X2=0.081 $Y2=0.0675
cc_72 N_B_c_87_n N_6_c_120_n 6.8292e-19 $X=0.351 $Y=0.135 $X2=0.36 $Y2=0.072
cc_73 N_B_M2_g N_6_c_122_n 2.65491e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_74 N_B_M3_g N_6_c_122_n 2.38942e-19 $X=0.351 $Y=0.054 $X2=0 $Y2=0
cc_75 B N_6_c_140_n 3.03334e-19 $X=0.35 $Y=0.135 $X2=0 $Y2=0
cc_76 VSS N_B_c_87_n 6.8292e-19 $X=0.351 $Y=0.135 $X2=0.395 $Y2=0.054
cc_77 VSS N_B_M2_g 2.90722e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_78 VSS N_6_c_141_p 0.00391186f $X=0.056 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_79 VSS N_6_c_120_n 0.00169333f $X=0.216 $Y=0.036 $X2=0.395 $Y2=0.054
cc_80 VSS N_6_c_143_p 6.5272e-19 $X=0.054 $Y=0.234 $X2=0 $Y2=0
cc_81 N_6_c_128_n N_Y_M6_d 3.80455e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_82 N_6_c_128_n N_Y_M13_d 3.80663e-19 $X=0.513 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_83 N_6_c_128_n N_Y_c_168_n 5.9618e-19 $X=0.513 $Y=0.135 $X2=0.361 $Y2=0.054
cc_84 N_6_c_128_n N_Y_c_169_n 8.00061e-19 $X=0.513 $Y=0.135 $X2=0.341 $Y2=0.2025
cc_85 N_6_c_148_p N_Y_c_169_n 0.00130196f $X=0.477 $Y=0.072 $X2=0.341 $Y2=0.2025
cc_86 N_6_c_149_p N_Y_c_169_n 3.88373e-19 $X=0.4745 $Y=0.072 $X2=0.341
+ $Y2=0.2025
cc_87 N_6_c_150_p N_Y_c_169_n 0.00147706f $X=0.486 $Y=0.107 $X2=0.341 $Y2=0.2025
cc_88 N_6_c_140_n N_Y_c_169_n 5.6276e-19 $X=0.486 $Y=0.126 $X2=0.341 $Y2=0.2025
cc_89 N_6_c_130_n N_Y_c_174_n 9.63474e-19 $X=0.423 $Y=0.036 $X2=0 $Y2=0
cc_90 N_6_c_149_p N_Y_c_174_n 0.00176732f $X=0.4745 $Y=0.072 $X2=0 $Y2=0
cc_91 N_6_M6_g N_Y_c_176_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.326 $Y2=0.2025
cc_92 N_6_c_128_n N_Y_c_176_n 3.25494e-19 $X=0.513 $Y=0.135 $X2=0.326 $Y2=0.2025
cc_93 N_6_c_135_n N_Y_c_163_n 3.89018e-19 $X=0.486 $Y=0.135 $X2=0.081 $Y2=0.135
cc_94 N_6_M6_g N_Y_c_179_n 4.59284e-19 $X=0.513 $Y=0.0675 $X2=0.302 $Y2=0.072
cc_95 N_6_c_128_n N_Y_c_179_n 3.25494e-19 $X=0.513 $Y=0.135 $X2=0.302 $Y2=0.072
cc_96 N_6_c_128_n Y 3.82643e-19 $X=0.513 $Y=0.135 $X2=0.144 $Y2=0.072
cc_97 N_6_c_140_n Y 9.11642e-19 $X=0.486 $Y=0.126 $X2=0.144 $Y2=0.072
cc_98 N_6_c_148_p N_Y_c_183_n 9.11642e-19 $X=0.477 $Y=0.072 $X2=0.311 $Y2=0.081
cc_99 VSS N_6_c_122_n 3.33359e-19 $X=0.392 $Y=0.036 $X2=0.081 $Y2=0.0675

* END of "./XNOR2x2_ASAP7_75t_R.pex.sp.XNOR2X2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: XNOR2xp5_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:07:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "XNOR2xp5_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./XNOR2xp5_ASAP7_75t_R.pex.sp.pex"
* File: XNOR2xp5_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:07:33 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_XNOR2XP5_ASAP7_75T_R%A 2 5 7 10 13 15 18 20 26 31 32 33 36 41 42 43
+ 44 45 48 51 53 VSS
c38 53 VSS 0.00754613f $X=0.018 $Y=0.135
c39 51 VSS 4.24224e-19 $X=0.351 $Y=0.128
c40 50 VSS 0.00154135f $X=0.351 $Y=0.121
c41 48 VSS 5.24005e-20 $X=0.351 $Y=0.135
c42 45 VSS 1.78615e-19 $X=0.3015 $Y=0.072
c43 44 VSS 0.0019627f $X=0.261 $Y=0.072
c44 43 VSS 1.80165e-19 $X=0.225 $Y=0.072
c45 42 VSS 0.00284881f $X=0.342 $Y=0.072
c46 41 VSS 6.38596e-24 $X=0.216 $Y=0.063
c47 36 VSS 0.00203697f $X=0.06 $Y=0.136
c48 33 VSS 0.00133719f $X=0.18 $Y=0.036
c49 32 VSS 0.00181942f $X=0.162 $Y=0.036
c50 31 VSS 0.00321912f $X=0.144 $Y=0.036
c51 30 VSS 0.00131186f $X=0.106 $Y=0.036
c52 29 VSS 0.00145201f $X=0.094 $Y=0.036
c53 28 VSS 0.00785083f $X=0.078 $Y=0.036
c54 27 VSS 0.0032309f $X=0.027 $Y=0.036
c55 26 VSS 0.00472496f $X=0.207 $Y=0.036
c56 20 VSS 8.69458e-19 $X=0.018 $Y=0.081
c57 19 VSS 6.58554e-19 $X=0.018 $Y=0.063
c58 18 VSS 0.00218042f $X=0.018 $Y=0.126
c59 13 VSS 0.00145322f $X=0.351 $Y=0.135
c60 10 VSS 0.0618866f $X=0.351 $Y=0.0675
c61 5 VSS 0.00580911f $X=0.081 $Y=0.135
c62 2 VSS 0.0638905f $X=0.081 $Y=0.0675
r63 50 51 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.121 $X2=0.351 $Y2=0.128
r64 48 51 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.128
r65 46 50 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.121
r66 44 45 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.261
+ $Y=0.072 $X2=0.3015 $Y2=0.072
r67 43 44 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.072 $X2=0.261 $Y2=0.072
r68 42 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.072 $X2=0.351 $Y2=0.081
r69 42 45 2.75 $w=1.8e-08 $l=4.05e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.072 $X2=0.3015 $Y2=0.072
r70 41 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.063 $X2=0.225 $Y2=0.072
r71 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.045 $X2=0.216 $Y2=0.063
r72 36 38 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r73 34 53 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r74 34 36 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.06 $Y2=0.135
r75 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r76 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.162 $Y2=0.036
r77 30 31 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.106
+ $Y=0.036 $X2=0.144 $Y2=0.036
r78 29 30 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.036 $X2=0.106 $Y2=0.036
r79 28 29 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.036 $X2=0.094 $Y2=0.036
r80 27 28 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.078 $Y2=0.036
r81 26 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.207 $Y=0.036 $X2=0.216 $Y2=0.045
r82 26 33 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.036 $X2=0.18 $Y2=0.036
r83 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.081
r84 18 53 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.135
r85 18 20 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.081
r86 17 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r87 17 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r88 13 48 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r89 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r90 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r91 5 38 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r92 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r93 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_XNOR2XP5_ASAP7_75T_R%B 2 7 10 13 15 24 VSS
c33 24 VSS 0.00331009f $X=0.136 $Y=0.135
c34 13 VSS 0.0170619f $X=0.297 $Y=0.135
c35 10 VSS 0.0656304f $X=0.297 $Y=0.0675
c36 2 VSS 0.0637809f $X=0.135 $Y=0.0675
r37 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r38 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r39 5 13 202.5 $w=1.6e-08 $l=1.62e-07 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.297 $Y2=0.135
r40 5 24 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r41 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r42 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_XNOR2XP5_ASAP7_75T_R%5 2 5 7 9 12 14 15 18 19 26 27 28 30 36 38 41 42
+ 43 44 49 53 54 VSS
c39 54 VSS 0.00205152f $X=0.171 $Y=0.198
c40 53 VSS 6.92425e-19 $X=0.405 $Y=0.1695
c41 49 VSS 4.12414e-19 $X=0.405 $Y=0.135
c42 47 VSS 9.17737e-19 $X=0.405 $Y=0.189
c43 46 VSS 1.56568e-19 $X=0.3915 $Y=0.198
c44 45 VSS 0.00223866f $X=0.387 $Y=0.198
c45 44 VSS 8.46035e-21 $X=0.36 $Y=0.198
c46 43 VSS 8.93197e-19 $X=0.342 $Y=0.198
c47 42 VSS 0.00278191f $X=0.256 $Y=0.198
c48 41 VSS 0.00149783f $X=0.207 $Y=0.198
c49 39 VSS 7.89418e-20 $X=0.396 $Y=0.198
c50 38 VSS 9.37882e-19 $X=0.171 $Y=0.225
c51 36 VSS 7.17067e-19 $X=0.171 $Y=0.1695
c52 30 VSS 0.00149298f $X=0.171 $Y=0.09
c53 28 VSS 2.52481e-19 $X=0.171 $Y=0.189
c54 27 VSS 0.00150698f $X=0.153 $Y=0.234
c55 26 VSS 0.00287092f $X=0.144 $Y=0.234
c56 21 VSS 0.00259482f $X=0.108 $Y=0.234
c57 19 VSS 0.00458651f $X=0.162 $Y=0.234
c58 18 VSS 0.00800631f $X=0.108 $Y=0.216
c59 14 VSS 6.05457e-19 $X=0.125 $Y=0.216
c60 12 VSS 0.0148676f $X=0.16 $Y=0.0675
c61 5 VSS 0.00172642f $X=0.405 $Y=0.135
c62 2 VSS 0.0664387f $X=0.405 $Y=0.0675
r63 52 53 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.15 $X2=0.405 $Y2=0.1695
r64 49 52 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.15
r65 47 53 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.1695
r66 45 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.387
+ $Y=0.198 $X2=0.3915 $Y2=0.198
r67 44 45 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.198 $X2=0.387 $Y2=0.198
r68 43 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r69 42 43 5.83951 $w=1.8e-08 $l=8.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.198 $X2=0.342 $Y2=0.198
r70 41 42 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.198 $X2=0.256 $Y2=0.198
r71 40 54 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.198 $X2=0.171 $Y2=0.198
r72 40 41 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.198 $X2=0.207 $Y2=0.198
r73 39 47 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.198 $X2=0.405 $Y2=0.189
r74 39 46 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.3915 $Y2=0.198
r75 37 54 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.207 $X2=0.171 $Y2=0.198
r76 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.207 $X2=0.171 $Y2=0.225
r77 35 36 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.15 $X2=0.171 $Y2=0.1695
r78 30 35 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.09 $X2=0.171 $Y2=0.15
r79 28 54 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.189 $X2=0.171 $Y2=0.198
r80 28 36 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.189 $X2=0.171 $Y2=0.1695
r81 26 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.153 $Y2=0.234
r82 21 26 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.144 $Y2=0.234
r83 19 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.234 $X2=0.171 $Y2=0.225
r84 19 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.153 $Y2=0.234
r85 18 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r86 15 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.216 $X2=0.108 $Y2=0.216
r87 14 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.216 $X2=0.108 $Y2=0.216
r88 12 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.171 $Y=0.09 $X2=0.171
+ $Y2=0.09
r89 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.16 $Y2=0.0675
r90 5 49 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r91 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r92 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_XNOR2XP5_ASAP7_75T_R%Y 1 6 9 11 14 24 29 31 36 39 VSS
c17 39 VSS 0.00328191f $X=0.45 $Y=0.036
c18 38 VSS 0.00277971f $X=0.459 $Y=0.036
c19 36 VSS 0.00294549f $X=0.432 $Y=0.036
c20 33 VSS 2.98008e-19 $X=0.459 $Y=0.216
c21 31 VSS 0.00258114f $X=0.459 $Y=0.121
c22 30 VSS 0.00102822f $X=0.459 $Y=0.063
c23 29 VSS 0.00366991f $X=0.457 $Y=0.135
c24 27 VSS 2.81452e-19 $X=0.459 $Y=0.225
c25 25 VSS 8.76814e-19 $X=0.423 $Y=0.234
c26 24 VSS 0.0162493f $X=0.414 $Y=0.234
c27 16 VSS 0.00607607f $X=0.45 $Y=0.234
c28 14 VSS 0.00704473f $X=0.43 $Y=0.2025
c29 9 VSS 0.00505246f $X=0.272 $Y=0.2025
c30 6 VSS 4.39464e-19 $X=0.287 $Y=0.2025
c31 4 VSS 3.25039e-19 $X=0.43 $Y=0.0675
r32 39 40 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r33 38 40 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r34 35 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r35 35 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r36 32 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.207 $X2=0.459 $Y2=0.216
r37 30 31 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.063 $X2=0.459 $Y2=0.121
r38 29 32 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.207
r39 29 31 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.121
r40 27 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.216
r41 26 38 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r42 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.063
r43 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.423 $Y2=0.234
r44 22 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.423 $Y2=0.234
r45 18 24 9.77778 $w=1.8e-08 $l=1.44e-07 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.414 $Y2=0.234
r46 16 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r47 16 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.432 $Y2=0.234
r48 14 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r49 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.43 $Y2=0.2025
r50 9 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r51 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.272 $Y2=0.2025
r52 4 36 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r53 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.43 $Y2=0.0675
.ends

.subckt PM_XNOR2XP5_ASAP7_75T_R%8 1 2 VSS
c1 1 VSS 0.0022361f $X=0.125 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends


* END of "./XNOR2xp5_ASAP7_75t_R.pex.sp.pex"
* 
.subckt XNOR2xp5_ASAP7_75t_R  VSS VDD A B Y
* 
* Y	Y
* B	B
* A	A
M0 N_8_M0_d N_A_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_5_M1_d N_B_M1_g N_8_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_B_M2_g noxref_6 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M3 noxref_6 N_A_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M4 N_Y_M4_d N_5_M4_g noxref_6 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 N_5_M5_d N_A_M5_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071 $Y=0.189
M6 VDD N_B_M6_g N_5_M6_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125 $Y=0.189
M7 noxref_9 N_B_M7_g N_Y_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M8 VDD N_A_M8_g noxref_9 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.162
M9 N_Y_M9_d N_5_M9_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.162
*
* 
* .include "XNOR2xp5_ASAP7_75t_R.pex.sp.XNOR2XP5_ASAP7_75T_R.pxi"
* BEGIN of "./XNOR2xp5_ASAP7_75t_R.pex.sp.XNOR2XP5_ASAP7_75T_R.pxi"
* File: XNOR2xp5_ASAP7_75t_R.pex.sp.XNOR2XP5_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:07:33 2017
* 
x_PM_XNOR2XP5_ASAP7_75T_R%A N_A_M0_g N_A_c_5_p N_A_M5_g N_A_M3_g N_A_c_6_p
+ N_A_M8_g N_A_c_9_p N_A_c_10_p N_A_c_7_p N_A_c_2_p N_A_c_18_p N_A_c_19_p A
+ N_A_c_20_p N_A_c_33_p N_A_c_8_p N_A_c_31_p N_A_c_4_p N_A_c_27_p N_A_c_28_p
+ N_A_c_14_p VSS PM_XNOR2XP5_ASAP7_75T_R%A
x_PM_XNOR2XP5_ASAP7_75T_R%B N_B_M1_g N_B_M6_g N_B_M2_g N_B_c_43_n N_B_M7_g B VSS
+ PM_XNOR2XP5_ASAP7_75T_R%B
x_PM_XNOR2XP5_ASAP7_75T_R%5 N_5_M4_g N_5_c_73_n N_5_M9_g N_5_M1_d N_5_c_74_n
+ N_5_M6_s N_5_M5_d N_5_c_89_n N_5_c_107_p N_5_c_90_n N_5_c_92_n N_5_c_93_n
+ N_5_c_78_n N_5_c_96_n N_5_c_103_p N_5_c_97_n N_5_c_81_n N_5_c_82_n N_5_c_83_n
+ N_5_c_85_n N_5_c_105_p N_5_c_99_n VSS PM_XNOR2XP5_ASAP7_75T_R%5
x_PM_XNOR2XP5_ASAP7_75T_R%Y N_Y_M4_d N_Y_M7_s N_Y_c_113_n N_Y_M9_d N_Y_c_119_n
+ N_Y_c_111_n Y N_Y_c_112_n N_Y_c_125_n N_Y_c_126_n VSS
+ PM_XNOR2XP5_ASAP7_75T_R%Y
x_PM_XNOR2XP5_ASAP7_75T_R%8 N_8_M1_s N_8_M0_d VSS PM_XNOR2XP5_ASAP7_75T_R%8
cc_1 N_A_M0_g N_B_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_M1_g 2.38942e-19 $X=0.144 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_3 N_A_M3_g N_B_M2_g 0.00323392f $X=0.351 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_4 N_A_c_4_p N_B_M2_g 2.9656e-19 $X=0.3015 $Y=0.072 $X2=0.297 $Y2=0.0675
cc_5 N_A_c_5_p N_B_c_43_n 8.12544e-19 $X=0.081 $Y=0.135 $X2=0.297 $Y2=0.135
cc_6 N_A_c_6_p N_B_c_43_n 0.00106649f $X=0.351 $Y=0.135 $X2=0.297 $Y2=0.135
cc_7 N_A_c_7_p N_B_c_43_n 3.32907e-19 $X=0.207 $Y=0.036 $X2=0.297 $Y2=0.135
cc_8 N_A_c_8_p N_B_c_43_n 0.00124812f $X=0.225 $Y=0.072 $X2=0.297 $Y2=0.135
cc_9 N_A_c_9_p B 2.57131e-19 $X=0.018 $Y=0.126 $X2=0.136 $Y2=0.135
cc_10 N_A_c_10_p B 2.3692e-19 $X=0.018 $Y=0.081 $X2=0.136 $Y2=0.135
cc_11 N_A_c_2_p B 0.00409303f $X=0.144 $Y=0.036 $X2=0.136 $Y2=0.135
cc_12 A B 4.29558e-19 $X=0.06 $Y=0.136 $X2=0.136 $Y2=0.135
cc_13 N_A_c_8_p B 3.32918e-19 $X=0.225 $Y=0.072 $X2=0.136 $Y2=0.135
cc_14 N_A_c_14_p B 8.13002e-19 $X=0.018 $Y=0.135 $X2=0.136 $Y2=0.135
cc_15 N_A_M3_g N_5_M4_g 0.00323392f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_16 N_A_c_6_p N_5_c_73_n 9.46013e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_17 N_A_c_7_p N_5_c_74_n 0.00142006f $X=0.207 $Y=0.036 $X2=0.297 $Y2=0.135
cc_18 N_A_c_18_p N_5_c_74_n 0.00161143f $X=0.162 $Y=0.036 $X2=0.297 $Y2=0.135
cc_19 N_A_c_19_p N_5_c_74_n 0.00130888f $X=0.18 $Y=0.036 $X2=0.297 $Y2=0.135
cc_20 N_A_c_20_p N_5_c_74_n 7.82924e-19 $X=0.216 $Y=0.063 $X2=0.297 $Y2=0.135
cc_21 N_A_c_19_p N_5_c_78_n 8.69266e-19 $X=0.18 $Y=0.036 $X2=0 $Y2=0
cc_22 N_A_c_8_p N_5_c_78_n 3.12063e-19 $X=0.225 $Y=0.072 $X2=0 $Y2=0
cc_23 N_A_c_14_p N_5_c_78_n 2.69986e-19 $X=0.018 $Y=0.135 $X2=0 $Y2=0
cc_24 N_A_c_8_p N_5_c_81_n 7.72163e-19 $X=0.225 $Y=0.072 $X2=0 $Y2=0
cc_25 N_A_c_4_p N_5_c_82_n 7.72163e-19 $X=0.3015 $Y=0.072 $X2=0 $Y2=0
cc_26 N_A_M3_g N_5_c_83_n 3.0688e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_A_c_27_p N_5_c_83_n 8.07817e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_28 N_A_c_28_p N_5_c_85_n 0.00118958f $X=0.351 $Y=0.128 $X2=0 $Y2=0
cc_29 VSS N_A_c_4_p 3.29233e-19 $X=0.3015 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_30 VSS N_A_c_7_p 7.39549e-19 $X=0.207 $Y=0.036 $X2=0.297 $Y2=0.135
cc_31 VSS N_A_c_31_p 4.94068e-19 $X=0.261 $Y=0.072 $X2=0.297 $Y2=0.135
cc_32 VSS N_A_c_4_p 0.00169244f $X=0.3015 $Y=0.072 $X2=0.297 $Y2=0.135
cc_33 VSS N_A_c_33_p 0.00158538f $X=0.342 $Y=0.072 $X2=0 $Y2=0
cc_34 VSS N_A_M3_g 2.34993e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_35 VSS N_A_c_7_p 8.81227e-19 $X=0.207 $Y=0.036 $X2=0 $Y2=0
cc_36 VSS N_A_c_4_p 0.00841951f $X=0.3015 $Y=0.072 $X2=0 $Y2=0
cc_37 N_A_M3_g N_Y_c_111_n 2.38303e-19 $X=0.351 $Y=0.0675 $X2=0.136 $Y2=0.135
cc_38 N_A_c_33_p N_Y_c_112_n 6.03287e-19 $X=0.342 $Y=0.072 $X2=0 $Y2=0
cc_39 N_B_M2_g N_5_M4_g 2.34385e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_40 N_B_c_43_n N_5_c_74_n 0.00369057f $X=0.297 $Y=0.135 $X2=0.351 $Y2=0.135
cc_41 B N_5_c_74_n 5.10449e-19 $X=0.136 $Y=0.135 $X2=0.351 $Y2=0.135
cc_42 B N_5_c_89_n 0.00184579f $X=0.136 $Y=0.135 $X2=0.018 $Y2=0.126
cc_43 N_B_M1_g N_5_c_90_n 2.35623e-19 $X=0.135 $Y=0.0675 $X2=0.207 $Y2=0.036
cc_44 B N_5_c_90_n 0.00374777f $X=0.136 $Y=0.135 $X2=0.207 $Y2=0.036
cc_45 N_B_c_43_n N_5_c_92_n 2.91977e-19 $X=0.297 $Y=0.135 $X2=0.027 $Y2=0.036
cc_46 B N_5_c_93_n 0.00183916f $X=0.136 $Y=0.135 $X2=0.078 $Y2=0.036
cc_47 N_B_c_43_n N_5_c_78_n 0.00250832f $X=0.297 $Y=0.135 $X2=0.106 $Y2=0.036
cc_48 B N_5_c_78_n 0.00551748f $X=0.136 $Y=0.135 $X2=0.106 $Y2=0.036
cc_49 B N_5_c_96_n 0.00183916f $X=0.136 $Y=0.135 $X2=0.06 $Y2=0.136
cc_50 N_B_c_43_n N_5_c_97_n 0.00135939f $X=0.297 $Y=0.135 $X2=0.216 $Y2=0.063
cc_51 N_B_M2_g N_5_c_82_n 4.09048e-19 $X=0.297 $Y=0.0675 $X2=0.225 $Y2=0.072
cc_52 B N_5_c_99_n 0.00183916f $X=0.136 $Y=0.135 $X2=0.064 $Y2=0.135
cc_53 VSS N_B_c_43_n 6.8292e-19 $X=0.297 $Y=0.135 $X2=0.351 $Y2=0.135
cc_54 VSS N_B_M2_g 2.65491e-19 $X=0.297 $Y=0.0675 $X2=0.018 $Y2=0.126
cc_55 N_B_c_43_n N_Y_c_113_n 6.8292e-19 $X=0.297 $Y=0.135 $X2=0.351 $Y2=0.0675
cc_56 N_B_M2_g N_Y_c_111_n 2.65491e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_57 B N_8_M1_s 2.02285e-19 $X=0.136 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_58 VSS N_5_c_74_n 0.0022753f $X=0.16 $Y=0.0675 $X2=0.351 $Y2=0.135
cc_59 N_5_c_82_n N_Y_M7_s 3.29233e-19 $X=0.342 $Y=0.198 $X2=0.081 $Y2=0.216
cc_60 N_5_c_96_n N_Y_c_113_n 5.55768e-19 $X=0.171 $Y=0.1695 $X2=0.351 $Y2=0.0675
cc_61 N_5_c_103_p N_Y_c_113_n 2.38811e-19 $X=0.171 $Y=0.225 $X2=0.351 $Y2=0.0675
cc_62 N_5_c_82_n N_Y_c_113_n 0.00284111f $X=0.342 $Y=0.198 $X2=0.351 $Y2=0.0675
cc_63 N_5_c_105_p N_Y_c_119_n 0.00135952f $X=0.405 $Y=0.1695 $X2=0.351
+ $Y2=0.2025
cc_64 N_5_M4_g N_Y_c_111_n 2.34993e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_65 N_5_c_107_p N_Y_c_111_n 5.49907e-19 $X=0.162 $Y=0.234 $X2=0 $Y2=0
cc_66 N_5_c_82_n N_Y_c_111_n 0.0133208f $X=0.342 $Y=0.198 $X2=0 $Y2=0
cc_67 N_5_c_85_n Y 0.0034418f $X=0.405 $Y=0.135 $X2=0.094 $Y2=0.036
cc_68 VSS N_5_c_82_n 5.15356e-19 $X=0.342 $Y=0.198 $X2=0.081 $Y2=0.0675
cc_69 VSS N_Y_c_113_n 0.00169333f $X=0.27 $Y=0.036 $X2=0.351 $Y2=0.0675
cc_70 VSS N_Y_c_125_n 0.00395939f $X=0.378 $Y=0.036 $X2=0.06 $Y2=0.136
cc_71 VSS N_Y_c_126_n 6.52162e-19 $X=0.378 $Y=0.036 $X2=0 $Y2=0
cc_72 VSS N_Y_c_111_n 3.33359e-19 $X=0.414 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./XNOR2xp5_ASAP7_75t_R.pex.sp.XNOR2XP5_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: MAJIxp5_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:36:51 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "MAJIxp5_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./MAJIxp5_ASAP7_75t_R.pex.sp.pex"
* File: MAJIxp5_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:36:51 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_MAJIXP5_ASAP7_75T_R%B 2 5 7 10 13 15 27 29 33 36 37 38 41 43 45 49
+ VSS
c31 49 VSS 0.00757186f $X=0.018 $Y=0.135
c32 45 VSS 0.00113888f $X=0.243 $Y=0.135
c33 43 VSS 3.12554e-20 $X=0.198 $Y=0.135
c34 42 VSS 6.79449e-19 $X=0.189 $Y=0.1765
c35 41 VSS 3.30052e-19 $X=0.189 $Y=0.164
c36 40 VSS 6.05864e-19 $X=0.189 $Y=0.189
c37 38 VSS 8.46035e-21 $X=0.144 $Y=0.198
c38 37 VSS 5.71746e-19 $X=0.126 $Y=0.198
c39 36 VSS 4.40637e-21 $X=0.095 $Y=0.198
c40 35 VSS 0.00502565f $X=0.094 $Y=0.198
c41 34 VSS 0.00194397f $X=0.027 $Y=0.198
c42 33 VSS 0.00237121f $X=0.18 $Y=0.198
c43 29 VSS 0.00350979f $X=0.081 $Y=0.135
c44 24 VSS 5.58698e-19 $X=0.018 $Y=0.1765
c45 23 VSS 8.46985e-19 $X=0.018 $Y=0.164
c46 22 VSS 4.47174e-19 $X=0.018 $Y=0.189
c47 13 VSS 0.00123068f $X=0.243 $Y=0.135
c48 10 VSS 0.0599814f $X=0.243 $Y=0.0675
c49 5 VSS 0.00262838f $X=0.081 $Y=0.135
c50 2 VSS 0.0597899f $X=0.081 $Y=0.0675
r51 43 45 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.135 $X2=0.243 $Y2=0.135
r52 41 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.1765
r53 40 42 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.1765
r54 39 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.144 $X2=0.198 $Y2=0.135
r55 39 41 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.164
r56 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.198 $X2=0.144 $Y2=0.198
r57 36 37 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.198 $X2=0.126 $Y2=0.198
r58 35 36 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.198 $X2=0.095 $Y2=0.198
r59 34 35 4.54938 $w=1.8e-08 $l=6.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.198 $X2=0.094 $Y2=0.198
r60 33 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.198 $X2=0.189 $Y2=0.189
r61 33 38 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.198 $X2=0.144 $Y2=0.198
r62 27 29 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.063
+ $Y=0.135 $X2=0.081 $Y2=0.135
r63 25 49 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r64 25 27 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.063 $Y2=0.135
r65 23 24 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.164 $X2=0.018 $Y2=0.1765
r66 22 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.189 $X2=0.027 $Y2=0.198
r67 22 24 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.189 $X2=0.018 $Y2=0.1765
r68 21 49 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.135
r69 21 23 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.144 $X2=0.018 $Y2=0.164
r70 13 45 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r71 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r72 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r73 5 29 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r74 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r75 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_MAJIXP5_ASAP7_75T_R%C 2 7 10 13 15 19 23 26 VSS
c26 26 VSS 1.44512e-20 $X=0.135 $Y=0.1305
c27 23 VSS 5.26174e-19 $X=0.135 $Y=0.135
c28 19 VSS 0.00354745f $X=0.138 $Y=0.116
c29 13 VSS 0.00960045f $X=0.189 $Y=0.135
c30 10 VSS 0.0609113f $X=0.189 $Y=0.0675
c31 2 VSS 0.0587452f $X=0.135 $Y=0.0675
r32 25 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.126 $X2=0.135 $Y2=0.1305
r33 23 26 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.1305
r34 19 25 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.116 $X2=0.135 $Y2=0.126
r35 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r36 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
r37 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.189 $Y2=0.135
r38 5 23 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r39 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r40 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_MAJIXP5_ASAP7_75T_R%A 2 5 7 10 13 16 VSS
c14 16 VSS 1.44512e-20 $X=0.297 $Y=0.1305
c15 13 VSS 3.17034e-19 $X=0.297 $Y=0.135
c16 10 VSS 3.4868e-19 $X=0.296 $Y=0.116
c17 5 VSS 0.00170066f $X=0.297 $Y=0.135
c18 2 VSS 0.0634749f $X=0.297 $Y=0.0675
r19 15 16 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.297 $Y2=0.1305
r20 13 16 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.1305
r21 10 15 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.116 $X2=0.297 $Y2=0.126
r22 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r23 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r24 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
.ends

.subckt PM_MAJIXP5_ASAP7_75T_R%6 1 2 6 9 13 18 19 21 22 23 VSS
c17 23 VSS 0.0027128f $X=0.2895 $Y=0.036
c18 22 VSS 0.00624731f $X=0.255 $Y=0.036
c19 21 VSS 0.00708303f $X=0.18 $Y=0.036
c20 20 VSS 0.00248077f $X=0.126 $Y=0.036
c21 19 VSS 0.00236594f $X=0.324 $Y=0.036
c22 18 VSS 0.00501912f $X=0.324 $Y=0.036
c23 13 VSS 0.00980178f $X=0.108 $Y=0.036
c24 12 VSS 0.00202752f $X=0.108 $Y=0.036
c25 9 VSS 2.69461e-19 $X=0.322 $Y=0.0675
c26 1 VSS 6.11334e-19 $X=0.125 $Y=0.0675
r27 22 23 2.34259 $w=1.8e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.255
+ $Y=0.036 $X2=0.2895 $Y2=0.036
r28 21 22 5.09259 $w=1.8e-08 $l=7.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.036 $X2=0.255 $Y2=0.036
r29 20 21 3.66667 $w=1.8e-08 $l=5.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.18 $Y2=0.036
r30 18 23 2.34259 $w=1.8e-08 $l=3.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.036 $X2=0.2895 $Y2=0.036
r31 18 19 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.036 $X2=0.324
+ $Y2=0.036
r32 12 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r33 12 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r34 9 19 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.324
+ $Y=0.0675 $X2=0.324 $Y2=0.036
r35 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.0675 $X2=0.322 $Y2=0.0675
r36 5 13 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r37 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
r38 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.108 $Y2=0.0675
.ends

.subckt PM_MAJIXP5_ASAP7_75T_R%7 1 2 5 6 9 16 18 19 VSS
c15 19 VSS 0.00476966f $X=0.255 $Y=0.234
c16 18 VSS 0.0122251f $X=0.198 $Y=0.234
c17 16 VSS 0.00773728f $X=0.324 $Y=0.234
c18 9 VSS 0.0026354f $X=0.322 $Y=0.2025
c19 5 VSS 0.00940011f $X=0.108 $Y=0.2025
c20 1 VSS 6.64569e-19 $X=0.125 $Y=0.2025
r21 18 19 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.234 $X2=0.255 $Y2=0.234
r22 16 19 4.68518 $w=1.8e-08 $l=6.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.234 $X2=0.255 $Y2=0.234
r23 12 18 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.198 $Y2=0.234
r24 9 16 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.324 $Y=0.234 $X2=0.324
+ $Y2=0.234
r25 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.307
+ $Y=0.2025 $X2=0.322 $Y2=0.2025
r26 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r27 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.091
+ $Y=0.2025 $X2=0.108 $Y2=0.2025
r28 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.2025 $X2=0.108 $Y2=0.2025
.ends

.subckt PM_MAJIXP5_ASAP7_75T_R%Y 1 2 5 6 7 10 13 18 19 20 24 30 31 36 37 38 VSS
c21 40 VSS 6.00064e-19 $X=0.352 $Y=0.1765
c22 38 VSS 5.78177e-19 $X=0.352 $Y=0.1185
c23 37 VSS 0.00122318f $X=0.352 $Y=0.106
c24 36 VSS 0.00208008f $X=0.354 $Y=0.131
c25 34 VSS 6.42831e-19 $X=0.352 $Y=0.189
c26 32 VSS 1.72289e-19 $X=0.3405 $Y=0.198
c27 31 VSS 3.67948e-19 $X=0.338 $Y=0.198
c28 30 VSS 8.46035e-21 $X=0.306 $Y=0.198
c29 29 VSS 3.18436e-19 $X=0.288 $Y=0.198
c30 24 VSS 2.24252e-19 $X=0.269 $Y=0.198
c31 22 VSS 0.00210789f $X=0.343 $Y=0.198
c32 21 VSS 1.72289e-19 $X=0.3405 $Y=0.072
c33 20 VSS 3.67948e-19 $X=0.338 $Y=0.072
c34 19 VSS 8.46035e-21 $X=0.306 $Y=0.072
c35 18 VSS 3.18436e-19 $X=0.288 $Y=0.072
c36 13 VSS 2.63633e-19 $X=0.269 $Y=0.072
c37 11 VSS 0.00210789f $X=0.343 $Y=0.072
c38 10 VSS 0.00350219f $X=0.27 $Y=0.2025
c39 6 VSS 6.10538e-19 $X=0.287 $Y=0.2025
c40 5 VSS 0.00366232f $X=0.27 $Y=0.0675
c41 1 VSS 6.12399e-19 $X=0.287 $Y=0.0675
r42 39 40 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.352
+ $Y=0.164 $X2=0.352 $Y2=0.1765
r43 37 38 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.352
+ $Y=0.106 $X2=0.352 $Y2=0.1185
r44 36 39 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.352
+ $Y=0.131 $X2=0.352 $Y2=0.164
r45 36 38 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.352
+ $Y=0.131 $X2=0.352 $Y2=0.1185
r46 34 40 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.352
+ $Y=0.189 $X2=0.352 $Y2=0.1765
r47 33 37 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.352
+ $Y=0.081 $X2=0.352 $Y2=0.106
r48 31 32 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.198 $X2=0.3405 $Y2=0.198
r49 30 31 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.198 $X2=0.338 $Y2=0.198
r50 29 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.198 $X2=0.306 $Y2=0.198
r51 24 29 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.269
+ $Y=0.198 $X2=0.288 $Y2=0.198
r52 22 34 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.343 $Y=0.198 $X2=0.352 $Y2=0.189
r53 22 32 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.343
+ $Y=0.198 $X2=0.3405 $Y2=0.198
r54 20 21 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.338
+ $Y=0.072 $X2=0.3405 $Y2=0.072
r55 19 20 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.306
+ $Y=0.072 $X2=0.338 $Y2=0.072
r56 18 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.288
+ $Y=0.072 $X2=0.306 $Y2=0.072
r57 13 18 1.29012 $w=1.8e-08 $l=1.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.269
+ $Y=0.072 $X2=0.288 $Y2=0.072
r58 11 33 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.343 $Y=0.072 $X2=0.352 $Y2=0.081
r59 11 21 0.169753 $w=1.8e-08 $l=2.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.343
+ $Y=0.072 $X2=0.3405 $Y2=0.072
r60 10 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.269 $Y=0.198 $X2=0.269
+ $Y2=0.198
r61 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r62 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r63 5 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.269 $Y=0.072 $X2=0.269
+ $Y2=0.072
r64 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.253
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
r65 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.0675 $X2=0.27 $Y2=0.0675
.ends

.subckt PM_MAJIXP5_ASAP7_75T_R%9 1 2 VSS
c2 1 VSS 0.00183233f $X=0.233 $Y=0.0675
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.0675 $X2=0.199 $Y2=0.0675
.ends

.subckt PM_MAJIXP5_ASAP7_75T_R%10 1 2 VSS
c2 1 VSS 0.00183233f $X=0.233 $Y=0.2025
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.233
+ $Y=0.2025 $X2=0.199 $Y2=0.2025
.ends


* END of "./MAJIxp5_ASAP7_75t_R.pex.sp.pex"
* 
.subckt MAJIxp5_ASAP7_75t_R  VSS VDD B C A Y
* 
* Y	Y
* A	A
* C	C
* B	B
M0 N_6_M0_d N_B_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 VSS N_C_M1_g N_6_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.027
M2 N_9_M2_d N_C_M2_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179 $Y=0.027
M3 N_Y_M3_d N_B_M3_g N_9_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 N_6_M4_d N_A_M4_g N_Y_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.027
M5 N_7_M5_d N_B_M5_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
M6 VDD N_C_M6_g N_7_M6_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125 $Y=0.162
M7 N_10_M7_d N_C_M7_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M8 N_Y_M8_d N_B_M8_g N_10_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M9 N_7_M9_d N_A_M9_g N_Y_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
*
* 
* .include "MAJIxp5_ASAP7_75t_R.pex.sp.MAJIXP5_ASAP7_75T_R.pxi"
* BEGIN of "./MAJIxp5_ASAP7_75t_R.pex.sp.MAJIXP5_ASAP7_75T_R.pxi"
* File: MAJIxp5_ASAP7_75t_R.pex.sp.MAJIXP5_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:36:51 2017
* 
x_PM_MAJIXP5_ASAP7_75T_R%B N_B_M0_g N_B_c_7_p N_B_M5_g N_B_M3_g N_B_c_8_p
+ N_B_M8_g B N_B_c_16_p N_B_c_9_p N_B_c_25_p N_B_c_24_p N_B_c_3_p N_B_c_10_p
+ N_B_c_6_p N_B_c_12_p N_B_c_13_p VSS PM_MAJIXP5_ASAP7_75T_R%B
x_PM_MAJIXP5_ASAP7_75T_R%C N_C_M1_g N_C_M6_g N_C_M2_g N_C_c_38_n N_C_M7_g C
+ N_C_c_45_n N_C_c_47_n VSS PM_MAJIXP5_ASAP7_75T_R%C
x_PM_MAJIXP5_ASAP7_75T_R%A N_A_M4_g N_A_c_59_n N_A_M9_g A N_A_c_60_n N_A_c_61_n
+ VSS PM_MAJIXP5_ASAP7_75T_R%A
x_PM_MAJIXP5_ASAP7_75T_R%6 N_6_M1_s N_6_M0_d N_6_M4_d N_6_c_85_p N_6_c_74_n
+ N_6_c_78_n N_6_c_80_p N_6_c_75_n N_6_c_72_n N_6_c_82_p VSS
+ PM_MAJIXP5_ASAP7_75T_R%6
x_PM_MAJIXP5_ASAP7_75T_R%7 N_7_M6_s N_7_M5_d N_7_c_89_n N_7_M9_d N_7_c_97_n
+ N_7_c_95_n N_7_c_90_n N_7_c_91_n VSS PM_MAJIXP5_ASAP7_75T_R%7
x_PM_MAJIXP5_ASAP7_75T_R%Y N_Y_M4_s N_Y_M3_d N_Y_c_113_n N_Y_M9_s N_Y_M8_d
+ N_Y_c_104_n N_Y_c_106_n N_Y_c_116_n N_Y_c_107_n N_Y_c_117_n N_Y_c_105_n
+ N_Y_c_109_n N_Y_c_123_n Y N_Y_c_119_n N_Y_c_112_n VSS PM_MAJIXP5_ASAP7_75T_R%Y
x_PM_MAJIXP5_ASAP7_75T_R%9 N_9_M3_s N_9_M2_d VSS PM_MAJIXP5_ASAP7_75T_R%9
x_PM_MAJIXP5_ASAP7_75T_R%10 N_10_M8_s N_10_M7_d VSS PM_MAJIXP5_ASAP7_75T_R%10
cc_1 N_B_M0_g N_C_M1_g 0.00316373f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_B_M3_g N_C_M1_g 2.13359e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_3 N_B_c_3_p N_C_M1_g 2.76185e-19 $X=0.144 $Y=0.198 $X2=0.135 $Y2=0.0675
cc_4 N_B_M0_g N_C_M2_g 2.13359e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_5 N_B_M3_g N_C_M2_g 0.00341068f $X=0.243 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_6 N_B_c_6_p N_C_M2_g 3.47593e-19 $X=0.198 $Y=0.135 $X2=0.189 $Y2=0.0675
cc_7 N_B_c_7_p N_C_c_38_n 0.00122296f $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.135
cc_8 N_B_c_8_p N_C_c_38_n 0.00148337f $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.135
cc_9 N_B_c_9_p N_C_c_38_n 4.36331e-19 $X=0.18 $Y=0.198 $X2=0.189 $Y2=0.135
cc_10 N_B_c_10_p N_C_c_38_n 4.74454e-19 $X=0.189 $Y=0.164 $X2=0.189 $Y2=0.135
cc_11 N_B_c_6_p N_C_c_38_n 0.00147533f $X=0.198 $Y=0.135 $X2=0.189 $Y2=0.135
cc_12 N_B_c_12_p N_C_c_38_n 3.58003e-19 $X=0.243 $Y=0.135 $X2=0.189 $Y2=0.135
cc_13 N_B_c_13_p C 6.03035e-19 $X=0.018 $Y=0.135 $X2=0.138 $Y2=0.116
cc_14 N_B_c_3_p N_C_c_45_n 0.00123353f $X=0.144 $Y=0.198 $X2=0.135 $Y2=0.135
cc_15 N_B_c_10_p N_C_c_45_n 8.0975e-19 $X=0.189 $Y=0.164 $X2=0.135 $Y2=0.135
cc_16 N_B_c_16_p N_C_c_47_n 8.78098e-19 $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.1305
cc_17 N_B_c_6_p N_C_c_47_n 8.0975e-19 $X=0.198 $Y=0.135 $X2=0.135 $Y2=0.1305
cc_18 N_B_M3_g N_A_M4_g 0.00355599f $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_19 N_B_c_8_p N_A_c_59_n 0.00118985f $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.135
cc_20 N_B_c_10_p N_A_c_60_n 4.37585e-19 $X=0.189 $Y=0.164 $X2=0.189 $Y2=0.135
cc_21 N_B_c_12_p N_A_c_61_n 8.76278e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_22 N_B_M3_g N_6_c_72_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_23 N_B_c_6_p N_6_c_72_n 0.00162183f $X=0.198 $Y=0.135 $X2=0.135 $Y2=0.135
cc_24 N_B_c_24_p N_7_c_89_n 0.00233206f $X=0.126 $Y=0.198 $X2=0.135 $Y2=0.135
cc_25 N_B_c_25_p N_7_c_90_n 0.00913202f $X=0.095 $Y=0.198 $X2=0.135 $Y2=0.116
cc_26 N_B_M3_g N_7_c_91_n 4.28653e-19 $X=0.243 $Y=0.0675 $X2=0.138 $Y2=0.116
cc_27 N_B_c_12_p N_7_c_91_n 0.00121779f $X=0.243 $Y=0.135 $X2=0.138 $Y2=0.116
cc_28 N_B_c_10_p N_Y_c_104_n 4.22488e-19 $X=0.189 $Y=0.164 $X2=0.189 $Y2=0.0675
cc_29 N_B_c_9_p N_Y_c_105_n 6.52936e-19 $X=0.18 $Y=0.198 $X2=0.135 $Y2=0.135
cc_30 N_B_c_12_p N_9_M3_s 4.4685e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_31 N_B_c_12_p N_10_M8_s 4.4685e-19 $X=0.243 $Y=0.135 $X2=0.135 $Y2=0.0675
cc_32 N_C_M2_g N_A_M4_g 2.82885e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_33 C A 2.40891e-19 $X=0.138 $Y=0.116 $X2=0.243 $Y2=0.0675
cc_34 C N_6_c_74_n 0.0015758f $X=0.138 $Y=0.116 $X2=0.243 $Y2=0.135
cc_35 N_C_M1_g N_6_c_75_n 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0.018 $Y2=0.144
cc_36 C N_6_c_75_n 0.00509708f $X=0.138 $Y=0.116 $X2=0.018 $Y2=0.144
cc_37 N_C_M2_g N_6_c_72_n 4.01862e-19 $X=0.189 $Y=0.0675 $X2=0.018 $Y2=0.189
cc_38 N_C_M1_g N_7_c_90_n 2.38303e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_C_M2_g N_7_c_90_n 2.34993e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_40 C N_Y_c_106_n 4.57752e-19 $X=0.138 $Y=0.116 $X2=0.243 $Y2=0.135
cc_41 N_A_M4_g N_6_c_78_n 2.15135e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_42 N_A_M4_g N_7_c_95_n 2.38303e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_43 N_A_M4_g N_Y_c_107_n 2.76185e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_44 A N_Y_c_107_n 0.00122099f $X=0.296 $Y=0.116 $X2=0 $Y2=0
cc_45 N_A_M4_g N_Y_c_109_n 2.76185e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_46 N_A_c_60_n N_Y_c_109_n 0.00122099f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_47 N_A_c_60_n Y 0.00138659f $X=0.297 $Y=0.135 $X2=0.095 $Y2=0.198
cc_48 A N_Y_c_112_n 0.00138659f $X=0.296 $Y=0.116 $X2=0.144 $Y2=0.198
cc_49 N_6_c_74_n N_7_c_89_n 0.00138157f $X=0.108 $Y=0.036 $X2=0.081 $Y2=0.135
cc_50 N_6_c_80_p N_7_c_97_n 0.00169333f $X=0.324 $Y=0.036 $X2=0.243 $Y2=0.0675
cc_51 N_6_c_80_p N_Y_c_113_n 0.00376964f $X=0.324 $Y=0.036 $X2=0.081 $Y2=0.135
cc_52 N_6_c_82_p N_Y_c_113_n 0.00284083f $X=0.2895 $Y=0.036 $X2=0.081 $Y2=0.135
cc_53 N_6_c_82_p N_Y_c_106_n 0.00353979f $X=0.2895 $Y=0.036 $X2=0.243 $Y2=0.135
cc_54 N_6_c_78_n N_Y_c_116_n 0.00353979f $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_55 N_6_c_85_p N_Y_c_117_n 2.45503e-19 $X=0.322 $Y=0.0675 $X2=0 $Y2=0
cc_56 N_6_c_80_p N_Y_c_117_n 0.00253233f $X=0.324 $Y=0.036 $X2=0 $Y2=0
cc_57 N_6_c_80_p N_Y_c_119_n 3.42083e-19 $X=0.324 $Y=0.036 $X2=0.126 $Y2=0.198
cc_58 N_6_c_72_n N_9_M3_s 4.63074e-19 $X=0.255 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_59 N_7_c_97_n N_Y_c_104_n 0.00376954f $X=0.322 $Y=0.2025 $X2=0.243 $Y2=0.0675
cc_60 N_7_c_95_n N_Y_c_104_n 0.00284083f $X=0.324 $Y=0.234 $X2=0.243 $Y2=0.0675
cc_61 N_7_c_95_n N_Y_c_105_n 0.00707944f $X=0.324 $Y=0.234 $X2=0.018 $Y2=0.1765
cc_62 N_7_c_97_n N_Y_c_123_n 0.00277783f $X=0.322 $Y=0.2025 $X2=0 $Y2=0
cc_63 N_7_c_97_n Y 3.32646e-19 $X=0.322 $Y=0.2025 $X2=0.095 $Y2=0.198
cc_64 N_7_c_91_n N_10_M8_s 4.63074e-19 $X=0.255 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./MAJIxp5_ASAP7_75t_R.pex.sp.MAJIXP5_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: MAJx2_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:37:13 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "MAJx2_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./MAJx2_ASAP7_75t_R.pex.sp.pex"
* File: MAJx2_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:37:13 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_MAJX2_ASAP7_75T_R%A 2 5 7 10 13 16 VSS
c13 16 VSS 1.44512e-20 $X=0.081 $Y=0.1305
c14 13 VSS 3.17034e-19 $X=0.081 $Y=0.135
c15 10 VSS 3.4868e-19 $X=0.082 $Y=0.116
c16 5 VSS 0.00170659f $X=0.081 $Y=0.135
c17 2 VSS 0.0634749f $X=0.081 $Y=0.0675
r18 15 16 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r19 13 16 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r20 10 15 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.116 $X2=0.081 $Y2=0.126
r21 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_MAJX2_ASAP7_75T_R%B 2 5 7 10 13 15 17 19 26 29 31 32 33 34 38 41 VSS
c41 41 VSS 0.00240496f $X=0.297 $Y=0.135
c42 39 VSS 0.00104593f $X=0.324 $Y=0.164
c43 38 VSS 5.33988e-20 $X=0.324 $Y=0.149
c44 37 VSS 0.00143326f $X=0.324 $Y=0.189
c45 35 VSS 4.40637e-21 $X=0.284 $Y=0.198
c46 34 VSS 5.22651e-19 $X=0.283 $Y=0.198
c47 33 VSS 8.46035e-21 $X=0.252 $Y=0.198
c48 32 VSS 0.0021192f $X=0.234 $Y=0.198
c49 29 VSS 3.26268e-19 $X=0.198 $Y=0.198
c50 28 VSS 0.00361589f $X=0.315 $Y=0.198
c51 27 VSS 6.38949e-19 $X=0.189 $Y=0.1765
c52 26 VSS 3.30052e-19 $X=0.189 $Y=0.164
c53 25 VSS 5.59921e-19 $X=0.189 $Y=0.189
c54 19 VSS 4.29576e-19 $X=0.135 $Y=0.135
c55 17 VSS 5.234e-19 $X=0.18 $Y=0.135
c56 13 VSS 0.00100977f $X=0.297 $Y=0.135
c57 10 VSS 0.0587302f $X=0.297 $Y=0.0675
c58 5 VSS 0.00119949f $X=0.135 $Y=0.135
c59 2 VSS 0.0599814f $X=0.135 $Y=0.0675
r60 41 43 1.32 $w=2.5e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.324 $Y2=0.126
r61 38 39 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.149 $X2=0.324 $Y2=0.164
r62 37 39 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.189 $X2=0.324 $Y2=0.164
r63 36 43 0.266695 $w=2.5e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.144 $X2=0.324 $Y2=0.126
r64 36 38 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.144 $X2=0.324 $Y2=0.149
r65 34 35 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.283
+ $Y=0.198 $X2=0.284 $Y2=0.198
r66 33 34 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.283 $Y2=0.198
r67 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.252 $Y2=0.198
r68 31 35 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.289
+ $Y=0.198 $X2=0.284 $Y2=0.198
r69 29 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.198 $X2=0.234 $Y2=0.198
r70 28 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.315 $Y=0.198 $X2=0.324 $Y2=0.189
r71 28 31 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.315
+ $Y=0.198 $X2=0.289 $Y2=0.198
r72 26 27 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.1765
r73 25 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.189 $X2=0.198 $Y2=0.198
r74 25 27 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.1765
r75 24 26 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.164
r76 17 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r77 17 19 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.135 $Y2=0.135
r78 13 41 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r79 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r80 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r81 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r82 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r83 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_MAJX2_ASAP7_75T_R%C 2 7 10 13 15 18 21 24 VSS
c28 24 VSS 1.44512e-20 $X=0.243 $Y=0.1305
c29 21 VSS 2.8151e-19 $X=0.243 $Y=0.135
c30 18 VSS 3.77468e-19 $X=0.24 $Y=0.116
c31 13 VSS 0.00942605f $X=0.243 $Y=0.135
c32 10 VSS 0.0583526f $X=0.243 $Y=0.0675
c33 2 VSS 0.0609465f $X=0.189 $Y=0.0675
r34 23 24 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.1305
r35 21 24 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.1305
r36 18 23 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.116 $X2=0.243 $Y2=0.126
r37 13 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r38 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r39 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r40 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r41 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r42 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_MAJX2_ASAP7_75T_R%6 2 7 10 13 15 17 18 21 22 23 26 29 30 31 37 38 41
+ 43 44 45 46 47 49 52 55 56 62 64 65 VSS
c53 65 VSS 2.72731e-19 $X=0.377 $Y=0.1205
c54 64 VSS 9.18711e-19 $X=0.377 $Y=0.106
c55 62 VSS 6.39194e-19 $X=0.377 $Y=0.135
c56 57 VSS 1.05074e-19 $X=0.0995 $Y=0.198
c57 56 VSS 8.46035e-21 $X=0.09 $Y=0.198
c58 55 VSS 4.41002e-19 $X=0.072 $Y=0.198
c59 54 VSS 3.80317e-19 $X=0.04 $Y=0.198
c60 52 VSS 4.23036e-19 $X=0.109 $Y=0.198
c61 50 VSS 0.00199912f $X=0.035 $Y=0.198
c62 49 VSS 1.36714e-20 $X=0.366 $Y=0.072
c63 48 VSS 0.00184044f $X=0.364 $Y=0.072
c64 47 VSS 0.0019689f $X=0.333 $Y=0.072
c65 46 VSS 0.0016201f $X=0.315 $Y=0.072
c66 45 VSS 4.40637e-21 $X=0.284 $Y=0.072
c67 44 VSS 5.22651e-19 $X=0.283 $Y=0.072
c68 43 VSS 8.46035e-21 $X=0.252 $Y=0.072
c69 42 VSS 0.00304109f $X=0.234 $Y=0.072
c70 41 VSS 2.51834e-19 $X=0.198 $Y=0.072
c71 40 VSS 2.61464e-19 $X=0.121 $Y=0.072
c72 39 VSS 1.05074e-19 $X=0.0995 $Y=0.072
c73 38 VSS 8.46035e-21 $X=0.09 $Y=0.072
c74 37 VSS 2.66799e-19 $X=0.072 $Y=0.072
c75 36 VSS 2.38309e-19 $X=0.04 $Y=0.072
c76 32 VSS 0.00206328f $X=0.035 $Y=0.072
c77 31 VSS 1.23404e-19 $X=0.368 $Y=0.072
c78 30 VSS 0.00267929f $X=0.026 $Y=0.164
c79 29 VSS 0.0010539f $X=0.026 $Y=0.106
c80 28 VSS 0.00124616f $X=0.026 $Y=0.189
c81 26 VSS 0.00350219f $X=0.108 $Y=0.2025
c82 22 VSS 6.10767e-19 $X=0.125 $Y=0.2025
c83 21 VSS 0.00357941f $X=0.108 $Y=0.0675
c84 17 VSS 6.22718e-19 $X=0.125 $Y=0.0675
c85 13 VSS 0.00452707f $X=0.405 $Y=0.135
c86 10 VSS 0.0639847f $X=0.405 $Y=0.0675
c87 2 VSS 0.0613943f $X=0.351 $Y=0.0675
r88 64 65 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.377
+ $Y=0.106 $X2=0.377 $Y2=0.1205
r89 62 65 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.377
+ $Y=0.135 $X2=0.377 $Y2=0.1205
r90 62 63 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.377 $Y=0.135 $X2=0.377
+ $Y2=0.135
r91 60 64 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.377
+ $Y=0.081 $X2=0.377 $Y2=0.106
r92 56 57 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.198 $X2=0.0995 $Y2=0.198
r93 55 56 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.198 $X2=0.09 $Y2=0.198
r94 54 55 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.198 $X2=0.072 $Y2=0.198
r95 52 57 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.198 $X2=0.0995 $Y2=0.198
r96 50 54 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.035
+ $Y=0.198 $X2=0.04 $Y2=0.198
r97 48 49 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.364
+ $Y=0.072 $X2=0.366 $Y2=0.072
r98 47 48 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.072 $X2=0.364 $Y2=0.072
r99 46 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.315
+ $Y=0.072 $X2=0.333 $Y2=0.072
r100 45 46 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.072 $X2=0.315 $Y2=0.072
r101 44 45 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.283
+ $Y=0.072 $X2=0.284 $Y2=0.072
r102 43 44 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.072 $X2=0.283 $Y2=0.072
r103 42 43 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.252 $Y2=0.072
r104 41 42 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.072 $X2=0.234 $Y2=0.072
r105 40 41 5.22839 $w=1.8e-08 $l=7.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.121
+ $Y=0.072 $X2=0.198 $Y2=0.072
r106 38 39 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.0995 $Y2=0.072
r107 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.072 $X2=0.09 $Y2=0.072
r108 36 37 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.072 $X2=0.072 $Y2=0.072
r109 34 40 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.072 $X2=0.121 $Y2=0.072
r110 34 39 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.072 $X2=0.0995 $Y2=0.072
r111 32 36 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.035
+ $Y=0.072 $X2=0.04 $Y2=0.072
r112 31 60 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.368 $Y=0.072 $X2=0.377 $Y2=0.081
r113 31 49 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.368
+ $Y=0.072 $X2=0.366 $Y2=0.072
r114 29 30 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.026
+ $Y=0.106 $X2=0.026 $Y2=0.164
r115 28 50 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.026 $Y=0.189 $X2=0.035 $Y2=0.198
r116 28 30 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.026
+ $Y=0.189 $X2=0.026 $Y2=0.164
r117 27 32 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.026 $Y=0.081 $X2=0.035 $Y2=0.072
r118 27 29 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.026
+ $Y=0.081 $X2=0.026 $Y2=0.106
r119 26 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.109 $Y=0.198
+ $X2=0.109 $Y2=0.198
r120 23 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r121 22 26 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r122 21 34 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.109 $Y=0.072
+ $X2=0.109 $Y2=0.072
r123 18 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r124 17 21 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r125 13 63 25.4545 $w=2.2e-08 $l=2.8e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.377 $Y2=0.135
r126 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r127 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r128 5 63 23.6364 $w=2.2e-08 $l=2.6e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.377 $Y2=0.135
r129 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r130 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_MAJX2_ASAP7_75T_R%7 1 6 7 13 16 17 VSS
c15 17 VSS 0.00954518f $X=0.27 $Y=0.036
c16 16 VSS 0.0247244f $X=0.27 $Y=0.036
c17 13 VSS 0.00237043f $X=0.054 $Y=0.036
c18 6 VSS 6.60818e-19 $X=0.287 $Y=0.0675
c19 1 VSS 2.69461e-19 $X=0.071 $Y=0.0675
r20 16 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r21 12 16 14.6667 $w=1.8e-08 $l=2.16e-07 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.27 $Y2=0.036
r22 12 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r23 10 17 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r24 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r25 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r26 4 13 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r27 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends

.subckt PM_MAJX2_ASAP7_75T_R%8 1 4 6 7 10 16 18 19 VSS
c17 19 VSS 0.00476966f $X=0.18 $Y=0.234
c18 18 VSS 0.00772545f $X=0.123 $Y=0.234
c19 16 VSS 0.0120511f $X=0.27 $Y=0.234
c20 10 VSS 0.00948401f $X=0.27 $Y=0.2025
c21 6 VSS 6.60818e-19 $X=0.287 $Y=0.2025
c22 4 VSS 0.00233685f $X=0.056 $Y=0.2025
c23 1 VSS 2.69461e-19 $X=0.071 $Y=0.2025
r24 18 19 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.123
+ $Y=0.234 $X2=0.18 $Y2=0.234
r25 16 19 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.18 $Y2=0.234
r26 12 18 4.68518 $w=1.8e-08 $l=6.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.123 $Y2=0.234
r27 10 16 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r28 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r29 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r30 4 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r31 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
.ends

.subckt PM_MAJX2_ASAP7_75T_R%Y 1 2 6 7 10 14 16 17 20 26 30 32 34 VSS
c20 34 VSS 0.00335843f $X=0.459 $Y=0.207
c21 32 VSS 0.00214572f $X=0.459 $Y=0.10525
c22 31 VSS 8.85605e-19 $X=0.459 $Y=0.063
c23 30 VSS 0.00202383f $X=0.459 $Y=0.1475
c24 28 VSS 8.85605e-19 $X=0.459 $Y=0.225
c25 26 VSS 0.00279029f $X=0.418 $Y=0.234
c26 25 VSS 0.00105488f $X=0.386 $Y=0.234
c27 20 VSS 0.00167554f $X=0.378 $Y=0.234
c28 18 VSS 0.00882372f $X=0.45 $Y=0.234
c29 17 VSS 0.00279029f $X=0.418 $Y=0.036
c30 16 VSS 0.00267863f $X=0.386 $Y=0.036
c31 14 VSS 0.0109023f $X=0.378 $Y=0.036
c32 11 VSS 0.00882372f $X=0.45 $Y=0.036
c33 10 VSS 0.00930355f $X=0.378 $Y=0.2025
c34 6 VSS 5.72268e-19 $X=0.395 $Y=0.2025
c35 1 VSS 5.92081e-19 $X=0.395 $Y=0.0675
r36 33 34 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.149 $X2=0.459 $Y2=0.207
r37 31 32 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.063 $X2=0.459 $Y2=0.10525
r38 30 33 0.101852 $w=1.8e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.1475 $X2=0.459 $Y2=0.149
r39 30 32 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.1475 $X2=0.459 $Y2=0.10525
r40 28 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.207
r41 27 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.063
r42 25 26 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.386
+ $Y=0.234 $X2=0.418 $Y2=0.234
r43 20 25 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.386 $Y2=0.234
r44 18 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r45 18 26 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.418 $Y2=0.234
r46 16 17 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.386
+ $Y=0.036 $X2=0.418 $Y2=0.036
r47 13 16 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.386 $Y2=0.036
r48 13 14 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r49 11 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.036 $X2=0.459 $Y2=0.045
r50 11 17 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.418 $Y2=0.036
r51 10 20 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r52 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r53 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r54 5 14 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r55 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.0675 $X2=0.378 $Y2=0.0675
r56 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.378 $Y2=0.0675
.ends

.subckt PM_MAJX2_ASAP7_75T_R%10 1 2 VSS
c3 1 VSS 0.00183233f $X=0.179 $Y=0.0675
r4 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.145 $Y2=0.0675
.ends

.subckt PM_MAJX2_ASAP7_75T_R%11 1 2 VSS
c2 1 VSS 0.00183233f $X=0.179 $Y=0.2025
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends


* END of "./MAJx2_ASAP7_75t_R.pex.sp.pex"
* 
.subckt MAJx2_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 N_6_M0_d N_A_M0_g N_7_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_10_M1_d N_B_M1_g N_6_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_C_M2_g N_10_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_7_M3_d N_C_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 VSS N_B_M4_g N_7_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_6_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_6_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_6_M7_d N_A_M7_g N_8_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M8 N_11_M8_d N_B_M8_g N_6_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M9 VDD N_C_M9_g N_11_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M10 N_8_M10_d N_C_M10_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M11 VDD N_B_M11_g N_8_M11_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M12 N_Y_M12_d N_6_M12_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M13 N_Y_M13_d N_6_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
*
* 
* .include "MAJx2_ASAP7_75t_R.pex.sp.MAJX2_ASAP7_75T_R.pxi"
* BEGIN of "./MAJx2_ASAP7_75t_R.pex.sp.MAJX2_ASAP7_75T_R.pxi"
* File: MAJx2_ASAP7_75t_R.pex.sp.MAJX2_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:37:13 2017
* 
x_PM_MAJX2_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M7_g A N_A_c_4_p N_A_c_3_p VSS
+ PM_MAJX2_ASAP7_75T_R%A
x_PM_MAJX2_ASAP7_75T_R%B N_B_M1_g N_B_c_15_n N_B_M8_g N_B_M4_g N_B_c_25_p
+ N_B_M11_g N_B_c_20_p N_B_c_16_n N_B_c_17_n N_B_c_44_p B N_B_c_28_p N_B_c_23_p
+ N_B_c_48_p N_B_c_32_p N_B_c_29_p VSS PM_MAJX2_ASAP7_75T_R%B
x_PM_MAJX2_ASAP7_75T_R%C N_C_M2_g N_C_M9_g N_C_M3_g N_C_c_63_n N_C_M10_g C
+ N_C_c_69_n N_C_c_72_n VSS PM_MAJX2_ASAP7_75T_R%C
x_PM_MAJX2_ASAP7_75T_R%6 N_6_M5_g N_6_M12_g N_6_M6_g N_6_c_90_n N_6_M13_g
+ N_6_M1_s N_6_M0_d N_6_c_106_p N_6_M8_s N_6_M7_d N_6_c_91_n N_6_c_107_p
+ N_6_c_83_n N_6_c_122_p N_6_c_105_p N_6_c_84_n N_6_c_92_n N_6_c_103_n
+ N_6_c_111_p N_6_c_94_n N_6_c_95_n N_6_c_96_n N_6_c_123_p N_6_c_97_n
+ N_6_c_112_p N_6_c_86_n N_6_c_98_n N_6_c_124_p N_6_c_99_n VSS
+ PM_MAJX2_ASAP7_75T_R%6
x_PM_MAJX2_ASAP7_75T_R%7 N_7_M0_s N_7_M4_s N_7_M3_d N_7_c_141_n N_7_c_136_n
+ N_7_c_146_n VSS PM_MAJX2_ASAP7_75T_R%7
x_PM_MAJX2_ASAP7_75T_R%8 N_8_M7_s N_8_c_159_n N_8_M11_s N_8_M10_d N_8_c_152_n
+ N_8_c_153_n N_8_c_151_n N_8_c_154_n VSS PM_MAJX2_ASAP7_75T_R%8
x_PM_MAJX2_ASAP7_75T_R%Y N_Y_M6_d N_Y_M5_d N_Y_M13_d N_Y_M12_d N_Y_c_171_n
+ N_Y_c_172_n N_Y_c_177_n N_Y_c_178_n N_Y_c_180_n N_Y_c_181_n Y N_Y_c_185_n
+ N_Y_c_168_n VSS PM_MAJX2_ASAP7_75T_R%Y
x_PM_MAJX2_ASAP7_75T_R%10 N_10_M2_s N_10_M1_d VSS PM_MAJX2_ASAP7_75T_R%10
x_PM_MAJX2_ASAP7_75T_R%11 N_11_M9_s N_11_M8_d VSS PM_MAJX2_ASAP7_75T_R%11
cc_1 N_A_M0_g N_B_M1_g 0.00355599f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_15_n 0.00118985f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A_c_3_p N_B_c_16_n 8.76278e-19 $X=0.081 $Y=0.1305 $X2=0.135 $Y2=0.135
cc_4 N_A_c_4_p N_B_c_17_n 4.37585e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.164
cc_5 N_A_M0_g N_C_M2_g 2.82885e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 A C 2.79894e-19 $X=0.082 $Y=0.116 $X2=0.135 $Y2=0.135
cc_7 A N_6_c_83_n 0.00278289f $X=0.082 $Y=0.116 $X2=0.289 $Y2=0.198
cc_8 N_A_M0_g N_6_c_84_n 2.68514e-19 $X=0.081 $Y=0.0675 $X2=0.324 $Y2=0.149
cc_9 A N_6_c_84_n 0.00120437f $X=0.082 $Y=0.116 $X2=0.324 $Y2=0.149
cc_10 N_A_M0_g N_6_c_86_n 2.68514e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_11 N_A_c_4_p N_6_c_86_n 0.00120437f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_12 N_A_M0_g N_7_c_136_n 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_13 N_A_M0_g N_8_c_151_n 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_14 N_B_M1_g N_C_M2_g 0.00341068f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_15 N_B_M4_g N_C_M2_g 2.13359e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_B_c_20_p N_C_M2_g 2.59444e-19 $X=0.18 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_17 N_B_M1_g N_C_M3_g 2.13359e-19 $X=0.135 $Y=0.0675 $X2=0.082 $Y2=0.116
cc_18 N_B_M4_g N_C_M3_g 0.00310096f $X=0.297 $Y=0.0675 $X2=0.082 $Y2=0.116
cc_19 N_B_c_23_p N_C_M3_g 2.76185e-19 $X=0.252 $Y=0.198 $X2=0.082 $Y2=0.116
cc_20 N_B_c_15_n N_C_c_63_n 0.00148337f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 N_B_c_25_p N_C_c_63_n 0.00113349f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 N_B_c_20_p N_C_c_63_n 0.00174199f $X=0.18 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 N_B_c_17_n N_C_c_63_n 4.74454e-19 $X=0.189 $Y=0.164 $X2=0.081 $Y2=0.135
cc_24 N_B_c_28_p N_C_c_63_n 4.36331e-19 $X=0.234 $Y=0.198 $X2=0.081 $Y2=0.135
cc_25 N_B_c_29_p C 6.76085e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_26 N_B_c_17_n N_C_c_69_n 8.92128e-19 $X=0.189 $Y=0.164 $X2=0 $Y2=0
cc_27 N_B_c_23_p N_C_c_69_n 0.00122099f $X=0.252 $Y=0.198 $X2=0 $Y2=0
cc_28 N_B_c_32_p N_C_c_69_n 6.40886e-19 $X=0.324 $Y=0.149 $X2=0 $Y2=0
cc_29 N_B_c_20_p N_C_c_72_n 8.92128e-19 $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_30 N_B_c_29_p N_C_c_72_n 8.67481e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_31 N_B_M4_g N_6_M5_g 0.00286002f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_32 N_B_M4_g N_6_M6_g 2.31381e-19 $X=0.297 $Y=0.0675 $X2=0.082 $Y2=0.116
cc_33 N_B_c_25_p N_6_c_90_n 9.42614e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_34 N_B_c_17_n N_6_c_91_n 4.22488e-19 $X=0.189 $Y=0.164 $X2=0 $Y2=0
cc_35 N_B_M1_g N_6_c_92_n 3.26592e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B_c_16_n N_6_c_92_n 0.00300955f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_37 N_B_c_29_p N_6_c_94_n 0.00106635f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_38 N_B_M4_g N_6_c_95_n 4.27107e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_B_c_29_p N_6_c_96_n 0.00104972f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_40 N_B_c_44_p N_6_c_97_n 6.50564e-19 $X=0.198 $Y=0.198 $X2=0 $Y2=0
cc_41 N_B_c_32_p N_6_c_98_n 0.00101322f $X=0.324 $Y=0.149 $X2=0 $Y2=0
cc_42 N_B_c_29_p N_6_c_99_n 0.00101322f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_43 N_B_M1_g N_7_c_136_n 2.64781e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.1305
cc_44 N_B_c_48_p N_8_c_152_n 0.00226064f $X=0.283 $Y=0.198 $X2=0.082 $Y2=0.116
cc_45 N_B_c_44_p N_8_c_153_n 0.00914072f $X=0.198 $Y=0.198 $X2=0.081 $Y2=0.1305
cc_46 N_B_M1_g N_8_c_154_n 4.28653e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_B_c_16_n N_8_c_154_n 0.00121846f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_48 N_B_c_29_p N_Y_c_168_n 5.35584e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_49 N_B_c_20_p N_10_M2_s 3.75655e-19 $X=0.18 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_50 N_B_c_20_p N_11_M9_s 4.4685e-19 $X=0.18 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_51 N_C_M3_g N_6_M5_g 2.13359e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_52 N_C_M2_g N_6_c_92_n 3.34646e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_53 N_C_c_63_n N_6_c_92_n 9.63103e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_54 N_C_M3_g N_6_c_103_n 2.76185e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_55 C N_6_c_103_n 0.00122099f $X=0.24 $Y=0.116 $X2=0 $Y2=0
cc_56 N_C_M2_g N_7_c_136_n 2.51542e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.1305
cc_57 N_C_M3_g N_7_c_136_n 2.38303e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.1305
cc_58 N_C_M2_g N_8_c_153_n 2.34993e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.1305
cc_59 N_C_M3_g N_8_c_153_n 2.38303e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.1305
cc_60 N_6_c_105_p N_7_M0_s 2.45503e-19 $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_61 N_6_c_106_p N_7_c_141_n 0.00376964f $X=0.108 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_62 N_6_c_107_p N_7_c_141_n 3.9292e-19 $X=0.026 $Y=0.106 $X2=0.081 $Y2=0.135
cc_63 N_6_c_105_p N_7_c_141_n 0.00242096f $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.135
cc_64 N_6_c_106_p N_7_c_136_n 0.00279121f $X=0.108 $Y=0.0675 $X2=0.081
+ $Y2=0.1305
cc_65 N_6_c_105_p N_7_c_136_n 0.0206416f $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.1305
cc_66 N_6_c_111_p N_7_c_146_n 0.00226064f $X=0.283 $Y=0.072 $X2=0 $Y2=0
cc_67 N_6_c_112_p N_8_M7_s 2.45503e-19 $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.0675
cc_68 N_6_c_91_n N_8_c_159_n 0.00376954f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_69 N_6_c_83_n N_8_c_159_n 3.31614e-19 $X=0.026 $Y=0.164 $X2=0.081 $Y2=0.135
cc_70 N_6_c_112_p N_8_c_159_n 0.00256506f $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.135
cc_71 N_6_c_91_n N_8_c_151_n 0.00279121f $X=0.108 $Y=0.2025 $X2=0 $Y2=0
cc_72 N_6_c_112_p N_8_c_151_n 0.00711303f $X=0.072 $Y=0.198 $X2=0 $Y2=0
cc_73 N_6_c_90_n N_Y_M6_d 3.80663e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_74 N_6_c_90_n N_Y_M13_d 3.80663e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.2025
cc_75 N_6_c_90_n N_Y_c_171_n 5.9618e-19 $X=0.405 $Y=0.135 $X2=0.082 $Y2=0.116
cc_76 N_6_c_90_n N_Y_c_172_n 8.00061e-19 $X=0.405 $Y=0.135 $X2=0.081 $Y2=0.135
cc_77 N_6_c_122_p N_Y_c_172_n 0.00123144f $X=0.368 $Y=0.072 $X2=0.081 $Y2=0.135
cc_78 N_6_c_123_p N_Y_c_172_n 3.88373e-19 $X=0.366 $Y=0.072 $X2=0.081 $Y2=0.135
cc_79 N_6_c_124_p N_Y_c_172_n 0.00118517f $X=0.377 $Y=0.106 $X2=0.081 $Y2=0.135
cc_80 N_6_c_99_n N_Y_c_172_n 6.41089e-19 $X=0.377 $Y=0.1205 $X2=0.081 $Y2=0.135
cc_81 N_6_c_123_p N_Y_c_177_n 0.00197206f $X=0.366 $Y=0.072 $X2=0.081 $Y2=0.1305
cc_82 N_6_M6_g N_Y_c_178_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_83 N_6_c_90_n N_Y_c_178_n 3.34995e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_84 N_6_c_98_n N_Y_c_180_n 3.75693e-19 $X=0.377 $Y=0.135 $X2=0 $Y2=0
cc_85 N_6_M6_g N_Y_c_181_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_86 N_6_c_90_n N_Y_c_181_n 3.34995e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_87 N_6_c_90_n Y 3.83961e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_88 N_6_c_99_n Y 8.61292e-19 $X=0.377 $Y=0.1205 $X2=0 $Y2=0
cc_89 N_6_c_122_p N_Y_c_185_n 8.61292e-19 $X=0.368 $Y=0.072 $X2=0 $Y2=0
cc_90 N_6_c_92_n N_10_M2_s 4.51066e-19 $X=0.198 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_91 N_7_c_141_n N_8_c_159_n 0.00154652f $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.135
cc_92 N_7_c_146_n N_8_c_152_n 0.00169333f $X=0.27 $Y=0.036 $X2=0.082 $Y2=0.116
cc_93 N_7_c_136_n N_Y_c_177_n 2.91377e-19 $X=0.27 $Y=0.036 $X2=0.081 $Y2=0.1305
cc_94 N_7_c_136_n N_10_M2_s 3.44107e-19 $X=0.27 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_95 N_8_c_153_n N_Y_c_180_n 2.91377e-19 $X=0.27 $Y=0.234 $X2=0 $Y2=0
cc_96 N_8_c_154_n N_11_M9_s 4.63074e-19 $X=0.18 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./MAJx2_ASAP7_75t_R.pex.sp.MAJX2_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: MAJx3_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:37:36 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "MAJx3_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./MAJx3_ASAP7_75t_R.pex.sp.pex"
* File: MAJx3_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:37:36 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_MAJX3_ASAP7_75T_R%A 2 5 7 10 13 16 VSS
c13 16 VSS 1.44512e-20 $X=0.081 $Y=0.1305
c14 13 VSS 3.17034e-19 $X=0.081 $Y=0.135
c15 10 VSS 3.4868e-19 $X=0.082 $Y=0.116
c16 5 VSS 0.00170659f $X=0.081 $Y=0.135
c17 2 VSS 0.0634749f $X=0.081 $Y=0.0675
r18 15 16 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.126 $X2=0.081 $Y2=0.1305
r19 13 16 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.1305
r20 10 15 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.116 $X2=0.081 $Y2=0.126
r21 5 13 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r22 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r23 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_MAJX3_ASAP7_75T_R%B 2 5 7 10 13 15 17 19 26 29 31 32 33 34 38 41 VSS
c41 41 VSS 0.00243687f $X=0.297 $Y=0.135
c42 39 VSS 0.00106497f $X=0.324 $Y=0.164
c43 38 VSS 6.22772e-20 $X=0.324 $Y=0.149
c44 37 VSS 0.00143326f $X=0.324 $Y=0.189
c45 35 VSS 4.40637e-21 $X=0.284 $Y=0.198
c46 34 VSS 5.22651e-19 $X=0.283 $Y=0.198
c47 33 VSS 8.46035e-21 $X=0.252 $Y=0.198
c48 32 VSS 0.0021192f $X=0.234 $Y=0.198
c49 29 VSS 3.26268e-19 $X=0.198 $Y=0.198
c50 28 VSS 0.00361589f $X=0.315 $Y=0.198
c51 27 VSS 6.38949e-19 $X=0.189 $Y=0.1765
c52 26 VSS 3.30052e-19 $X=0.189 $Y=0.164
c53 25 VSS 5.59921e-19 $X=0.189 $Y=0.189
c54 19 VSS 4.29576e-19 $X=0.135 $Y=0.135
c55 17 VSS 5.234e-19 $X=0.18 $Y=0.135
c56 13 VSS 0.00100977f $X=0.297 $Y=0.135
c57 10 VSS 0.0592658f $X=0.297 $Y=0.0675
c58 5 VSS 0.00119949f $X=0.135 $Y=0.135
c59 2 VSS 0.0599814f $X=0.135 $Y=0.0675
r60 41 43 1.32 $w=2.5e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.297
+ $Y=0.126 $X2=0.324 $Y2=0.126
r61 38 39 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.149 $X2=0.324 $Y2=0.164
r62 37 39 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.189 $X2=0.324 $Y2=0.164
r63 36 43 0.266695 $w=2.5e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.144 $X2=0.324 $Y2=0.126
r64 36 38 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.324
+ $Y=0.144 $X2=0.324 $Y2=0.149
r65 34 35 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.283
+ $Y=0.198 $X2=0.284 $Y2=0.198
r66 33 34 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.198 $X2=0.283 $Y2=0.198
r67 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.198 $X2=0.252 $Y2=0.198
r68 31 35 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.289
+ $Y=0.198 $X2=0.284 $Y2=0.198
r69 29 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.198 $X2=0.234 $Y2=0.198
r70 28 37 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.315 $Y=0.198 $X2=0.324 $Y2=0.189
r71 28 31 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.315
+ $Y=0.198 $X2=0.289 $Y2=0.198
r72 26 27 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.164 $X2=0.189 $Y2=0.1765
r73 25 29 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.189 $Y=0.189 $X2=0.198 $Y2=0.198
r74 25 27 0.848765 $w=1.8e-08 $l=1.25e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.189 $X2=0.189 $Y2=0.1765
r75 24 26 1.35802 $w=1.8e-08 $l=2e-08 $layer=M1 $thickness=3.6e-08 $X=0.189
+ $Y=0.144 $X2=0.189 $Y2=0.164
r76 17 24 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.18 $Y=0.135 $X2=0.189 $Y2=0.144
r77 17 19 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.135 $X2=0.135 $Y2=0.135
r78 13 41 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r79 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r80 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r81 5 19 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r82 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.2025
r83 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_MAJX3_ASAP7_75T_R%C 2 7 10 13 15 18 21 24 VSS
c28 24 VSS 1.44512e-20 $X=0.243 $Y=0.1305
c29 21 VSS 2.8151e-19 $X=0.243 $Y=0.135
c30 18 VSS 3.77468e-19 $X=0.24 $Y=0.116
c31 13 VSS 0.00942715f $X=0.243 $Y=0.135
c32 10 VSS 0.0583526f $X=0.243 $Y=0.0675
c33 2 VSS 0.0609465f $X=0.189 $Y=0.0675
r34 23 24 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.126 $X2=0.243 $Y2=0.1305
r35 21 24 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.1305
r36 18 23 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.243
+ $Y=0.116 $X2=0.243 $Y2=0.126
r37 13 21 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r38 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r39 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
r40 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.189
+ $Y=0.135 $X2=0.243 $Y2=0.135
r41 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r42 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_MAJX3_ASAP7_75T_R%6 2 7 10 15 18 21 23 25 26 29 30 31 34 37 38 39 45
+ 46 49 51 52 53 54 55 57 60 63 64 70 72 73 VSS
c55 73 VSS 2.58515e-19 $X=0.377 $Y=0.1205
c56 72 VSS 9.18711e-19 $X=0.377 $Y=0.106
c57 70 VSS 6.03793e-19 $X=0.377 $Y=0.135
c58 65 VSS 1.05074e-19 $X=0.0995 $Y=0.198
c59 64 VSS 8.46035e-21 $X=0.09 $Y=0.198
c60 63 VSS 4.41002e-19 $X=0.072 $Y=0.198
c61 62 VSS 3.80317e-19 $X=0.04 $Y=0.198
c62 60 VSS 4.23036e-19 $X=0.109 $Y=0.198
c63 58 VSS 0.00199912f $X=0.035 $Y=0.198
c64 57 VSS 1.36714e-20 $X=0.366 $Y=0.072
c65 56 VSS 0.00184044f $X=0.364 $Y=0.072
c66 55 VSS 0.0019689f $X=0.333 $Y=0.072
c67 54 VSS 0.0016201f $X=0.315 $Y=0.072
c68 53 VSS 4.40637e-21 $X=0.284 $Y=0.072
c69 52 VSS 5.22651e-19 $X=0.283 $Y=0.072
c70 51 VSS 8.46035e-21 $X=0.252 $Y=0.072
c71 50 VSS 0.00304109f $X=0.234 $Y=0.072
c72 49 VSS 2.51834e-19 $X=0.198 $Y=0.072
c73 48 VSS 2.61464e-19 $X=0.121 $Y=0.072
c74 47 VSS 1.05074e-19 $X=0.0995 $Y=0.072
c75 46 VSS 8.46035e-21 $X=0.09 $Y=0.072
c76 45 VSS 2.66799e-19 $X=0.072 $Y=0.072
c77 44 VSS 2.38309e-19 $X=0.04 $Y=0.072
c78 40 VSS 0.00206328f $X=0.035 $Y=0.072
c79 39 VSS 1.23404e-19 $X=0.368 $Y=0.072
c80 38 VSS 0.00267929f $X=0.026 $Y=0.164
c81 37 VSS 0.0010539f $X=0.026 $Y=0.106
c82 36 VSS 0.00124616f $X=0.026 $Y=0.189
c83 34 VSS 0.00350219f $X=0.108 $Y=0.2025
c84 30 VSS 6.10767e-19 $X=0.125 $Y=0.2025
c85 29 VSS 0.00357941f $X=0.108 $Y=0.0675
c86 25 VSS 6.22718e-19 $X=0.125 $Y=0.0675
c87 21 VSS 0.0137244f $X=0.459 $Y=0.135
c88 18 VSS 0.0682225f $X=0.459 $Y=0.0675
c89 10 VSS 0.0643964f $X=0.405 $Y=0.0675
c90 2 VSS 0.0617078f $X=0.351 $Y=0.0675
r91 72 73 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.377
+ $Y=0.106 $X2=0.377 $Y2=0.1205
r92 70 73 0.984568 $w=1.8e-08 $l=1.45e-08 $layer=M1 $thickness=3.6e-08 $X=0.377
+ $Y=0.135 $X2=0.377 $Y2=0.1205
r93 70 71 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.377 $Y=0.135 $X2=0.377
+ $Y2=0.135
r94 68 72 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.377
+ $Y=0.081 $X2=0.377 $Y2=0.106
r95 64 65 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.198 $X2=0.0995 $Y2=0.198
r96 63 64 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.198 $X2=0.09 $Y2=0.198
r97 62 63 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.198 $X2=0.072 $Y2=0.198
r98 60 65 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.198 $X2=0.0995 $Y2=0.198
r99 58 62 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.035
+ $Y=0.198 $X2=0.04 $Y2=0.198
r100 56 57 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.364
+ $Y=0.072 $X2=0.366 $Y2=0.072
r101 55 56 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.072 $X2=0.364 $Y2=0.072
r102 54 55 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.315
+ $Y=0.072 $X2=0.333 $Y2=0.072
r103 53 54 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.284
+ $Y=0.072 $X2=0.315 $Y2=0.072
r104 52 53 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.283
+ $Y=0.072 $X2=0.284 $Y2=0.072
r105 51 52 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.072 $X2=0.283 $Y2=0.072
r106 50 51 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.072 $X2=0.252 $Y2=0.072
r107 49 50 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.072 $X2=0.234 $Y2=0.072
r108 48 49 5.22839 $w=1.8e-08 $l=7.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.121
+ $Y=0.072 $X2=0.198 $Y2=0.072
r109 46 47 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.072 $X2=0.0995 $Y2=0.072
r110 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.072 $X2=0.09 $Y2=0.072
r111 44 45 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.04
+ $Y=0.072 $X2=0.072 $Y2=0.072
r112 42 48 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.072 $X2=0.121 $Y2=0.072
r113 42 47 0.645062 $w=1.8e-08 $l=9.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.109
+ $Y=0.072 $X2=0.0995 $Y2=0.072
r114 40 44 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.035
+ $Y=0.072 $X2=0.04 $Y2=0.072
r115 39 68 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.368 $Y=0.072 $X2=0.377 $Y2=0.081
r116 39 57 0.135802 $w=1.8e-08 $l=2e-09 $layer=M1 $thickness=3.6e-08 $X=0.368
+ $Y=0.072 $X2=0.366 $Y2=0.072
r117 37 38 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.026
+ $Y=0.106 $X2=0.026 $Y2=0.164
r118 36 58 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.026 $Y=0.189 $X2=0.035 $Y2=0.198
r119 36 38 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.026
+ $Y=0.189 $X2=0.026 $Y2=0.164
r120 35 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.026 $Y=0.081 $X2=0.035 $Y2=0.072
r121 35 37 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.026
+ $Y=0.081 $X2=0.026 $Y2=0.106
r122 34 60 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.109 $Y=0.198
+ $X2=0.109 $Y2=0.198
r123 31 34 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.108 $Y2=0.2025
r124 30 34 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.2025 $X2=0.108 $Y2=0.2025
r125 29 42 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.109 $Y=0.072
+ $X2=0.109 $Y2=0.072
r126 26 29 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.108 $Y2=0.0675
r127 25 29 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.0675 $X2=0.108 $Y2=0.0675
r128 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.135 $X2=0.459 $Y2=0.2025
r129 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.459 $Y=0.0675 $X2=0.459 $Y2=0.135
r130 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.459 $Y2=0.135
r131 13 71 25.4545 $w=2.2e-08 $l=2.8e-08 $layer=LIG $thickness=5e-08 $X=0.405
+ $Y=0.135 $X2=0.377 $Y2=0.135
r132 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r133 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r134 5 71 23.6364 $w=2.2e-08 $l=2.6e-08 $layer=LIG $thickness=5e-08 $X=0.351
+ $Y=0.135 $X2=0.377 $Y2=0.135
r135 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r136 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
.ends

.subckt PM_MAJX3_ASAP7_75T_R%7 1 6 7 13 16 17 VSS
c15 17 VSS 0.00954518f $X=0.27 $Y=0.036
c16 16 VSS 0.0245056f $X=0.27 $Y=0.036
c17 13 VSS 0.00237043f $X=0.054 $Y=0.036
c18 6 VSS 6.60818e-19 $X=0.287 $Y=0.0675
c19 1 VSS 2.69461e-19 $X=0.071 $Y=0.0675
r20 16 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r21 12 16 14.6667 $w=1.8e-08 $l=2.16e-07 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.27 $Y2=0.036
r22 12 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r23 10 17 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r24 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r25 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r26 4 13 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r27 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends

.subckt PM_MAJX3_ASAP7_75T_R%8 1 4 6 7 10 16 18 19 VSS
c17 19 VSS 0.00476966f $X=0.18 $Y=0.234
c18 18 VSS 0.00772545f $X=0.123 $Y=0.234
c19 16 VSS 0.0120511f $X=0.27 $Y=0.234
c20 10 VSS 0.00948401f $X=0.27 $Y=0.2025
c21 6 VSS 6.60818e-19 $X=0.287 $Y=0.2025
c22 4 VSS 0.00233685f $X=0.056 $Y=0.2025
c23 1 VSS 2.69461e-19 $X=0.071 $Y=0.2025
r24 18 19 3.87037 $w=1.8e-08 $l=5.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.123
+ $Y=0.234 $X2=0.18 $Y2=0.234
r25 16 19 6.11111 $w=1.8e-08 $l=9e-08 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.18 $Y2=0.234
r26 12 18 4.68518 $w=1.8e-08 $l=6.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.123 $Y2=0.234
r27 10 16 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r28 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r29 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r30 4 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r31 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
.ends

.subckt PM_MAJX3_ASAP7_75T_R%Y 1 2 6 11 12 15 16 24 26 27 30 36 40 42 44 VSS
c22 56 VSS 0.00177111f $X=0.459 $Y=0.234
c23 55 VSS 0.00177111f $X=0.459 $Y=0.036
c24 52 VSS 0.00491044f $X=0.486 $Y=0.234
c25 48 VSS 0.00614864f $X=0.486 $Y=0.036
c26 47 VSS 0.00491044f $X=0.486 $Y=0.036
c27 44 VSS 0.0022902f $X=0.459 $Y=0.207
c28 42 VSS 0.00157632f $X=0.459 $Y=0.10525
c29 41 VSS 1.4615e-20 $X=0.459 $Y=0.063
c30 40 VSS 7.28605e-19 $X=0.459 $Y=0.1475
c31 38 VSS 1.4615e-20 $X=0.459 $Y=0.225
c32 36 VSS 0.00279445f $X=0.418 $Y=0.234
c33 35 VSS 0.00105488f $X=0.386 $Y=0.234
c34 30 VSS 0.00167797f $X=0.378 $Y=0.234
c35 28 VSS 0.0052909f $X=0.45 $Y=0.234
c36 27 VSS 0.00279445f $X=0.418 $Y=0.036
c37 26 VSS 0.00268106f $X=0.386 $Y=0.036
c38 24 VSS 0.0108653f $X=0.378 $Y=0.036
c39 21 VSS 0.0052909f $X=0.45 $Y=0.036
c40 19 VSS 0.00649424f $X=0.484 $Y=0.2025
c41 15 VSS 0.00927982f $X=0.378 $Y=0.2025
c42 11 VSS 5.72268e-19 $X=0.395 $Y=0.2025
c43 9 VSS 3.45593e-19 $X=0.484 $Y=0.0675
c44 1 VSS 5.92081e-19 $X=0.395 $Y=0.0675
r45 50 56 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.459 $Y2=0.234
r46 50 52 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.234 $X2=0.486 $Y2=0.234
r47 47 48 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.036 $X2=0.486
+ $Y2=0.036
r48 45 55 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.459 $Y2=0.036
r49 45 47 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.486 $Y2=0.036
r50 43 44 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.149 $X2=0.459 $Y2=0.207
r51 41 42 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.063 $X2=0.459 $Y2=0.10525
r52 40 43 0.101852 $w=1.8e-08 $l=1.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.1475 $X2=0.459 $Y2=0.149
r53 40 42 2.86883 $w=1.8e-08 $l=4.225e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.1475 $X2=0.459 $Y2=0.10525
r54 38 56 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.234
r55 38 44 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.207
r56 37 55 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r57 37 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.063
r58 35 36 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.386
+ $Y=0.234 $X2=0.418 $Y2=0.234
r59 30 35 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.234 $X2=0.386 $Y2=0.234
r60 28 56 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.459 $Y2=0.234
r61 28 36 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.418 $Y2=0.234
r62 26 27 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.386
+ $Y=0.036 $X2=0.418 $Y2=0.036
r63 23 26 0.54321 $w=1.8e-08 $l=8e-09 $layer=M1 $thickness=3.6e-08 $X=0.378
+ $Y=0.036 $X2=0.386 $Y2=0.036
r64 23 24 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.036 $X2=0.378
+ $Y2=0.036
r65 21 55 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.459 $Y2=0.036
r66 21 27 2.17284 $w=1.8e-08 $l=3.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.418 $Y2=0.036
r67 19 52 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.234 $X2=0.486
+ $Y2=0.234
r68 16 19 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.484 $Y2=0.2025
r69 15 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.378 $Y=0.234 $X2=0.378
+ $Y2=0.234
r70 12 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.361 $Y=0.2025 $X2=0.378 $Y2=0.2025
r71 11 15 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.395 $Y=0.2025 $X2=0.378 $Y2=0.2025
r72 9 48 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.486
+ $Y=0.0675 $X2=0.486 $Y2=0.036
r73 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.469
+ $Y=0.0675 $X2=0.484 $Y2=0.0675
r74 5 24 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.378
+ $Y=0.0675 $X2=0.378 $Y2=0.036
r75 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.361
+ $Y=0.0675 $X2=0.378 $Y2=0.0675
r76 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.378 $Y2=0.0675
.ends

.subckt PM_MAJX3_ASAP7_75T_R%10 1 2 VSS
c3 1 VSS 0.00183233f $X=0.179 $Y=0.0675
r4 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.145 $Y2=0.0675
.ends

.subckt PM_MAJX3_ASAP7_75T_R%11 1 2 VSS
c2 1 VSS 0.00183233f $X=0.179 $Y=0.2025
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends


* END of "./MAJx3_ASAP7_75t_R.pex.sp.pex"
* 
.subckt MAJx3_ASAP7_75t_R  VSS VDD A B C Y
* 
* Y	Y
* C	C
* B	B
* A	A
M0 N_6_M0_d N_A_M0_g N_7_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.027
M1 N_10_M1_d N_B_M1_g N_6_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_C_M2_g N_10_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_7_M3_d N_C_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233 $Y=0.027
M4 VSS N_B_M4_g N_7_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_Y_M5_d N_6_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M6 N_Y_M6_d N_6_M6_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395 $Y=0.027
M7 N_Y_M7_d N_6_M7_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449 $Y=0.027
M8 N_6_M8_d N_A_M8_g N_8_M8_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M9 N_11_M9_d N_B_M9_g N_6_M9_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M10 VDD N_C_M10_g N_11_M10_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.162
M11 N_8_M11_d N_C_M11_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.162
M12 VDD N_B_M12_g N_8_M12_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M13 N_Y_M13_d N_6_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M14 N_Y_M14_d N_6_M14_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
M15 N_Y_M15_d N_6_M15_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.162
*
* 
* .include "MAJx3_ASAP7_75t_R.pex.sp.MAJX3_ASAP7_75T_R.pxi"
* BEGIN of "./MAJx3_ASAP7_75t_R.pex.sp.MAJX3_ASAP7_75T_R.pxi"
* File: MAJx3_ASAP7_75t_R.pex.sp.MAJX3_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:37:36 2017
* 
x_PM_MAJX3_ASAP7_75T_R%A N_A_M0_g N_A_c_2_p N_A_M8_g A N_A_c_4_p N_A_c_3_p VSS
+ PM_MAJX3_ASAP7_75T_R%A
x_PM_MAJX3_ASAP7_75T_R%B N_B_M1_g N_B_c_15_n N_B_M9_g N_B_M4_g N_B_c_25_p
+ N_B_M12_g N_B_c_20_p N_B_c_16_n N_B_c_17_n N_B_c_44_p B N_B_c_28_p N_B_c_23_p
+ N_B_c_48_p N_B_c_32_p N_B_c_29_p VSS PM_MAJX3_ASAP7_75T_R%B
x_PM_MAJX3_ASAP7_75T_R%C N_C_M2_g N_C_M10_g N_C_M3_g N_C_c_63_n N_C_M11_g C
+ N_C_c_69_n N_C_c_72_n VSS PM_MAJX3_ASAP7_75T_R%C
x_PM_MAJX3_ASAP7_75T_R%6 N_6_M5_g N_6_M13_g N_6_M6_g N_6_M14_g N_6_M7_g
+ N_6_c_90_n N_6_M15_g N_6_M1_s N_6_M0_d N_6_c_106_p N_6_M9_s N_6_M8_d
+ N_6_c_91_n N_6_c_107_p N_6_c_83_n N_6_c_122_p N_6_c_105_p N_6_c_84_n
+ N_6_c_92_n N_6_c_103_n N_6_c_111_p N_6_c_94_n N_6_c_95_n N_6_c_96_n
+ N_6_c_123_p N_6_c_97_n N_6_c_112_p N_6_c_86_n N_6_c_98_n N_6_c_124_p
+ N_6_c_99_n VSS PM_MAJX3_ASAP7_75T_R%6
x_PM_MAJX3_ASAP7_75T_R%7 N_7_M0_s N_7_M4_s N_7_M3_d N_7_c_143_n N_7_c_138_n
+ N_7_c_148_n VSS PM_MAJX3_ASAP7_75T_R%7
x_PM_MAJX3_ASAP7_75T_R%8 N_8_M8_s N_8_c_161_n N_8_M12_s N_8_M11_d N_8_c_154_n
+ N_8_c_155_n N_8_c_153_n N_8_c_156_n VSS PM_MAJX3_ASAP7_75T_R%8
x_PM_MAJX3_ASAP7_75T_R%Y N_Y_M6_d N_Y_M5_d N_Y_M7_d N_Y_M14_d N_Y_M13_d
+ N_Y_c_173_n N_Y_M15_d N_Y_c_174_n N_Y_c_179_n N_Y_c_180_n N_Y_c_182_n
+ N_Y_c_183_n Y N_Y_c_187_n N_Y_c_170_n VSS PM_MAJX3_ASAP7_75T_R%Y
x_PM_MAJX3_ASAP7_75T_R%10 N_10_M2_s N_10_M1_d VSS PM_MAJX3_ASAP7_75T_R%10
x_PM_MAJX3_ASAP7_75T_R%11 N_11_M10_s N_11_M9_d VSS PM_MAJX3_ASAP7_75T_R%11
cc_1 N_A_M0_g N_B_M1_g 0.00355599f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_c_15_n 0.00118985f $X=0.081 $Y=0.135 $X2=0.135 $Y2=0.135
cc_3 N_A_c_3_p N_B_c_16_n 8.76278e-19 $X=0.081 $Y=0.1305 $X2=0.135 $Y2=0.135
cc_4 N_A_c_4_p N_B_c_17_n 4.37585e-19 $X=0.081 $Y=0.135 $X2=0.189 $Y2=0.164
cc_5 N_A_M0_g N_C_M2_g 2.82885e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_6 A C 2.79894e-19 $X=0.082 $Y=0.116 $X2=0.135 $Y2=0.135
cc_7 A N_6_c_83_n 0.00278289f $X=0.082 $Y=0.116 $X2=0.324 $Y2=0.149
cc_8 N_A_M0_g N_6_c_84_n 2.68514e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_9 A N_6_c_84_n 0.00120437f $X=0.082 $Y=0.116 $X2=0 $Y2=0
cc_10 N_A_M0_g N_6_c_86_n 2.68514e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_11 N_A_c_4_p N_6_c_86_n 0.00120437f $X=0.081 $Y=0.135 $X2=0 $Y2=0
cc_12 N_A_M0_g N_7_c_138_n 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_13 N_A_M0_g N_8_c_153_n 2.38303e-19 $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.135
cc_14 N_B_M1_g N_C_M2_g 0.00341068f $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_15 N_B_M4_g N_C_M2_g 2.13359e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_16 N_B_c_20_p N_C_M2_g 2.59444e-19 $X=0.18 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_17 N_B_M1_g N_C_M3_g 2.13359e-19 $X=0.135 $Y=0.0675 $X2=0.082 $Y2=0.116
cc_18 N_B_M4_g N_C_M3_g 0.0030905f $X=0.297 $Y=0.0675 $X2=0.082 $Y2=0.116
cc_19 N_B_c_23_p N_C_M3_g 2.76185e-19 $X=0.252 $Y=0.198 $X2=0.082 $Y2=0.116
cc_20 N_B_c_15_n N_C_c_63_n 0.00148337f $X=0.135 $Y=0.135 $X2=0.081 $Y2=0.135
cc_21 N_B_c_25_p N_C_c_63_n 0.00113349f $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_22 N_B_c_20_p N_C_c_63_n 0.00174199f $X=0.18 $Y=0.135 $X2=0.081 $Y2=0.135
cc_23 N_B_c_17_n N_C_c_63_n 4.74454e-19 $X=0.189 $Y=0.164 $X2=0.081 $Y2=0.135
cc_24 N_B_c_28_p N_C_c_63_n 4.36331e-19 $X=0.234 $Y=0.198 $X2=0.081 $Y2=0.135
cc_25 N_B_c_29_p C 6.76085e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_26 N_B_c_17_n N_C_c_69_n 8.92128e-19 $X=0.189 $Y=0.164 $X2=0 $Y2=0
cc_27 N_B_c_23_p N_C_c_69_n 0.00122099f $X=0.252 $Y=0.198 $X2=0 $Y2=0
cc_28 N_B_c_32_p N_C_c_69_n 6.40886e-19 $X=0.324 $Y=0.149 $X2=0 $Y2=0
cc_29 N_B_c_20_p N_C_c_72_n 8.92128e-19 $X=0.18 $Y=0.135 $X2=0 $Y2=0
cc_30 N_B_c_29_p N_C_c_72_n 8.67481e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_31 N_B_M4_g N_6_M5_g 0.00288928f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_32 N_B_M4_g N_6_M6_g 2.34385e-19 $X=0.297 $Y=0.0675 $X2=0.082 $Y2=0.116
cc_33 N_B_c_25_p N_6_c_90_n 9.41786e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_34 N_B_c_17_n N_6_c_91_n 4.22488e-19 $X=0.189 $Y=0.164 $X2=0 $Y2=0
cc_35 N_B_M1_g N_6_c_92_n 3.26592e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_36 N_B_c_16_n N_6_c_92_n 0.00300955f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_37 N_B_c_29_p N_6_c_94_n 0.00106635f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_38 N_B_M4_g N_6_c_95_n 4.27107e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_39 N_B_c_29_p N_6_c_96_n 0.00104972f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_40 N_B_c_44_p N_6_c_97_n 6.50564e-19 $X=0.198 $Y=0.198 $X2=0 $Y2=0
cc_41 N_B_c_32_p N_6_c_98_n 0.00101681f $X=0.324 $Y=0.149 $X2=0 $Y2=0
cc_42 N_B_c_29_p N_6_c_99_n 0.00101681f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_43 N_B_M1_g N_7_c_138_n 2.64781e-19 $X=0.135 $Y=0.0675 $X2=0.081 $Y2=0.1305
cc_44 N_B_c_48_p N_8_c_154_n 0.00226064f $X=0.283 $Y=0.198 $X2=0.082 $Y2=0.116
cc_45 N_B_c_44_p N_8_c_155_n 0.00914072f $X=0.198 $Y=0.198 $X2=0.081 $Y2=0.1305
cc_46 N_B_M1_g N_8_c_156_n 4.28653e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_47 N_B_c_16_n N_8_c_156_n 0.00121846f $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_48 N_B_c_29_p N_Y_c_170_n 5.37696e-19 $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_49 N_B_c_20_p N_10_M2_s 3.75655e-19 $X=0.18 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_50 N_B_c_20_p N_11_M10_s 4.4685e-19 $X=0.18 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_51 N_C_M3_g N_6_M5_g 2.13359e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_52 N_C_M2_g N_6_c_92_n 3.34646e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_53 N_C_c_63_n N_6_c_92_n 9.63103e-19 $X=0.243 $Y=0.135 $X2=0 $Y2=0
cc_54 N_C_M3_g N_6_c_103_n 2.76185e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_55 C N_6_c_103_n 0.00122099f $X=0.24 $Y=0.116 $X2=0 $Y2=0
cc_56 N_C_M2_g N_7_c_138_n 2.51542e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.1305
cc_57 N_C_M3_g N_7_c_138_n 2.38303e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.1305
cc_58 N_C_M2_g N_8_c_155_n 2.34993e-19 $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.1305
cc_59 N_C_M3_g N_8_c_155_n 2.38303e-19 $X=0.243 $Y=0.0675 $X2=0.081 $Y2=0.1305
cc_60 N_6_c_105_p N_7_M0_s 2.45503e-19 $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_61 N_6_c_106_p N_7_c_143_n 0.00376964f $X=0.108 $Y=0.0675 $X2=0.081 $Y2=0.135
cc_62 N_6_c_107_p N_7_c_143_n 3.9292e-19 $X=0.026 $Y=0.106 $X2=0.081 $Y2=0.135
cc_63 N_6_c_105_p N_7_c_143_n 0.00242096f $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.135
cc_64 N_6_c_106_p N_7_c_138_n 0.00279121f $X=0.108 $Y=0.0675 $X2=0.081
+ $Y2=0.1305
cc_65 N_6_c_105_p N_7_c_138_n 0.0206416f $X=0.072 $Y=0.072 $X2=0.081 $Y2=0.1305
cc_66 N_6_c_111_p N_7_c_148_n 0.00226064f $X=0.283 $Y=0.072 $X2=0 $Y2=0
cc_67 N_6_c_112_p N_8_M8_s 2.45503e-19 $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.0675
cc_68 N_6_c_91_n N_8_c_161_n 0.00376954f $X=0.108 $Y=0.2025 $X2=0.081 $Y2=0.135
cc_69 N_6_c_83_n N_8_c_161_n 3.31614e-19 $X=0.026 $Y=0.164 $X2=0.081 $Y2=0.135
cc_70 N_6_c_112_p N_8_c_161_n 0.00256506f $X=0.072 $Y=0.198 $X2=0.081 $Y2=0.135
cc_71 N_6_c_91_n N_8_c_153_n 0.00279121f $X=0.108 $Y=0.2025 $X2=0 $Y2=0
cc_72 N_6_c_112_p N_8_c_153_n 0.00711303f $X=0.072 $Y=0.198 $X2=0 $Y2=0
cc_73 N_6_c_90_n N_Y_M6_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_74 N_6_c_90_n N_Y_M14_d 3.80663e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_75 N_6_c_90_n N_Y_c_173_n 5.9618e-19 $X=0.459 $Y=0.135 $X2=0.081 $Y2=0.126
cc_76 N_6_c_90_n N_Y_c_174_n 8.00061e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_77 N_6_c_122_p N_Y_c_174_n 0.00123144f $X=0.368 $Y=0.072 $X2=0 $Y2=0
cc_78 N_6_c_123_p N_Y_c_174_n 3.88373e-19 $X=0.366 $Y=0.072 $X2=0 $Y2=0
cc_79 N_6_c_124_p N_Y_c_174_n 0.00118517f $X=0.377 $Y=0.106 $X2=0 $Y2=0
cc_80 N_6_c_99_n N_Y_c_174_n 6.41089e-19 $X=0.377 $Y=0.1205 $X2=0 $Y2=0
cc_81 N_6_c_123_p N_Y_c_179_n 0.00197206f $X=0.366 $Y=0.072 $X2=0 $Y2=0
cc_82 N_6_M6_g N_Y_c_180_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_83 N_6_c_90_n N_Y_c_180_n 9.12592e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_84 N_6_c_98_n N_Y_c_182_n 3.75693e-19 $X=0.377 $Y=0.135 $X2=0 $Y2=0
cc_85 N_6_M6_g N_Y_c_183_n 4.59284e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_86 N_6_c_90_n N_Y_c_183_n 9.12592e-19 $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_87 N_6_c_90_n Y 0.00231288f $X=0.459 $Y=0.135 $X2=0 $Y2=0
cc_88 N_6_c_99_n Y 8.82689e-19 $X=0.377 $Y=0.1205 $X2=0 $Y2=0
cc_89 N_6_M7_g N_Y_c_187_n 3.01078e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_90 N_6_c_122_p N_Y_c_187_n 8.82689e-19 $X=0.368 $Y=0.072 $X2=0 $Y2=0
cc_91 N_6_M7_g N_Y_c_170_n 5.00993e-19 $X=0.459 $Y=0.0675 $X2=0 $Y2=0
cc_92 N_6_c_92_n N_10_M2_s 4.51066e-19 $X=0.198 $Y=0.072 $X2=0.081 $Y2=0.0675
cc_93 N_7_c_143_n N_8_c_161_n 0.00154652f $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.135
cc_94 N_7_c_148_n N_8_c_154_n 0.00169333f $X=0.27 $Y=0.036 $X2=0.082 $Y2=0.116
cc_95 N_7_c_138_n N_Y_c_179_n 3.02563e-19 $X=0.27 $Y=0.036 $X2=0 $Y2=0
cc_96 N_7_c_138_n N_10_M2_s 3.44107e-19 $X=0.27 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_97 N_8_c_155_n N_Y_c_182_n 3.02563e-19 $X=0.27 $Y=0.234 $X2=0 $Y2=0
cc_98 N_8_c_156_n N_11_M10_s 4.63074e-19 $X=0.18 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./MAJx3_ASAP7_75t_R.pex.sp.MAJX3_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: FAx1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:29:22 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "FAx1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./FAx1_ASAP7_75t_R.pex.sp.pex"
* File: FAx1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:29:22 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_FAX1_ASAP7_75T_R%A 2 7 10 13 15 18 21 23 26 29 31 33 40 44 47 53 56
+ 59 60 61 64 65 66 68 69 VSS
c83 69 VSS 0.00101542f $X=0.613 $Y=0.189
c84 68 VSS 0.00805156f $X=0.613 $Y=0.189
c85 66 VSS 0.00218299f $X=0.282 $Y=0.189
c86 65 VSS 0.00125538f $X=0.167 $Y=0.189
c87 64 VSS 3.89469e-19 $X=0.397 $Y=0.189
c88 61 VSS 4.1112e-19 $X=0.1345 $Y=0.189
c89 60 VSS 0.0023718f $X=0.128 $Y=0.189
c90 56 VSS 6.39294e-19 $X=0.073 $Y=0.189
c91 53 VSS 5.27129e-19 $X=0.621 $Y=0.167
c92 47 VSS 3.68638e-19 $X=0.621 $Y=0.135
c93 45 VSS 6.17151e-19 $X=0.621 $Y=0.18
c94 44 VSS 1.08645e-20 $X=0.405 $Y=0.1645
c95 40 VSS 9.20344e-20 $X=0.405 $Y=0.135
c96 38 VSS 6.62732e-20 $X=0.405 $Y=0.18
c97 33 VSS 0.00101019f $X=0.081 $Y=0.18
c98 29 VSS 0.00121021f $X=0.621 $Y=0.135
c99 26 VSS 0.0559973f $X=0.621 $Y=0.0675
c100 21 VSS 0.00113621f $X=0.405 $Y=0.135
c101 18 VSS 0.0594487f $X=0.405 $Y=0.0675
c102 13 VSS 0.010661f $X=0.135 $Y=0.135
c103 10 VSS 0.0624462f $X=0.135 $Y=0.0675
c104 2 VSS 0.0657415f $X=0.081 $Y=0.0675
r105 68 69 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.613 $Y=0.189 $X2=0.613
+ $Y2=0.189
r106 65 66 7.80864 $w=1.8e-08 $l=1.15e-07 $layer=M2 $thickness=3.6e-08 $X=0.167
+ $Y=0.189 $X2=0.282 $Y2=0.189
r107 63 68 14.6667 $w=1.8e-08 $l=2.16e-07 $layer=M2 $thickness=3.6e-08 $X=0.397
+ $Y=0.189 $X2=0.613 $Y2=0.189
r108 63 66 7.80864 $w=1.8e-08 $l=1.15e-07 $layer=M2 $thickness=3.6e-08 $X=0.397
+ $Y=0.189 $X2=0.282 $Y2=0.189
r109 63 64 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.397 $Y=0.189 $X2=0.397
+ $Y2=0.189
r110 60 61 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M2 $thickness=3.6e-08 $X=0.128
+ $Y=0.189 $X2=0.1345 $Y2=0.189
r111 59 65 1.76543 $w=1.8e-08 $l=2.6e-08 $layer=M2 $thickness=3.6e-08 $X=0.141
+ $Y=0.189 $X2=0.167 $Y2=0.189
r112 59 61 0.441358 $w=1.8e-08 $l=6.5e-09 $layer=M2 $thickness=3.6e-08 $X=0.141
+ $Y=0.189 $X2=0.1345 $Y2=0.189
r113 55 60 3.73457 $w=1.8e-08 $l=5.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.073
+ $Y=0.189 $X2=0.128 $Y2=0.189
r114 55 56 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.073 $Y=0.189 $X2=0.073
+ $Y2=0.189
r115 52 53 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.149 $X2=0.621 $Y2=0.167
r116 47 52 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.135 $X2=0.621 $Y2=0.149
r117 45 69 0.0717796 $w=1.8e-08 $l=1.23693e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.621 $Y=0.18 $X2=0.613 $Y2=0.189
r118 45 53 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.621
+ $Y=0.18 $X2=0.621 $Y2=0.167
r119 43 44 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.149 $X2=0.405 $Y2=0.1645
r120 40 43 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.149
r121 38 64 0.0717796 $w=1.8e-08 $l=1.23693e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.405 $Y=0.18 $X2=0.397 $Y2=0.189
r122 38 44 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.18 $X2=0.405 $Y2=0.1645
r123 33 56 0.0717796 $w=1.8e-08 $l=1.23693e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.081 $Y=0.18 $X2=0.073 $Y2=0.189
r124 33 35 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.18 $X2=0.081 $Y2=0.135
r125 29 47 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.621 $Y=0.135 $X2=0.621
+ $Y2=0.135
r126 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.135 $X2=0.621 $Y2=0.2025
r127 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.621 $Y=0.0675 $X2=0.621 $Y2=0.135
r128 21 40 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r129 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.135 $X2=0.405 $Y2=0.2025
r130 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.405 $Y=0.0675 $X2=0.405 $Y2=0.135
r131 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.135 $X2=0.135 $Y2=0.2025
r132 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08
+ $X=0.135 $Y=0.0675 $X2=0.135 $Y2=0.135
r133 5 13 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.135 $Y2=0.135
r134 5 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.135 $X2=0.081
+ $Y2=0.135
r135 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.2025
r136 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_FAX1_ASAP7_75T_R%B 2 5 7 10 15 18 21 23 26 29 31 37 41 42 44 46 47 51
+ 56 62 VSS
c64 62 VSS 0.00171728f $X=0.675 $Y=0.135
c65 56 VSS 0.0011733f $X=0.297 $Y=0.135
c66 51 VSS 5.90416e-19 $X=0.189 $Y=0.135
c67 47 VSS 0.00119634f $X=0.627 $Y=0.153
c68 46 VSS 0.00170571f $X=0.587 $Y=0.153
c69 44 VSS 0.00328347f $X=0.675 $Y=0.153
c70 42 VSS 2.11722e-19 $X=0.263 $Y=0.153
c71 41 VSS 4.68017e-19 $X=0.229 $Y=0.153
c72 29 VSS 0.00240665f $X=0.675 $Y=0.135
c73 26 VSS 0.0594173f $X=0.675 $Y=0.0675
c74 21 VSS 0.0115418f $X=0.351 $Y=0.135
c75 18 VSS 0.0628164f $X=0.351 $Y=0.0675
c76 10 VSS 0.0620159f $X=0.297 $Y=0.0675
c77 5 VSS 9.23882e-19 $X=0.189 $Y=0.135
c78 2 VSS 0.0585278f $X=0.189 $Y=0.0675
r79 46 47 2.71605 $w=1.8e-08 $l=4e-08 $layer=M2 $thickness=3.6e-08 $X=0.587
+ $Y=0.153 $X2=0.627 $Y2=0.153
r80 44 47 3.25926 $w=1.8e-08 $l=4.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.675
+ $Y=0.153 $X2=0.627 $Y2=0.153
r81 44 62 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.675 $Y=0.153 $X2=0.675
+ $Y2=0.153
r82 41 42 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.229
+ $Y=0.153 $X2=0.263 $Y2=0.153
r83 39 46 19.6914 $w=1.8e-08 $l=2.9e-07 $layer=M2 $thickness=3.6e-08 $X=0.297
+ $Y=0.153 $X2=0.587 $Y2=0.153
r84 39 42 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.297
+ $Y=0.153 $X2=0.263 $Y2=0.153
r85 39 56 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.297 $Y=0.153 $X2=0.297
+ $Y2=0.153
r86 37 41 3.25926 $w=1.8e-08 $l=4.8e-08 $layer=M2 $thickness=3.6e-08 $X=0.181
+ $Y=0.153 $X2=0.229 $Y2=0.153
r87 37 51 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.181 $Y=0.153 $X2=0.181
+ $Y2=0.153
r88 29 62 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.675 $Y=0.135 $X2=0.675
+ $Y2=0.135
r89 29 31 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.135 $X2=0.675 $Y2=0.2025
r90 26 29 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.675
+ $Y=0.0675 $X2=0.675 $Y2=0.135
r91 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r92 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r93 13 21 49.0909 $w=2.2e-08 $l=5.4e-08 $layer=LIG $thickness=5e-08 $X=0.297
+ $Y=0.135 $X2=0.351 $Y2=0.135
r94 13 56 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.297 $Y=0.135 $X2=0.297
+ $Y2=0.135
r95 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r96 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r97 5 51 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.189 $Y=0.135 $X2=0.189
+ $Y2=0.135
r98 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.135 $X2=0.189 $Y2=0.2025
r99 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.189
+ $Y=0.0675 $X2=0.189 $Y2=0.135
.ends

.subckt PM_FAX1_ASAP7_75T_R%CI 2 5 7 10 13 15 18 21 23 27 29 32 34 35 36 37 VSS
c56 37 VSS 4.89992e-19 $X=0.558 $Y=0.117
c57 36 VSS 0.00178225f $X=0.543 $Y=0.117
c58 35 VSS 0.00106902f $X=0.573 $Y=0.117
c59 34 VSS 3.37716e-19 $X=0.573 $Y=0.117
c60 32 VSS 8.05158e-19 $X=0.459 $Y=0.117
c61 27 VSS 0.0013451f $X=0.243 $Y=0.117
c62 21 VSS 0.00107594f $X=0.567 $Y=0.135
c63 18 VSS 0.0573918f $X=0.567 $Y=0.0675
c64 13 VSS 0.00113412f $X=0.459 $Y=0.135
c65 10 VSS 0.0589683f $X=0.459 $Y=0.0675
c66 5 VSS 0.00103426f $X=0.243 $Y=0.135
c67 2 VSS 0.0587152f $X=0.243 $Y=0.0675
r68 36 37 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.543
+ $Y=0.117 $X2=0.558 $Y2=0.117
r69 34 37 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.573
+ $Y=0.117 $X2=0.558 $Y2=0.117
r70 34 35 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.573 $Y=0.117 $X2=0.573
+ $Y2=0.117
r71 31 36 5.7037 $w=1.8e-08 $l=8.4e-08 $layer=M2 $thickness=3.6e-08 $X=0.459
+ $Y=0.117 $X2=0.543 $Y2=0.117
r72 31 32 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.459 $Y=0.117 $X2=0.459
+ $Y2=0.117
r73 29 31 14.6667 $w=1.8e-08 $l=2.16e-07 $layer=M2 $thickness=3.6e-08 $X=0.243
+ $Y=0.117 $X2=0.459 $Y2=0.117
r74 27 29 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.243 $Y=0.117 $X2=0.243
+ $Y2=0.117
r75 21 35 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.567 $Y=0.135 $X2=0.567
+ $Y2=0.135
r76 21 23 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.135 $X2=0.567 $Y2=0.2025
r77 18 21 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.567
+ $Y=0.0675 $X2=0.567 $Y2=0.135
r78 13 32 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.459 $Y=0.135 $X2=0.459
+ $Y2=0.135
r79 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.2025
r80 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.459
+ $Y=0.0675 $X2=0.459 $Y2=0.135
r81 5 27 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.243 $Y=0.135 $X2=0.243
+ $Y2=0.135
r82 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.135 $X2=0.243 $Y2=0.2025
r83 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.243
+ $Y=0.0675 $X2=0.243 $Y2=0.135
.ends

.subckt PM_FAX1_ASAP7_75T_R%CON 2 5 7 9 10 13 14 15 18 22 23 24 26 27 29 31 32
+ 35 37 43 46 47 48 50 62 66 67 68 VSS
c59 69 VSS 1.88705e-19 $X=0.207 $Y=0.081
c60 68 VSS 1.44512e-20 $X=0.198 $Y=0.081
c61 67 VSS 1.80896e-19 $X=0.18 $Y=0.081
c62 66 VSS 4.94527e-19 $X=0.167 $Y=0.081
c63 62 VSS 4.37092e-19 $X=0.216 $Y=0.081
c64 50 VSS 0.00684598f $X=0.529 $Y=0.081
c65 48 VSS 8.89976e-20 $X=0.229 $Y=0.081
c66 47 VSS 2.53984e-20 $X=0.167 $Y=0.081
c67 43 VSS 6.86259e-19 $X=0.142 $Y=0.081
c68 37 VSS 3.0085e-19 $X=0.513 $Y=0.135
c69 35 VSS 0.00267479f $X=0.513 $Y=0.108
c70 32 VSS 8.60543e-20 $X=0.198 $Y=0.198
c71 31 VSS 3.0894e-19 $X=0.167 $Y=0.198
c72 29 VSS 3.35608e-19 $X=0.216 $Y=0.198
c73 27 VSS 0.0010257f $X=0.142 $Y=0.198
c74 26 VSS 4.61302e-19 $X=0.133 $Y=0.178
c75 25 VSS 2.0145e-19 $X=0.133 $Y=0.167
c76 24 VSS 1.57245e-19 $X=0.133 $Y=0.162
c77 23 VSS 7.5088e-20 $X=0.133 $Y=0.144
c78 22 VSS 5.02107e-19 $X=0.133 $Y=0.121
c79 21 VSS 6.81772e-19 $X=0.133 $Y=0.108
c80 20 VSS 8.56715e-19 $X=0.133 $Y=0.189
c81 18 VSS 0.00399904f $X=0.216 $Y=0.2025
c82 14 VSS 6.36664e-19 $X=0.233 $Y=0.2025
c83 13 VSS 0.00396593f $X=0.216 $Y=0.0675
c84 9 VSS 6.47503e-19 $X=0.233 $Y=0.0675
c85 5 VSS 0.00131393f $X=0.513 $Y=0.135
c86 2 VSS 0.0599437f $X=0.513 $Y=0.0675
r87 68 69 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.198
+ $Y=0.081 $X2=0.207 $Y2=0.081
r88 67 68 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.081 $X2=0.198 $Y2=0.081
r89 66 67 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.167
+ $Y=0.081 $X2=0.18 $Y2=0.081
r90 62 69 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.081 $X2=0.207 $Y2=0.081
r91 50 51 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.529 $Y=0.081 $X2=0.529
+ $Y2=0.081
r92 47 48 4.20988 $w=1.8e-08 $l=6.2e-08 $layer=M2 $thickness=3.6e-08 $X=0.167
+ $Y=0.081 $X2=0.229 $Y2=0.081
r93 46 50 16.2284 $w=1.8e-08 $l=2.39e-07 $layer=M2 $thickness=3.6e-08 $X=0.29
+ $Y=0.081 $X2=0.529 $Y2=0.081
r94 46 48 4.14198 $w=1.8e-08 $l=6.1e-08 $layer=M2 $thickness=3.6e-08 $X=0.29
+ $Y=0.081 $X2=0.229 $Y2=0.081
r95 43 66 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.142
+ $Y=0.081 $X2=0.167 $Y2=0.081
r96 42 47 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M2 $thickness=3.6e-08 $X=0.142
+ $Y=0.081 $X2=0.167 $Y2=0.081
r97 42 43 8.97531 $a=3.24e-16 $layer=V1 $count=1 $X=0.142 $Y=0.081 $X2=0.142
+ $Y2=0.081
r98 35 51 1.32303 $w=2.85e-08 $l=3.18198e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.513 $Y=0.108 $X2=0.5235 $Y2=0.081
r99 35 37 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.513
+ $Y=0.108 $X2=0.513 $Y2=0.135
r100 31 32 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.167
+ $Y=0.198 $X2=0.198 $Y2=0.198
r101 29 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.198 $X2=0.198 $Y2=0.198
r102 27 31 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.142
+ $Y=0.198 $X2=0.167 $Y2=0.198
r103 25 26 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.133
+ $Y=0.167 $X2=0.133 $Y2=0.178
r104 24 25 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.133
+ $Y=0.162 $X2=0.133 $Y2=0.167
r105 23 24 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.133
+ $Y=0.144 $X2=0.133 $Y2=0.162
r106 22 23 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.133
+ $Y=0.121 $X2=0.133 $Y2=0.144
r107 21 22 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.133
+ $Y=0.108 $X2=0.133 $Y2=0.121
r108 20 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.133 $Y=0.189 $X2=0.142 $Y2=0.198
r109 20 26 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.133
+ $Y=0.189 $X2=0.133 $Y2=0.178
r110 19 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.133 $Y=0.09 $X2=0.142 $Y2=0.081
r111 19 21 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.133
+ $Y=0.09 $X2=0.133 $Y2=0.108
r112 18 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.198
+ $X2=0.216 $Y2=0.198
r113 15 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.2025 $X2=0.216 $Y2=0.2025
r114 14 18 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.2025 $X2=0.216 $Y2=0.2025
r115 13 62 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.216 $Y=0.081
+ $X2=0.216 $Y2=0.081
r116 10 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.199 $Y=0.0675 $X2=0.216 $Y2=0.0675
r117 9 13 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.233 $Y=0.0675 $X2=0.216 $Y2=0.0675
r118 5 37 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.513 $Y=0.135 $X2=0.513
+ $Y2=0.135
r119 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.135 $X2=0.513 $Y2=0.2025
r120 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.513
+ $Y=0.0675 $X2=0.513 $Y2=0.135
.ends

.subckt PM_FAX1_ASAP7_75T_R%7 1 6 7 13 16 17 20 21 VSS
c17 21 VSS 0.00588628f $X=0.124 $Y=0.036
c18 20 VSS 0.00142972f $X=0.09 $Y=0.036
c19 19 VSS 0.00127429f $X=0.072 $Y=0.036
c20 18 VSS 0.00320092f $X=0.059 $Y=0.036
c21 17 VSS 0.00567313f $X=0.27 $Y=0.036
c22 16 VSS 0.0137438f $X=0.27 $Y=0.036
c23 13 VSS 0.00565136f $X=0.054 $Y=0.036
c24 6 VSS 6.59235e-19 $X=0.287 $Y=0.0675
c25 1 VSS 2.69461e-19 $X=0.071 $Y=0.0675
r26 20 21 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.036 $X2=0.124 $Y2=0.036
r27 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.072
+ $Y=0.036 $X2=0.09 $Y2=0.036
r28 18 19 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.059
+ $Y=0.036 $X2=0.072 $Y2=0.036
r29 16 21 9.91358 $w=1.8e-08 $l=1.46e-07 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.036 $X2=0.124 $Y2=0.036
r30 16 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.036 $X2=0.27
+ $Y2=0.036
r31 12 18 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.059 $Y2=0.036
r32 12 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r33 10 17 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.27
+ $Y=0.0675 $X2=0.27 $Y2=0.036
r34 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.0675 $X2=0.27 $Y2=0.0675
r35 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.0675 $X2=0.27 $Y2=0.0675
r36 4 13 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.054
+ $Y=0.0675 $X2=0.054 $Y2=0.036
r37 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.0675 $X2=0.056 $Y2=0.0675
.ends

.subckt PM_FAX1_ASAP7_75T_R%8 1 4 6 7 10 16 19 20 21 22 23 25 VSS
c23 25 VSS 3.80702e-19 $X=0.2665 $Y=0.234
c24 24 VSS 0.00100634f $X=0.263 $Y=0.234
c25 23 VSS 0.00146362f $X=0.252 $Y=0.234
c26 22 VSS 3.67066e-19 $X=0.234 $Y=0.234
c27 21 VSS 0.00852672f $X=0.23 $Y=0.234
c28 20 VSS 0.00583598f $X=0.124 $Y=0.234
c29 19 VSS 0.00248313f $X=0.09 $Y=0.234
c30 18 VSS 0.00318704f $X=0.059 $Y=0.234
c31 16 VSS 0.00236354f $X=0.27 $Y=0.234
c32 10 VSS 0.00618666f $X=0.27 $Y=0.2025
c33 6 VSS 6.49491e-19 $X=0.287 $Y=0.2025
c34 4 VSS 0.00619865f $X=0.056 $Y=0.2025
c35 1 VSS 3.0531e-19 $X=0.071 $Y=0.2025
r36 24 25 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.263
+ $Y=0.234 $X2=0.2665 $Y2=0.234
r37 23 24 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.252
+ $Y=0.234 $X2=0.263 $Y2=0.234
r38 22 23 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.234
+ $Y=0.234 $X2=0.252 $Y2=0.234
r39 21 22 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.23
+ $Y=0.234 $X2=0.234 $Y2=0.234
r40 20 21 7.19753 $w=1.8e-08 $l=1.06e-07 $layer=M1 $thickness=3.6e-08 $X=0.124
+ $Y=0.234 $X2=0.23 $Y2=0.234
r41 19 20 2.30864 $w=1.8e-08 $l=3.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.09
+ $Y=0.234 $X2=0.124 $Y2=0.234
r42 18 19 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.059
+ $Y=0.234 $X2=0.09 $Y2=0.234
r43 16 25 0.237654 $w=1.8e-08 $l=3.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.2665 $Y2=0.234
r44 12 18 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.059 $Y2=0.234
r45 10 16 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r46 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.253 $Y=0.2025 $X2=0.27 $Y2=0.2025
r47 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.287 $Y=0.2025 $X2=0.27 $Y2=0.2025
r48 4 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r49 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.071
+ $Y=0.2025 $X2=0.056 $Y2=0.2025
.ends

.subckt PM_FAX1_ASAP7_75T_R%SN 1 2 5 6 7 10 14 17 18 20 21 22 23 24 28 29 31 32
+ 33 35 36 37 38 39 40 43 46 VSS
c46 49 VSS 2.602e-19 $X=0.486 $Y=0.054
c47 46 VSS 0.00203263f $X=0.486 $Y=0.036
c48 43 VSS 6.3239e-20 $X=0.486 $Y=0.198
c49 40 VSS 0.00164171f $X=0.468 $Y=0.234
c50 39 VSS 0.003286f $X=0.45 $Y=0.234
c51 38 VSS 0.00261714f $X=0.414 $Y=0.234
c52 37 VSS 0.00385212f $X=0.383 $Y=0.234
c53 36 VSS 0.0038898f $X=0.342 $Y=0.234
c54 35 VSS 0.00279621f $X=0.477 $Y=0.234
c55 34 VSS 4.60225e-19 $X=0.4725 $Y=0.036
c56 33 VSS 0.00145884f $X=0.468 $Y=0.036
c57 32 VSS 0.00332824f $X=0.45 $Y=0.036
c58 31 VSS 0.00142972f $X=0.414 $Y=0.036
c59 30 VSS 0.00139575f $X=0.396 $Y=0.036
c60 29 VSS 0.00377613f $X=0.383 $Y=0.036
c61 28 VSS 0.0038898f $X=0.342 $Y=0.036
c62 27 VSS 3.27473e-19 $X=0.477 $Y=0.036
c63 26 VSS 3.72558e-19 $X=0.333 $Y=0.211
c64 25 VSS 4.67328e-19 $X=0.333 $Y=0.207
c65 24 VSS 5.52181e-19 $X=0.333 $Y=0.198
c66 23 VSS 5.85069e-19 $X=0.333 $Y=0.189
c67 22 VSS 0.00113024f $X=0.333 $Y=0.18
c68 21 VSS 6.94044e-19 $X=0.333 $Y=0.167
c69 20 VSS 5.46546e-19 $X=0.333 $Y=0.121
c70 19 VSS 5.69494e-19 $X=0.333 $Y=0.108
c71 18 VSS 0.00108154f $X=0.333 $Y=0.103
c72 17 VSS 4.34944e-19 $X=0.333 $Y=0.09
c73 16 VSS 4.05732e-19 $X=0.333 $Y=0.072
c74 15 VSS 0.00206372f $X=0.333 $Y=0.068
c75 14 VSS 0.00125738f $X=0.334 $Y=0.215
c76 10 VSS 0.0028356f $X=0.486 $Y=0.2025
c77 6 VSS 5.945e-19 $X=0.503 $Y=0.2025
c78 5 VSS 0.00282385f $X=0.486 $Y=0.0675
c79 1 VSS 5.81027e-19 $X=0.503 $Y=0.0675
r80 51 52 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.045 $X2=0.486 $Y2=0.0495
r81 49 52 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.054 $X2=0.486 $Y2=0.0495
r82 46 51 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.036 $X2=0.486 $Y2=0.045
r83 41 43 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.486
+ $Y=0.225 $X2=0.486 $Y2=0.198
r84 39 40 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.468 $Y2=0.234
r85 38 39 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.45 $Y2=0.234
r86 37 38 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.383
+ $Y=0.234 $X2=0.414 $Y2=0.234
r87 36 37 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.234 $X2=0.383 $Y2=0.234
r88 35 41 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.477 $Y=0.234 $X2=0.486 $Y2=0.225
r89 35 40 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.477
+ $Y=0.234 $X2=0.468 $Y2=0.234
r90 33 34 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.468
+ $Y=0.036 $X2=0.4725 $Y2=0.036
r91 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.468 $Y2=0.036
r92 31 32 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.036 $X2=0.45 $Y2=0.036
r93 30 31 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.036 $X2=0.414 $Y2=0.036
r94 29 30 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.383
+ $Y=0.036 $X2=0.396 $Y2=0.036
r95 28 29 2.78395 $w=1.8e-08 $l=4.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.036 $X2=0.383 $Y2=0.036
r96 27 46 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.477
+ $Y=0.036 $X2=0.486 $Y2=0.036
r97 27 34 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.477
+ $Y=0.036 $X2=0.4725 $Y2=0.036
r98 25 26 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.207 $X2=0.333 $Y2=0.211
r99 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.198 $X2=0.333 $Y2=0.207
r100 23 24 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.189 $X2=0.333 $Y2=0.198
r101 22 23 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.18 $X2=0.333 $Y2=0.189
r102 21 22 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.167 $X2=0.333 $Y2=0.18
r103 20 21 3.12346 $w=1.8e-08 $l=4.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.121 $X2=0.333 $Y2=0.167
r104 19 20 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.108 $X2=0.333 $Y2=0.121
r105 18 19 0.339506 $w=1.8e-08 $l=5e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.103 $X2=0.333 $Y2=0.108
r106 17 18 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.09 $X2=0.333 $Y2=0.103
r107 16 17 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.072 $X2=0.333 $Y2=0.09
r108 15 16 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.068 $X2=0.333 $Y2=0.072
r109 14 26 0.271605 $w=1.8e-08 $l=4e-09 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.215 $X2=0.333 $Y2=0.211
r110 12 36 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.333 $Y=0.225 $X2=0.342 $Y2=0.234
r111 12 14 0.679012 $w=1.8e-08 $l=1e-08 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.225 $X2=0.333 $Y2=0.215
r112 11 28 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.333 $Y=0.045 $X2=0.342 $Y2=0.036
r113 11 15 1.56173 $w=1.8e-08 $l=2.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.333
+ $Y=0.045 $X2=0.333 $Y2=0.068
r114 10 43 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.198
+ $X2=0.486 $Y2=0.198
r115 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.2025 $X2=0.486 $Y2=0.2025
r116 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.2025 $X2=0.486 $Y2=0.2025
r117 5 49 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.486 $Y=0.054 $X2=0.486
+ $Y2=0.054
r118 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.469 $Y=0.0675 $X2=0.486 $Y2=0.0675
r119 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.503 $Y=0.0675 $X2=0.486 $Y2=0.0675
.ends

.subckt PM_FAX1_ASAP7_75T_R%10 1 2 6 7 13 16 17 18 20 21 23 VSS
c16 23 VSS 0.00147038f $X=0.63 $Y=0.036
c17 22 VSS 0.0021772f $X=0.612 $Y=0.036
c18 21 VSS 0.00206834f $X=0.599 $Y=0.036
c19 20 VSS 0.00310894f $X=0.587 $Y=0.036
c20 19 VSS 0.00156875f $X=0.558 $Y=0.036
c21 18 VSS 0.00179868f $X=0.543 $Y=0.036
c22 17 VSS 0.00854116f $X=0.648 $Y=0.036
c23 16 VSS 0.0041274f $X=0.648 $Y=0.036
c24 13 VSS 0.00645597f $X=0.54 $Y=0.036
c25 6 VSS 5.72268e-19 $X=0.665 $Y=0.0675
c26 1 VSS 6.15477e-19 $X=0.557 $Y=0.0675
r27 22 23 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.612
+ $Y=0.036 $X2=0.63 $Y2=0.036
r28 21 22 0.882716 $w=1.8e-08 $l=1.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.599
+ $Y=0.036 $X2=0.612 $Y2=0.036
r29 20 21 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.587
+ $Y=0.036 $X2=0.599 $Y2=0.036
r30 19 20 1.96914 $w=1.8e-08 $l=2.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.036 $X2=0.587 $Y2=0.036
r31 18 19 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.543
+ $Y=0.036 $X2=0.558 $Y2=0.036
r32 16 23 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.036 $X2=0.63 $Y2=0.036
r33 16 17 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.036 $X2=0.648
+ $Y2=0.036
r34 12 18 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.036 $X2=0.543 $Y2=0.036
r35 12 13 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.036 $X2=0.54
+ $Y2=0.036
r36 10 17 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.648
+ $Y=0.0675 $X2=0.648 $Y2=0.036
r37 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.0675 $X2=0.648 $Y2=0.0675
r38 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.0675 $X2=0.648 $Y2=0.0675
r39 5 13 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.54
+ $Y=0.0675 $X2=0.54 $Y2=0.036
r40 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.523
+ $Y=0.0675 $X2=0.54 $Y2=0.0675
r41 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=N_src_drn $thickness=1e-09 $X=0.557
+ $Y=0.0675 $X2=0.54 $Y2=0.0675
.ends

.subckt PM_FAX1_ASAP7_75T_R%11 1 2 5 6 7 10 12 18 22 25 VSS
c15 25 VSS 0.00345866f $X=0.63 $Y=0.234
c16 24 VSS 0.0019857f $X=0.599 $Y=0.234
c17 23 VSS 0.00181262f $X=0.587 $Y=0.234
c18 22 VSS 0.00142296f $X=0.576 $Y=0.234
c19 21 VSS 0.00135758f $X=0.558 $Y=0.234
c20 20 VSS 5.29738e-19 $X=0.543 $Y=0.234
c21 18 VSS 0.00411198f $X=0.648 $Y=0.234
c22 12 VSS 0.00148269f $X=0.54 $Y=0.234
c23 10 VSS 0.00988919f $X=0.648 $Y=0.2025
c24 6 VSS 5.72268e-19 $X=0.665 $Y=0.2025
c25 5 VSS 0.00636683f $X=0.54 $Y=0.2025
c26 1 VSS 5.72268e-19 $X=0.557 $Y=0.2025
r27 24 25 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.599
+ $Y=0.234 $X2=0.63 $Y2=0.234
r28 23 24 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.587
+ $Y=0.234 $X2=0.599 $Y2=0.234
r29 22 23 0.746914 $w=1.8e-08 $l=1.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.576
+ $Y=0.234 $X2=0.587 $Y2=0.234
r30 21 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.558
+ $Y=0.234 $X2=0.576 $Y2=0.234
r31 20 21 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.543
+ $Y=0.234 $X2=0.558 $Y2=0.234
r32 18 25 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.648
+ $Y=0.234 $X2=0.63 $Y2=0.234
r33 12 20 0.203704 $w=1.8e-08 $l=3e-09 $layer=M1 $thickness=3.6e-08 $X=0.54
+ $Y=0.234 $X2=0.543 $Y2=0.234
r34 10 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.648 $Y=0.234 $X2=0.648
+ $Y2=0.234
r35 7 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.631 $Y=0.2025 $X2=0.648 $Y2=0.2025
r36 6 10 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.665 $Y=0.2025 $X2=0.648 $Y2=0.2025
r37 5 12 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.54 $Y=0.234 $X2=0.54
+ $Y2=0.234
r38 2 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.523
+ $Y=0.2025 $X2=0.54 $Y2=0.2025
r39 1 5 8.39506 $w=8.1e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09 $X=0.557
+ $Y=0.2025 $X2=0.54 $Y2=0.2025
.ends

.subckt PM_FAX1_ASAP7_75T_R%12 1 2 VSS
c1 1 VSS 0.00226413f $X=0.179 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.0675 $X2=0.145 $Y2=0.0675
.ends

.subckt PM_FAX1_ASAP7_75T_R%13 1 2 VSS
c1 1 VSS 0.001961f $X=0.395 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.0675 $X2=0.361 $Y2=0.0675
.ends

.subckt PM_FAX1_ASAP7_75T_R%14 1 2 VSS
c1 1 VSS 0.00183233f $X=0.449 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.449
+ $Y=0.0675 $X2=0.415 $Y2=0.0675
.ends

.subckt PM_FAX1_ASAP7_75T_R%15 1 2 VSS
c1 1 VSS 0.00223579f $X=0.179 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.179
+ $Y=0.2025 $X2=0.145 $Y2=0.2025
.ends

.subckt PM_FAX1_ASAP7_75T_R%16 1 2 VSS
c2 1 VSS 0.00191352f $X=0.395 $Y=0.2025
r3 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.395
+ $Y=0.2025 $X2=0.361 $Y2=0.2025
.ends

.subckt PM_FAX1_ASAP7_75T_R%17 1 2 VSS
c1 1 VSS 0.00183233f $X=0.449 $Y=0.2025
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=P_src_drn $thickness=1e-09 $X=0.449
+ $Y=0.2025 $X2=0.415 $Y2=0.2025
.ends


* END of "./FAx1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt FAx1_ASAP7_75t_R  VSS VDD A B CI CON SN
* 
* SN	SN
* CON	CON
* CI	CI
* B	B
* A	A
M0 VSS N_A_M0_g N_7_M0_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_12_M1_d N_A_M1_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 N_CON_M2_d N_B_M2_g N_12_M2_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.179
+ $Y=0.027
M3 N_7_M3_d N_CI_M3_g N_CON_M3_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.233
+ $Y=0.027
M4 VSS N_B_M4_g N_7_M4_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M5 N_13_M5_d N_B_M5_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.027
M6 N_14_M6_d N_A_M6_g N_13_M6_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M7 N_SN_M7_d N_CI_M7_g N_14_M7_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.449
+ $Y=0.027
M8 N_10_M8_d N_CON_M8_g N_SN_M8_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.503
+ $Y=0.027
M9 VSS N_CI_M9_g N_10_M9_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.027
M10 N_10_M10_d N_A_M10_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.027
M11 VSS N_B_M11_g N_10_M11_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.027
M12 VDD N_A_M12_g N_8_M12_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071
+ $Y=0.162
M13 N_15_M13_d N_A_M13_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.162
M14 N_CON_M14_d N_B_M14_g N_15_M14_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.179 $Y=0.162
M15 N_8_M15_d N_CI_M15_g N_CON_M15_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.233 $Y=0.162
M16 VDD N_B_M16_g N_8_M16_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M17 N_16_M17_d N_B_M17_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341
+ $Y=0.162
M18 N_17_M18_d N_A_M18_g N_16_M18_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.395 $Y=0.162
M19 N_SN_M19_d N_CI_M19_g N_17_M19_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.449 $Y=0.162
M20 N_11_M20_d N_CON_M20_g N_SN_M20_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3
+ $X=0.503 $Y=0.162
M21 VDD N_CI_M21_g N_11_M21_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.557
+ $Y=0.162
M22 N_11_M22_d N_A_M22_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.611
+ $Y=0.162
M23 VDD N_B_M23_g N_11_M23_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.665
+ $Y=0.162
*
* 
* .include "FAx1_ASAP7_75t_R.pex.sp.FAX1_ASAP7_75T_R.pxi"
* BEGIN of "./FAx1_ASAP7_75t_R.pex.sp.FAX1_ASAP7_75T_R.pxi"
* File: FAx1_ASAP7_75t_R.pex.sp.FAX1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:29:22 2017
* 
x_PM_FAX1_ASAP7_75T_R%A N_A_M0_g N_A_M12_g N_A_M1_g N_A_c_3_p N_A_M13_g N_A_M6_g
+ N_A_c_6_p N_A_M18_g N_A_M10_g N_A_c_9_p N_A_M22_g N_A_c_34_p N_A_c_11_p
+ N_A_c_12_p N_A_c_15_p N_A_c_16_p N_A_c_36_p A N_A_c_47_p N_A_c_42_p N_A_c_13_p
+ N_A_c_39_p N_A_c_10_p N_A_c_7_p N_A_c_17_p VSS PM_FAX1_ASAP7_75T_R%A
x_PM_FAX1_ASAP7_75T_R%B N_B_M2_g N_B_c_86_n N_B_M14_g N_B_M4_g N_B_M16_g
+ N_B_M5_g N_B_c_89_n N_B_M17_g N_B_M11_g N_B_c_92_n N_B_M23_g B N_B_c_93_n
+ N_B_c_111_p N_B_c_143_p N_B_c_94_n N_B_c_98_n N_B_c_101_n N_B_c_102_n
+ N_B_c_103_n VSS PM_FAX1_ASAP7_75T_R%B
x_PM_FAX1_ASAP7_75T_R%CI N_CI_M3_g N_CI_c_161_n N_CI_M15_g N_CI_M7_g
+ N_CI_c_150_n N_CI_M19_g N_CI_M9_g N_CI_c_152_n N_CI_M21_g N_CI_c_165_n CI
+ N_CI_c_153_n N_CI_c_200_p N_CI_c_154_n N_CI_c_155_n N_CI_c_157_n VSS
+ PM_FAX1_ASAP7_75T_R%CI
x_PM_FAX1_ASAP7_75T_R%CON N_CON_M8_g N_CON_c_231_n N_CON_M20_g N_CON_M3_s
+ N_CON_M2_d N_CON_c_245_p N_CON_M15_s N_CON_M14_d N_CON_c_251_p N_CON_c_233_n
+ N_CON_c_206_n N_CON_c_208_n N_CON_c_209_n N_CON_c_210_n N_CON_c_211_n
+ N_CON_c_212_n N_CON_c_213_n N_CON_c_234_n N_CON_c_221_n N_CON_c_214_n CON
+ N_CON_c_215_n N_CON_c_222_n N_CON_c_224_n N_CON_c_242_n N_CON_c_248_p
+ N_CON_c_226_n N_CON_c_227_n VSS PM_FAX1_ASAP7_75T_R%CON
x_PM_FAX1_ASAP7_75T_R%7 N_7_M0_s N_7_M4_s N_7_M3_d N_7_c_276_p N_7_c_263_n
+ N_7_c_274_n N_7_c_264_n N_7_c_266_n VSS PM_FAX1_ASAP7_75T_R%7
x_PM_FAX1_ASAP7_75T_R%8 N_8_M12_s N_8_c_280_n N_8_M16_s N_8_M15_d N_8_c_283_n
+ N_8_c_301_p N_8_c_284_n N_8_c_287_n N_8_c_289_n N_8_c_290_n N_8_c_293_n
+ N_8_c_291_n VSS PM_FAX1_ASAP7_75T_R%8
x_PM_FAX1_ASAP7_75T_R%SN N_SN_M8_s N_SN_M7_d N_SN_c_332_n N_SN_M20_s N_SN_M19_d
+ N_SN_c_303_n SN N_SN_c_318_n N_SN_c_319_n N_SN_c_320_n N_SN_c_304_n
+ N_SN_c_305_n N_SN_c_306_n N_SN_c_308_n N_SN_c_337_n N_SN_c_325_n N_SN_c_309_n
+ N_SN_c_346_p N_SN_c_329_n N_SN_c_344_p N_SN_c_338_n N_SN_c_311_n N_SN_c_312_n
+ N_SN_c_315_n N_SN_c_331_n N_SN_c_316_n N_SN_c_341_p VSS PM_FAX1_ASAP7_75T_R%SN
x_PM_FAX1_ASAP7_75T_R%10 N_10_M9_s N_10_M8_d N_10_M11_s N_10_M10_d N_10_c_357_n
+ N_10_c_351_n N_10_c_352_n N_10_c_358_n N_10_c_354_n N_10_c_353_n N_10_c_349_n
+ VSS PM_FAX1_ASAP7_75T_R%10
x_PM_FAX1_ASAP7_75T_R%11 N_11_M21_s N_11_M20_d N_11_c_365_n N_11_M23_s
+ N_11_M22_d N_11_c_366_n N_11_c_367_n N_11_c_372_n N_11_c_373_n N_11_c_368_n
+ VSS PM_FAX1_ASAP7_75T_R%11
x_PM_FAX1_ASAP7_75T_R%12 N_12_M2_s N_12_M1_d VSS PM_FAX1_ASAP7_75T_R%12
x_PM_FAX1_ASAP7_75T_R%13 N_13_M6_s N_13_M5_d VSS PM_FAX1_ASAP7_75T_R%13
x_PM_FAX1_ASAP7_75T_R%14 N_14_M7_s N_14_M6_d VSS PM_FAX1_ASAP7_75T_R%14
x_PM_FAX1_ASAP7_75T_R%15 N_15_M14_s N_15_M13_d VSS PM_FAX1_ASAP7_75T_R%15
x_PM_FAX1_ASAP7_75T_R%16 N_16_M18_s N_16_M17_d VSS PM_FAX1_ASAP7_75T_R%16
x_PM_FAX1_ASAP7_75T_R%17 N_17_M19_s N_17_M18_d VSS PM_FAX1_ASAP7_75T_R%17
cc_1 N_A_M0_g N_B_M2_g 2.13359e-19 $X=0.081 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_2 N_A_M1_g N_B_M2_g 0.00341068f $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_3 N_A_c_3_p N_B_c_86_n 9.57863e-19 $X=0.135 $Y=0.135 $X2=0.189 $Y2=0.135
cc_4 N_A_M6_g N_B_M4_g 2.13359e-19 $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_5 N_A_M6_g N_B_M5_g 0.00341068f $X=0.405 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_6 N_A_c_6_p N_B_c_89_n 0.00119274f $X=0.405 $Y=0.135 $X2=0.351 $Y2=0.135
cc_7 N_A_c_7_p N_B_c_89_n 2.21426e-19 $X=0.613 $Y=0.189 $X2=0.351 $Y2=0.135
cc_8 N_A_M10_g N_B_M11_g 0.00316373f $X=0.621 $Y=0.0675 $X2=0.675 $Y2=0.0675
cc_9 N_A_c_9_p N_B_c_92_n 0.00101372f $X=0.621 $Y=0.135 $X2=0.675 $Y2=0.135
cc_10 N_A_c_10_p N_B_c_93_n 0.0189567f $X=0.282 $Y=0.189 $X2=0.229 $Y2=0.153
cc_11 N_A_c_11_p N_B_c_94_n 3.42042e-19 $X=0.405 $Y=0.135 $X2=0.587 $Y2=0.153
cc_12 N_A_c_12_p N_B_c_94_n 8.42075e-19 $X=0.405 $Y=0.1645 $X2=0.587 $Y2=0.153
cc_13 N_A_c_13_p N_B_c_94_n 2.46239e-19 $X=0.397 $Y=0.189 $X2=0.587 $Y2=0.153
cc_14 N_A_c_7_p N_B_c_94_n 0.0189567f $X=0.613 $Y=0.189 $X2=0.587 $Y2=0.153
cc_15 N_A_c_15_p N_B_c_98_n 4.12584e-19 $X=0.621 $Y=0.135 $X2=0.627 $Y2=0.153
cc_16 N_A_c_16_p N_B_c_98_n 5.8113e-19 $X=0.621 $Y=0.167 $X2=0.627 $Y2=0.153
cc_17 N_A_c_17_p N_B_c_98_n 2.46239e-19 $X=0.613 $Y=0.189 $X2=0.627 $Y2=0.153
cc_18 N_A_c_10_p N_B_c_101_n 3.67071e-19 $X=0.282 $Y=0.189 $X2=0.189 $Y2=0.135
cc_19 N_A_c_7_p N_B_c_102_n 2.46239e-19 $X=0.613 $Y=0.189 $X2=0.297 $Y2=0.135
cc_20 N_A_c_15_p N_B_c_103_n 0.00204558f $X=0.621 $Y=0.135 $X2=0.675 $Y2=0.135
cc_21 N_A_M1_g N_CI_M3_g 2.82885e-19 $X=0.135 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_22 N_A_M6_g N_CI_M7_g 0.00355599f $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_23 N_A_c_6_p N_CI_c_150_n 0.00105615f $X=0.405 $Y=0.135 $X2=0.297 $Y2=0.135
cc_24 N_A_M10_g N_CI_M9_g 0.00268443f $X=0.621 $Y=0.0675 $X2=0.351 $Y2=0.0675
cc_25 N_A_c_9_p N_CI_c_152_n 9.85642e-19 $X=0.621 $Y=0.135 $X2=0.351 $Y2=0.135
cc_26 N_A_c_11_p N_CI_c_153_n 0.00130629f $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_27 N_A_c_15_p N_CI_c_154_n 0.00118368f $X=0.621 $Y=0.135 $X2=0.181 $Y2=0.153
cc_28 N_A_c_11_p N_CI_c_155_n 5.49899e-19 $X=0.405 $Y=0.135 $X2=0 $Y2=0
cc_29 N_A_c_10_p N_CI_c_155_n 8.21999e-19 $X=0.282 $Y=0.189 $X2=0 $Y2=0
cc_30 N_A_c_7_p N_CI_c_157_n 8.21999e-19 $X=0.613 $Y=0.189 $X2=0.187 $Y2=0.153
cc_31 N_A_M6_g N_CON_M8_g 2.94371e-19 $X=0.405 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_32 N_A_M10_g N_CON_M8_g 2.13359e-19 $X=0.621 $Y=0.0675 $X2=0.189 $Y2=0.0675
cc_33 N_A_c_3_p N_CON_c_206_n 0.00173267f $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.2025
cc_34 N_A_c_34_p N_CON_c_206_n 0.00182504f $X=0.081 $Y=0.18 $X2=0.351 $Y2=0.2025
cc_35 N_A_c_3_p N_CON_c_208_n 4.53041e-19 $X=0.135 $Y=0.135 $X2=0 $Y2=0
cc_36 N_A_c_36_p N_CON_c_209_n 0.00182504f $X=0.073 $Y=0.189 $X2=0.675
+ $Y2=0.0675
cc_37 N_A_M1_g N_CON_c_210_n 2.0706e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_38 N_A_c_10_p N_CON_c_211_n 9.26735e-19 $X=0.282 $Y=0.189 $X2=0.675 $Y2=0.135
cc_39 N_A_c_39_p N_CON_c_212_n 6.49221e-19 $X=0.167 $Y=0.189 $X2=0.675
+ $Y2=0.2025
cc_40 N_A_c_10_p N_CON_c_213_n 7.75952e-19 $X=0.282 $Y=0.189 $X2=0 $Y2=0
cc_41 N_A_M1_g N_CON_c_214_n 2.79555e-19 $X=0.135 $Y=0.0675 $X2=0.675 $Y2=0.153
cc_42 N_A_c_42_p N_CON_c_215_n 9.27014e-19 $X=0.1345 $Y=0.189 $X2=0.627
+ $Y2=0.153
cc_43 N_A_M1_g N_7_c_263_n 2.97734e-19 $X=0.135 $Y=0.0675 $X2=0 $Y2=0
cc_44 N_A_M0_g N_7_c_264_n 3.65337e-19 $X=0.081 $Y=0.0675 $X2=0.351 $Y2=0.135
cc_45 N_A_c_34_p N_7_c_264_n 3.92093e-19 $X=0.081 $Y=0.18 $X2=0.351 $Y2=0.135
cc_46 N_A_c_3_p N_7_c_266_n 5.39672e-19 $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.135
cc_47 N_A_c_47_p N_7_c_266_n 2.96111e-19 $X=0.128 $Y=0.189 $X2=0.351 $Y2=0.135
cc_48 N_A_c_34_p N_8_c_280_n 3.30809e-19 $X=0.081 $Y=0.18 $X2=0.189 $Y2=0.135
cc_49 N_A_c_36_p N_8_c_280_n 0.00111813f $X=0.073 $Y=0.189 $X2=0.189 $Y2=0.135
cc_50 N_A_c_47_p N_8_c_280_n 6.70163e-19 $X=0.128 $Y=0.189 $X2=0.189 $Y2=0.135
cc_51 N_A_c_10_p N_8_c_283_n 2.53993e-19 $X=0.282 $Y=0.189 $X2=0.297 $Y2=0.0675
cc_52 N_A_M0_g N_8_c_284_n 2.65139e-19 $X=0.081 $Y=0.0675 $X2=0 $Y2=0
cc_53 N_A_c_36_p N_8_c_284_n 0.00233137f $X=0.073 $Y=0.189 $X2=0 $Y2=0
cc_54 N_A_c_47_p N_8_c_284_n 4.02121e-19 $X=0.128 $Y=0.189 $X2=0 $Y2=0
cc_55 N_A_c_3_p N_8_c_287_n 3.99058e-19 $X=0.135 $Y=0.135 $X2=0.351 $Y2=0.135
cc_56 N_A_c_47_p N_8_c_287_n 4.59935e-19 $X=0.128 $Y=0.189 $X2=0.351 $Y2=0.135
cc_57 N_A_M1_g N_8_c_289_n 2.61721e-19 $X=0.135 $Y=0.0675 $X2=0.351 $Y2=0.135
cc_58 N_A_c_10_p N_8_c_290_n 3.97613e-19 $X=0.282 $Y=0.189 $X2=0.351 $Y2=0.2025
cc_59 N_A_c_7_p N_8_c_291_n 3.97613e-19 $X=0.613 $Y=0.189 $X2=0.675 $Y2=0.0675
cc_60 N_A_c_12_p N_SN_c_303_n 7.36961e-19 $X=0.405 $Y=0.1645 $X2=0.297
+ $Y2=0.0675
cc_61 N_A_c_11_p N_SN_c_304_n 7.25277e-19 $X=0.405 $Y=0.135 $X2=0.351 $Y2=0.135
cc_62 N_A_c_12_p N_SN_c_305_n 7.25277e-19 $X=0.405 $Y=0.1645 $X2=0.351
+ $Y2=0.2025
cc_63 N_A_c_13_p N_SN_c_306_n 6.4841e-19 $X=0.397 $Y=0.189 $X2=0.351 $Y2=0.2025
cc_64 N_A_c_7_p N_SN_c_306_n 3.63178e-19 $X=0.613 $Y=0.189 $X2=0.351 $Y2=0.2025
cc_65 N_A_c_7_p N_SN_c_308_n 4.8223e-19 $X=0.613 $Y=0.189 $X2=0 $Y2=0
cc_66 N_A_M6_g N_SN_c_309_n 4.454e-19 $X=0.405 $Y=0.0675 $X2=0.675 $Y2=0.2025
cc_67 N_A_c_11_p N_SN_c_309_n 2.37545e-19 $X=0.405 $Y=0.135 $X2=0.675 $Y2=0.2025
cc_68 N_A_c_7_p N_SN_c_311_n 4.80144e-19 $X=0.613 $Y=0.189 $X2=0.187 $Y2=0.153
cc_69 N_A_M6_g N_SN_c_312_n 3.54161e-19 $X=0.405 $Y=0.0675 $X2=0.297 $Y2=0.153
cc_70 N_A_c_13_p N_SN_c_312_n 0.00244608f $X=0.397 $Y=0.189 $X2=0.297 $Y2=0.153
cc_71 N_A_c_7_p N_SN_c_312_n 4.0401e-19 $X=0.613 $Y=0.189 $X2=0.297 $Y2=0.153
cc_72 N_A_c_7_p N_SN_c_315_n 9.18278e-19 $X=0.613 $Y=0.189 $X2=0.297 $Y2=0.153
cc_73 N_A_c_13_p N_SN_c_316_n 3.23777e-19 $X=0.397 $Y=0.189 $X2=0.675 $Y2=0.153
cc_74 N_A_c_7_p N_SN_c_316_n 7.30118e-19 $X=0.613 $Y=0.189 $X2=0.675 $Y2=0.153
cc_75 N_A_M10_g N_10_c_349_n 3.6141e-19 $X=0.621 $Y=0.0675 $X2=0.351 $Y2=0.2025
cc_76 N_A_c_15_p N_10_c_349_n 3.82303e-19 $X=0.621 $Y=0.135 $X2=0.351 $Y2=0.2025
cc_77 N_A_c_7_p N_11_c_365_n 3.28479e-19 $X=0.613 $Y=0.189 $X2=0.189 $Y2=0.135
cc_78 N_A_c_16_p N_11_c_366_n 7.14055e-19 $X=0.621 $Y=0.167 $X2=0.297 $Y2=0.0675
cc_79 N_A_c_7_p N_11_c_367_n 0.00102531f $X=0.613 $Y=0.189 $X2=0.297 $Y2=0.135
cc_80 N_A_M10_g N_11_c_368_n 2.57834e-19 $X=0.621 $Y=0.0675 $X2=0.675 $Y2=0.0675
cc_81 N_A_c_7_p N_11_c_368_n 3.62477e-19 $X=0.613 $Y=0.189 $X2=0.675 $Y2=0.0675
cc_82 N_A_c_17_p N_11_c_368_n 0.00235846f $X=0.613 $Y=0.189 $X2=0.675 $Y2=0.0675
cc_83 N_A_c_13_p N_16_M18_s 2.50766e-19 $X=0.397 $Y=0.189 $X2=0.189 $Y2=0.0675
cc_84 N_B_M2_g N_CI_M3_g 0.00345435f $X=0.189 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_85 N_B_M4_g N_CI_M3_g 0.00341068f $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_86 N_B_M5_g N_CI_M3_g 2.13359e-19 $X=0.351 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_87 N_B_c_86_n N_CI_c_161_n 9.87435e-19 $X=0.189 $Y=0.135 $X2=0.081 $Y2=0.135
cc_88 N_B_c_89_n N_CI_c_161_n 0.00108306f $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_89 N_B_M5_g N_CI_M7_g 2.82885e-19 $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_90 N_B_M11_g N_CI_M9_g 2.13359e-19 $X=0.675 $Y=0.0675 $X2=0.405 $Y2=0.0675
cc_91 N_B_c_111_p N_CI_c_165_n 9.02142e-19 $X=0.263 $Y=0.153 $X2=0 $Y2=0
cc_92 N_B_c_101_n N_CI_c_165_n 0.00135898f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_93 N_B_c_102_n N_CI_c_165_n 0.00130683f $X=0.297 $Y=0.135 $X2=0 $Y2=0
cc_94 N_B_c_94_n N_CI_c_153_n 8.03561e-19 $X=0.587 $Y=0.153 $X2=0 $Y2=0
cc_95 N_B_c_94_n N_CI_c_154_n 8.69174e-19 $X=0.587 $Y=0.153 $X2=0.081 $Y2=0.135
cc_96 N_B_c_89_n N_CI_c_155_n 5.08852e-19 $X=0.351 $Y=0.135 $X2=0.081 $Y2=0.135
cc_97 N_B_c_111_p N_CI_c_155_n 0.0145012f $X=0.263 $Y=0.153 $X2=0.081 $Y2=0.135
cc_98 N_B_c_102_n N_CI_c_155_n 6.15506e-19 $X=0.297 $Y=0.135 $X2=0.081 $Y2=0.135
cc_99 N_B_c_94_n N_CI_c_157_n 0.0145012f $X=0.587 $Y=0.153 $X2=0 $Y2=0
cc_100 N_B_c_101_n N_CON_c_206_n 7.38096e-19 $X=0.189 $Y=0.135 $X2=0.405
+ $Y2=0.2025
cc_101 N_B_c_93_n N_CON_c_208_n 2.41745e-19 $X=0.229 $Y=0.153 $X2=0 $Y2=0
cc_102 N_B_c_101_n N_CON_c_208_n 0.00123511f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_103 N_B_M2_g N_CON_c_213_n 2.66072e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_104 N_B_c_101_n N_CON_c_213_n 0.00229458f $X=0.189 $Y=0.135 $X2=0 $Y2=0
cc_105 N_B_c_94_n N_CON_c_221_n 5.81489e-19 $X=0.587 $Y=0.153 $X2=0 $Y2=0
cc_106 N_B_c_93_n N_CON_c_222_n 0.00162526f $X=0.229 $Y=0.153 $X2=0.621
+ $Y2=0.135
cc_107 N_B_c_101_n N_CON_c_222_n 2.08291e-19 $X=0.189 $Y=0.135 $X2=0.621
+ $Y2=0.135
cc_108 N_B_c_89_n N_CON_c_224_n 2.21426e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_109 N_B_c_111_p N_CON_c_224_n 0.00162526f $X=0.263 $Y=0.153 $X2=0 $Y2=0
cc_110 N_B_c_101_n N_CON_c_226_n 3.92726e-19 $X=0.189 $Y=0.135 $X2=0.613
+ $Y2=0.189
cc_111 N_B_M2_g N_CON_c_227_n 2.61197e-19 $X=0.189 $Y=0.0675 $X2=0.613 $Y2=0.189
cc_112 N_B_c_101_n N_CON_c_227_n 8.73546e-19 $X=0.189 $Y=0.135 $X2=0.613
+ $Y2=0.189
cc_113 N_B_M2_g N_7_c_263_n 2.69932e-19 $X=0.189 $Y=0.0675 $X2=0 $Y2=0
cc_114 N_B_M2_g N_8_c_289_n 2.50481e-19 $X=0.189 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_115 N_B_M5_g N_SN_c_318_n 3.51587e-19 $X=0.351 $Y=0.0675 $X2=0.405 $Y2=0.0675
cc_116 N_B_M5_g N_SN_c_319_n 2.93361e-19 $X=0.351 $Y=0.0675 $X2=0.405 $Y2=0.0675
cc_117 N_B_M5_g N_SN_c_320_n 2.22452e-19 $X=0.351 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_118 N_B_M5_g N_SN_c_304_n 2.87785e-19 $X=0.351 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_119 N_B_c_89_n N_SN_c_304_n 0.00275831f $X=0.351 $Y=0.135 $X2=0.405 $Y2=0.135
cc_120 N_B_c_94_n N_SN_c_304_n 9.34039e-19 $X=0.587 $Y=0.153 $X2=0.405 $Y2=0.135
cc_121 N_B_c_102_n N_SN_c_304_n 0.00464886f $X=0.297 $Y=0.135 $X2=0.405
+ $Y2=0.135
cc_122 N_B_M5_g N_SN_c_325_n 2.35304e-19 $X=0.351 $Y=0.0675 $X2=0.621 $Y2=0.135
cc_123 N_B_c_143_p N_10_c_351_n 3.84788e-19 $X=0.675 $Y=0.153 $X2=0 $Y2=0
cc_124 N_B_c_143_p N_10_c_352_n 2.54113e-19 $X=0.675 $Y=0.153 $X2=0.405
+ $Y2=0.0675
cc_125 N_B_c_98_n N_10_c_353_n 2.91793e-19 $X=0.627 $Y=0.153 $X2=0.405 $Y2=0.135
cc_126 N_B_c_143_p N_11_c_366_n 3.0124e-19 $X=0.675 $Y=0.153 $X2=0.135
+ $Y2=0.0675
cc_127 N_B_c_143_p N_11_c_372_n 3.60542e-19 $X=0.675 $Y=0.153 $X2=0.405
+ $Y2=0.0675
cc_128 N_CI_M7_g N_CON_M8_g 0.00355599f $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_129 N_CI_M9_g N_CON_M8_g 0.00341068f $X=0.567 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_130 N_CI_c_150_n N_CON_c_231_n 0.00104908f $X=0.459 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_131 N_CI_c_152_n N_CON_c_231_n 0.00104908f $X=0.567 $Y=0.135 $X2=0.081
+ $Y2=0.135
cc_132 N_CI_c_165_n N_CON_c_233_n 3.29605e-19 $X=0.243 $Y=0.117 $X2=0.405
+ $Y2=0.2025
cc_133 N_CI_c_153_n N_CON_c_234_n 0.00101491f $X=0.459 $Y=0.117 $X2=0.081
+ $Y2=0.135
cc_134 N_CI_c_155_n N_CON_c_234_n 5.52177e-19 $X=0.543 $Y=0.117 $X2=0.081
+ $Y2=0.135
cc_135 N_CI_c_153_n N_CON_c_221_n 0.00120173f $X=0.459 $Y=0.117 $X2=0 $Y2=0
cc_136 N_CI_c_154_n N_CON_c_221_n 0.00184494f $X=0.573 $Y=0.117 $X2=0 $Y2=0
cc_137 N_CI_c_155_n N_CON_c_221_n 7.65244e-19 $X=0.543 $Y=0.117 $X2=0 $Y2=0
cc_138 N_CI_c_165_n N_CON_c_224_n 4.67307e-19 $X=0.243 $Y=0.117 $X2=0 $Y2=0
cc_139 N_CI_c_153_n N_CON_c_224_n 2.46239e-19 $X=0.459 $Y=0.117 $X2=0 $Y2=0
cc_140 N_CI_c_155_n N_CON_c_224_n 0.0258835f $X=0.543 $Y=0.117 $X2=0 $Y2=0
cc_141 N_CI_M3_g N_CON_c_242_n 2.14046e-19 $X=0.243 $Y=0.0675 $X2=0.397
+ $Y2=0.189
cc_142 N_CI_c_165_n N_CON_c_242_n 0.00386666f $X=0.243 $Y=0.117 $X2=0.397
+ $Y2=0.189
cc_143 N_CI_c_155_n N_CON_c_242_n 2.25232e-19 $X=0.543 $Y=0.117 $X2=0.397
+ $Y2=0.189
cc_144 N_CI_M3_g N_7_c_263_n 2.69932e-19 $X=0.243 $Y=0.0675 $X2=0 $Y2=0
cc_145 N_CI_M3_g N_8_c_293_n 3.77795e-19 $X=0.243 $Y=0.0675 $X2=0.405 $Y2=0.2025
cc_146 N_CI_c_165_n N_8_c_293_n 2.5254e-19 $X=0.243 $Y=0.117 $X2=0.405
+ $Y2=0.2025
cc_147 N_CI_c_165_n N_SN_c_320_n 3.55713e-19 $X=0.243 $Y=0.117 $X2=0.405
+ $Y2=0.135
cc_148 N_CI_c_155_n N_SN_c_320_n 8.18111e-19 $X=0.543 $Y=0.117 $X2=0.405
+ $Y2=0.135
cc_149 N_CI_c_155_n N_SN_c_304_n 3.20746e-19 $X=0.543 $Y=0.117 $X2=0.405
+ $Y2=0.135
cc_150 N_CI_M7_g N_SN_c_329_n 3.40089e-19 $X=0.459 $Y=0.0675 $X2=0.081 $Y2=0.18
cc_151 N_CI_c_153_n N_SN_c_329_n 3.40112e-19 $X=0.459 $Y=0.117 $X2=0.081
+ $Y2=0.18
cc_152 N_CI_M7_g N_SN_c_331_n 2.43117e-19 $X=0.459 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_153 N_CI_M9_g N_10_c_354_n 3.55467e-19 $X=0.567 $Y=0.0675 $X2=0.405 $Y2=0.135
cc_154 N_CI_c_200_p N_10_c_354_n 2.36327e-19 $X=0.573 $Y=0.117 $X2=0.405
+ $Y2=0.135
cc_155 N_CI_c_154_n N_10_c_354_n 7.31385e-19 $X=0.573 $Y=0.117 $X2=0.405
+ $Y2=0.135
cc_156 N_CI_M9_g N_11_c_373_n 3.67301e-19 $X=0.567 $Y=0.0675 $X2=0.405
+ $Y2=0.2025
cc_157 N_CI_c_154_n N_11_c_373_n 2.49583e-19 $X=0.573 $Y=0.117 $X2=0.405
+ $Y2=0.2025
cc_158 N_CON_c_245_p N_7_c_263_n 0.00286336f $X=0.216 $Y=0.0675 $X2=0 $Y2=0
cc_159 N_CON_c_214_n N_7_c_263_n 0.00883203f $X=0.142 $Y=0.081 $X2=0 $Y2=0
cc_160 N_CON_c_215_n N_7_c_263_n 0.00200331f $X=0.167 $Y=0.081 $X2=0 $Y2=0
cc_161 N_CON_c_248_p N_7_c_263_n 2.904e-19 $X=0.167 $Y=0.081 $X2=0 $Y2=0
cc_162 N_CON_c_245_p N_7_c_274_n 0.00358071f $X=0.216 $Y=0.0675 $X2=0.405
+ $Y2=0.0675
cc_163 N_CON_c_242_n N_7_c_274_n 0.00234221f $X=0.216 $Y=0.081 $X2=0.405
+ $Y2=0.0675
cc_164 N_CON_c_251_p N_8_c_283_n 0.00392408f $X=0.216 $Y=0.2025 $X2=0.135
+ $Y2=0.0675
cc_165 N_CON_c_211_n N_8_c_283_n 2.99306e-19 $X=0.216 $Y=0.198 $X2=0.135
+ $Y2=0.0675
cc_166 N_CON_c_251_p N_8_c_289_n 0.00278257f $X=0.216 $Y=0.2025 $X2=0.405
+ $Y2=0.135
cc_167 N_CON_c_210_n N_8_c_289_n 0.0094783f $X=0.142 $Y=0.198 $X2=0.405
+ $Y2=0.135
cc_168 N_CON_c_234_n N_SN_c_332_n 8.24577e-19 $X=0.513 $Y=0.108 $X2=0.081
+ $Y2=0.135
cc_169 N_CON_c_224_n N_SN_c_332_n 2.5959e-19 $X=0.529 $Y=0.081 $X2=0.081
+ $Y2=0.135
cc_170 N_CON_c_224_n N_SN_c_318_n 8.52063e-19 $X=0.529 $Y=0.081 $X2=0.405
+ $Y2=0.0675
cc_171 N_CON_c_242_n N_SN_c_318_n 4.38451e-19 $X=0.216 $Y=0.081 $X2=0.405
+ $Y2=0.0675
cc_172 N_CON_c_224_n N_SN_c_325_n 0.00280769f $X=0.529 $Y=0.081 $X2=0.621
+ $Y2=0.135
cc_173 N_CON_c_234_n N_10_c_357_n 0.00254473f $X=0.513 $Y=0.108 $X2=0.135
+ $Y2=0.135
cc_174 N_CON_c_234_n N_10_c_358_n 0.00126513f $X=0.513 $Y=0.108 $X2=0.405
+ $Y2=0.0675
cc_175 N_CON_c_224_n N_10_c_358_n 2.21727e-19 $X=0.529 $Y=0.081 $X2=0.405
+ $Y2=0.0675
cc_176 N_7_c_276_p N_8_c_280_n 0.00116479f $X=0.054 $Y=0.036 $X2=0.081 $Y2=0.135
cc_177 N_7_c_274_n N_8_c_283_n 0.00147414f $X=0.27 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_178 N_7_c_263_n N_SN_c_337_n 8.74938e-19 $X=0.27 $Y=0.036 $X2=0.621 $Y2=0.135
cc_179 N_7_c_263_n N_12_M2_s 2.75371e-19 $X=0.27 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_180 N_8_c_301_p N_SN_c_338_n 8.74938e-19 $X=0.27 $Y=0.234 $X2=0.081 $Y2=0.135
cc_181 N_8_c_289_n N_15_M14_s 2.23186e-19 $X=0.23 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_182 N_SN_c_332_n N_10_c_357_n 0.00401761f $X=0.486 $Y=0.0675 $X2=0.135
+ $Y2=0.135
cc_183 N_SN_c_332_n N_10_c_358_n 2.41445e-19 $X=0.486 $Y=0.0675 $X2=0.405
+ $Y2=0.0675
cc_184 N_SN_c_341_p N_10_c_358_n 0.00113918f $X=0.486 $Y=0.036 $X2=0.405
+ $Y2=0.0675
cc_185 N_SN_c_303_n N_11_c_365_n 0.00388565f $X=0.486 $Y=0.2025 $X2=0.081
+ $Y2=0.135
cc_186 N_SN_c_303_n N_11_c_367_n 2.41445e-19 $X=0.486 $Y=0.2025 $X2=0.135
+ $Y2=0.135
cc_187 N_SN_c_344_p N_11_c_367_n 0.00113918f $X=0.477 $Y=0.234 $X2=0.135
+ $Y2=0.135
cc_188 N_SN_c_325_n N_13_M6_s 2.96298e-19 $X=0.383 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_189 N_SN_c_346_p N_14_M7_s 4.56941e-19 $X=0.45 $Y=0.036 $X2=0.081 $Y2=0.0675
cc_190 N_SN_c_311_n N_16_M18_s 2.96298e-19 $X=0.383 $Y=0.234 $X2=0.081
+ $Y2=0.0675
cc_191 N_SN_c_315_n N_17_M19_s 4.56941e-19 $X=0.45 $Y=0.234 $X2=0.081 $Y2=0.0675
cc_192 N_10_c_357_n N_11_c_365_n 0.00147747f $X=0.54 $Y=0.036 $X2=0.081
+ $Y2=0.135
cc_193 N_10_c_352_n N_11_c_366_n 0.0013067f $X=0.648 $Y=0.036 $X2=0.135
+ $Y2=0.0675

* END of "./FAx1_ASAP7_75t_R.pex.sp.FAX1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: HAxp5_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 12:29:45 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "HAxp5_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./HAxp5_ASAP7_75t_R.pex.sp.pex"
* File: HAxp5_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 12:29:45 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_HAXP5_ASAP7_75T_R%A 2 5 7 10 13 15 18 20 26 31 32 33 36 41 42 43 45
+ 48 51 53 VSS
c37 53 VSS 0.00754613f $X=0.018 $Y=0.135
c38 51 VSS 4.24224e-19 $X=0.351 $Y=0.128
c39 50 VSS 0.00154135f $X=0.351 $Y=0.121
c40 48 VSS 5.24005e-20 $X=0.351 $Y=0.135
c41 45 VSS 2.41739e-19 $X=0.299 $Y=0.072
c42 44 VSS 0.00174705f $X=0.256 $Y=0.072
c43 43 VSS 1.80165e-19 $X=0.225 $Y=0.072
c44 42 VSS 0.00292169f $X=0.342 $Y=0.072
c45 41 VSS 6.38596e-24 $X=0.216 $Y=0.063
c46 36 VSS 0.00203697f $X=0.06 $Y=0.136
c47 33 VSS 0.00133719f $X=0.18 $Y=0.036
c48 32 VSS 0.00181942f $X=0.162 $Y=0.036
c49 31 VSS 0.00321912f $X=0.144 $Y=0.036
c50 30 VSS 0.00131186f $X=0.106 $Y=0.036
c51 29 VSS 0.00145201f $X=0.094 $Y=0.036
c52 28 VSS 0.00785083f $X=0.078 $Y=0.036
c53 27 VSS 0.0032309f $X=0.027 $Y=0.036
c54 26 VSS 0.00486444f $X=0.207 $Y=0.036
c55 20 VSS 8.69458e-19 $X=0.018 $Y=0.081
c56 19 VSS 6.58554e-19 $X=0.018 $Y=0.063
c57 18 VSS 0.00218042f $X=0.018 $Y=0.126
c58 13 VSS 0.00145322f $X=0.351 $Y=0.135
c59 10 VSS 0.0618866f $X=0.351 $Y=0.0675
c60 5 VSS 0.00580911f $X=0.081 $Y=0.135
c61 2 VSS 0.0638905f $X=0.081 $Y=0.0675
r62 50 51 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.121 $X2=0.351 $Y2=0.128
r63 48 51 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.128
r64 46 50 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.351
+ $Y=0.081 $X2=0.351 $Y2=0.121
r65 44 45 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.256
+ $Y=0.072 $X2=0.299 $Y2=0.072
r66 43 44 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.225
+ $Y=0.072 $X2=0.256 $Y2=0.072
r67 42 46 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.342 $Y=0.072 $X2=0.351 $Y2=0.081
r68 42 45 2.91975 $w=1.8e-08 $l=4.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.072 $X2=0.299 $Y2=0.072
r69 41 43 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.216 $Y=0.063 $X2=0.225 $Y2=0.072
r70 40 41 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.216
+ $Y=0.045 $X2=0.216 $Y2=0.063
r71 36 38 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.064 $Y=0.135 $X2=0.064
+ $Y2=0.135
r72 34 53 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.018 $Y2=0.135
r73 34 36 2.24074 $w=1.8e-08 $l=3.3e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.135 $X2=0.06 $Y2=0.135
r74 32 33 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.036 $X2=0.18 $Y2=0.036
r75 31 32 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.036 $X2=0.162 $Y2=0.036
r76 30 31 2.58025 $w=1.8e-08 $l=3.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.106
+ $Y=0.036 $X2=0.144 $Y2=0.036
r77 29 30 0.814815 $w=1.8e-08 $l=1.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.094
+ $Y=0.036 $X2=0.106 $Y2=0.036
r78 28 29 1.08642 $w=1.8e-08 $l=1.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.078
+ $Y=0.036 $X2=0.094 $Y2=0.036
r79 27 28 3.46296 $w=1.8e-08 $l=5.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.078 $Y2=0.036
r80 26 40 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.207 $Y=0.036 $X2=0.216 $Y2=0.045
r81 26 33 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.036 $X2=0.18 $Y2=0.036
r82 19 20 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.063 $X2=0.018 $Y2=0.081
r83 18 53 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.135
r84 18 20 3.05556 $w=1.8e-08 $l=4.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.126 $X2=0.018 $Y2=0.081
r85 17 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.018 $Y=0.045 $X2=0.027 $Y2=0.036
r86 17 19 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.018
+ $Y=0.045 $X2=0.018 $Y2=0.063
r87 13 48 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.351 $Y=0.135 $X2=0.351
+ $Y2=0.135
r88 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.135 $X2=0.351 $Y2=0.2025
r89 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.351
+ $Y=0.0675 $X2=0.351 $Y2=0.135
r90 5 38 15.4545 $w=2.2e-08 $l=1.7e-08 $layer=LIG $thickness=5e-08 $X=0.081
+ $Y=0.135 $X2=0.064 $Y2=0.135
r91 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.135 $X2=0.081 $Y2=0.216
r92 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.135
.ends

.subckt PM_HAXP5_ASAP7_75T_R%B 2 7 10 13 15 24 VSS
c33 24 VSS 0.00331009f $X=0.136 $Y=0.135
c34 13 VSS 0.0170781f $X=0.297 $Y=0.135
c35 10 VSS 0.0656969f $X=0.297 $Y=0.0675
c36 2 VSS 0.0637809f $X=0.135 $Y=0.0675
r37 13 15 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.135 $X2=0.297 $Y2=0.2025
r38 10 13 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.297
+ $Y=0.0675 $X2=0.297 $Y2=0.135
r39 5 13 202.5 $w=1.6e-08 $l=1.62e-07 $layer=LIG $thickness=5e-08 $X=0.135
+ $Y=0.135 $X2=0.297 $Y2=0.135
r40 5 24 6.82986 $a=2.88e-16 $layer=V0LIG $count=1 $X=0.135 $Y=0.135 $X2=0.135
+ $Y2=0.135
r41 5 7 303.467 $w=2e-08 $l=8.1e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.135 $X2=0.135 $Y2=0.216
r42 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.135
+ $Y=0.0675 $X2=0.135 $Y2=0.135
.ends

.subckt PM_HAXP5_ASAP7_75T_R%CON 2 5 7 9 12 14 15 18 19 26 27 28 30 36 38 42 43
+ 44 45 46 51 55 56 VSS
c39 56 VSS 0.00205152f $X=0.171 $Y=0.198
c40 55 VSS 6.92425e-19 $X=0.405 $Y=0.1695
c41 51 VSS 4.12414e-19 $X=0.405 $Y=0.135
c42 49 VSS 9.17737e-19 $X=0.405 $Y=0.189
c43 48 VSS 1.56568e-19 $X=0.3915 $Y=0.198
c44 47 VSS 0.00218422f $X=0.387 $Y=0.198
c45 46 VSS 8.46035e-21 $X=0.36 $Y=0.198
c46 45 VSS 9.56695e-19 $X=0.342 $Y=0.198
c47 44 VSS 0.00278191f $X=0.256 $Y=0.198
c48 43 VSS 0.00149783f $X=0.207 $Y=0.198
c49 39 VSS 7.89418e-20 $X=0.396 $Y=0.198
c50 38 VSS 9.37882e-19 $X=0.171 $Y=0.225
c51 36 VSS 7.17067e-19 $X=0.171 $Y=0.1695
c52 30 VSS 0.00149298f $X=0.171 $Y=0.09
c53 28 VSS 2.52481e-19 $X=0.171 $Y=0.189
c54 27 VSS 0.00150698f $X=0.153 $Y=0.234
c55 26 VSS 0.00287092f $X=0.144 $Y=0.234
c56 21 VSS 0.00259482f $X=0.108 $Y=0.234
c57 19 VSS 0.00458651f $X=0.162 $Y=0.234
c58 18 VSS 0.00800631f $X=0.108 $Y=0.216
c59 14 VSS 6.05457e-19 $X=0.125 $Y=0.216
c60 12 VSS 0.0148719f $X=0.16 $Y=0.0675
c61 5 VSS 0.00172642f $X=0.405 $Y=0.135
c62 2 VSS 0.0664387f $X=0.405 $Y=0.0675
r63 54 55 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.15 $X2=0.405 $Y2=0.1695
r64 51 54 1.01852 $w=1.8e-08 $l=1.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.15
r65 49 55 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.405
+ $Y=0.189 $X2=0.405 $Y2=0.1695
r66 47 48 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.387
+ $Y=0.198 $X2=0.3915 $Y2=0.198
r67 46 47 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.36
+ $Y=0.198 $X2=0.387 $Y2=0.198
r68 45 46 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.342
+ $Y=0.198 $X2=0.36 $Y2=0.198
r69 43 44 3.32716 $w=1.8e-08 $l=4.9e-08 $layer=M1 $thickness=3.6e-08 $X=0.207
+ $Y=0.198 $X2=0.256 $Y2=0.198
r70 42 45 5.77161 $w=1.8e-08 $l=8.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.257
+ $Y=0.198 $X2=0.342 $Y2=0.198
r71 42 44 0.0679012 $w=1.8e-08 $l=1e-09 $layer=M1 $thickness=3.6e-08 $X=0.257
+ $Y=0.198 $X2=0.256 $Y2=0.198
r72 40 56 0.134501 $w=3.6e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.198 $X2=0.171 $Y2=0.198
r73 40 43 1.83333 $w=1.8e-08 $l=2.7e-08 $layer=M1 $thickness=3.6e-08 $X=0.18
+ $Y=0.198 $X2=0.207 $Y2=0.198
r74 39 49 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.396 $Y=0.198 $X2=0.405 $Y2=0.189
r75 39 48 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.396
+ $Y=0.198 $X2=0.3915 $Y2=0.198
r76 37 56 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.207 $X2=0.171 $Y2=0.198
r77 37 38 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.207 $X2=0.171 $Y2=0.225
r78 35 36 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.15 $X2=0.171 $Y2=0.1695
r79 30 35 4.07407 $w=1.8e-08 $l=6e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.09 $X2=0.171 $Y2=0.15
r80 28 56 0.517544 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.189 $X2=0.171 $Y2=0.198
r81 28 36 1.32407 $w=1.8e-08 $l=1.95e-08 $layer=M1 $thickness=3.6e-08 $X=0.171
+ $Y=0.189 $X2=0.171 $Y2=0.1695
r82 26 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.144
+ $Y=0.234 $X2=0.153 $Y2=0.234
r83 21 26 2.44444 $w=1.8e-08 $l=3.6e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.144 $Y2=0.234
r84 19 38 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.162 $Y=0.234 $X2=0.171 $Y2=0.225
r85 19 27 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.162
+ $Y=0.234 $X2=0.153 $Y2=0.234
r86 18 21 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r87 15 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.216 $X2=0.108 $Y2=0.216
r88 14 18 12.5926 $w=5.4e-08 $l=1.7e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.125 $Y=0.216 $X2=0.108 $Y2=0.216
r89 12 30 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.171 $Y=0.09 $X2=0.171
+ $Y2=0.09
r90 9 12 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.145 $Y=0.0675 $X2=0.16 $Y2=0.0675
r91 5 51 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.405 $Y=0.135 $X2=0.405
+ $Y2=0.135
r92 5 7 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.135 $X2=0.405 $Y2=0.2025
r93 2 5 252.889 $w=2e-08 $l=6.75e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.405
+ $Y=0.0675 $X2=0.405 $Y2=0.135
.ends

.subckt PM_HAXP5_ASAP7_75T_R%SN 1 6 9 11 14 24 29 31 36 39 VSS
c17 39 VSS 0.00328191f $X=0.45 $Y=0.036
c18 38 VSS 0.00277971f $X=0.459 $Y=0.036
c19 36 VSS 0.00294528f $X=0.432 $Y=0.036
c20 33 VSS 2.98008e-19 $X=0.459 $Y=0.216
c21 31 VSS 0.00258114f $X=0.459 $Y=0.121
c22 30 VSS 0.00102822f $X=0.459 $Y=0.063
c23 29 VSS 0.00366991f $X=0.457 $Y=0.135
c24 27 VSS 2.81452e-19 $X=0.459 $Y=0.225
c25 25 VSS 8.76814e-19 $X=0.423 $Y=0.234
c26 24 VSS 0.0160774f $X=0.414 $Y=0.234
c27 16 VSS 0.00607607f $X=0.45 $Y=0.234
c28 14 VSS 0.00704473f $X=0.43 $Y=0.2025
c29 9 VSS 0.00505246f $X=0.272 $Y=0.2025
c30 6 VSS 4.39464e-19 $X=0.287 $Y=0.2025
c31 4 VSS 3.25039e-19 $X=0.43 $Y=0.0675
r32 39 40 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r33 38 40 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.036 $X2=0.4545 $Y2=0.036
r34 35 39 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.036 $X2=0.45 $Y2=0.036
r35 35 36 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.036 $X2=0.432
+ $Y2=0.036
r36 32 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.207 $X2=0.459 $Y2=0.216
r37 30 31 3.93827 $w=1.8e-08 $l=5.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.063 $X2=0.459 $Y2=0.121
r38 29 32 4.88889 $w=1.8e-08 $l=7.2e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.207
r39 29 31 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.135 $X2=0.459 $Y2=0.121
r40 27 33 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.225 $X2=0.459 $Y2=0.216
r41 26 38 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.036
r42 26 30 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.459
+ $Y=0.045 $X2=0.459 $Y2=0.063
r43 24 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.414
+ $Y=0.234 $X2=0.423 $Y2=0.234
r44 22 25 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.432
+ $Y=0.234 $X2=0.423 $Y2=0.234
r45 18 24 9.77778 $w=1.8e-08 $l=1.44e-07 $layer=M1 $thickness=3.6e-08 $X=0.27
+ $Y=0.234 $X2=0.414 $Y2=0.234
r46 16 27 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.45 $Y=0.234 $X2=0.459 $Y2=0.225
r47 16 22 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.45
+ $Y=0.234 $X2=0.432 $Y2=0.234
r48 14 22 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.432 $Y=0.234 $X2=0.432
+ $Y2=0.234
r49 11 14 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.415 $Y=0.2025 $X2=0.43 $Y2=0.2025
r50 9 18 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.27 $Y=0.234 $X2=0.27
+ $Y2=0.234
r51 6 9 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09 $X=0.287
+ $Y=0.2025 $X2=0.272 $Y2=0.2025
r52 4 36 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.432
+ $Y=0.0675 $X2=0.432 $Y2=0.036
r53 1 4 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09 $X=0.415
+ $Y=0.0675 $X2=0.43 $Y2=0.0675
.ends

.subckt PM_HAXP5_ASAP7_75T_R%8 1 2 VSS
c1 1 VSS 0.0022361f $X=0.125 $Y=0.0675
r2 1 2 16.7901 $w=8.1e-08 $l=3.4e-08 $layer=N_src_drn $thickness=1e-09 $X=0.125
+ $Y=0.0675 $X2=0.091 $Y2=0.0675
.ends


* END of "./HAxp5_ASAP7_75t_R.pex.sp.pex"
* 
.subckt HAxp5_ASAP7_75t_R  VSS VDD A B CON SN
* 
* SN	SN
* CON	CON
* B	B
* A	A
M0 N_8_M0_d N_A_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 N_CON_M1_d N_B_M1_g N_8_M1_s VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.125
+ $Y=0.027
M2 VSS N_B_M2_g noxref_6 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287 $Y=0.027
M3 noxref_6 N_A_M3_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.027
M4 N_SN_M4_d N_CON_M4_g noxref_6 VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.027
M5 N_CON_M5_d N_A_M5_g VDD VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.071
+ $Y=0.189
M6 VDD N_B_M6_g N_CON_M6_s VDD PMOS_RVT L=2e-08 W=5.4e-08 NFIN=2 $X=0.125
+ $Y=0.189
M7 noxref_9 N_B_M7_g N_SN_M7_s VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.287
+ $Y=0.162
M8 VDD N_A_M8_g noxref_9 VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.341 $Y=0.162
M9 N_SN_M9_d N_CON_M9_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.395
+ $Y=0.162
*
* 
* .include "HAxp5_ASAP7_75t_R.pex.sp.HAXP5_ASAP7_75T_R.pxi"
* BEGIN of "./HAxp5_ASAP7_75t_R.pex.sp.HAXP5_ASAP7_75T_R.pxi"
* File: HAxp5_ASAP7_75t_R.pex.sp.HAXP5_ASAP7_75T_R.pxi
* Created: Tue Sep  5 12:29:45 2017
* 
x_PM_HAXP5_ASAP7_75T_R%A N_A_M0_g N_A_c_5_p N_A_M5_g N_A_M3_g N_A_c_6_p N_A_M8_g
+ N_A_c_9_p N_A_c_10_p N_A_c_7_p N_A_c_2_p N_A_c_18_p N_A_c_19_p A N_A_c_20_p
+ N_A_c_32_p N_A_c_8_p N_A_c_4_p N_A_c_27_p N_A_c_28_p N_A_c_14_p VSS
+ PM_HAXP5_ASAP7_75T_R%A
x_PM_HAXP5_ASAP7_75T_R%B N_B_M1_g N_B_M6_g N_B_M2_g N_B_c_42_n N_B_M7_g B VSS
+ PM_HAXP5_ASAP7_75T_R%B
x_PM_HAXP5_ASAP7_75T_R%CON N_CON_M4_g N_CON_c_72_n N_CON_M9_g N_CON_M1_d
+ N_CON_c_73_n N_CON_M6_s N_CON_M5_d N_CON_c_88_n N_CON_c_106_p N_CON_c_89_n
+ N_CON_c_91_n N_CON_c_92_n N_CON_c_77_n N_CON_c_95_n N_CON_c_102_p CON
+ N_CON_c_96_n N_CON_c_80_n N_CON_c_81_n N_CON_c_82_n N_CON_c_84_n N_CON_c_104_p
+ N_CON_c_98_n VSS PM_HAXP5_ASAP7_75T_R%CON
x_PM_HAXP5_ASAP7_75T_R%SN N_SN_M4_d N_SN_M7_s N_SN_c_112_n N_SN_M9_d
+ N_SN_c_118_n N_SN_c_110_n SN N_SN_c_111_n N_SN_c_124_n N_SN_c_125_n VSS
+ PM_HAXP5_ASAP7_75T_R%SN
x_PM_HAXP5_ASAP7_75T_R%8 N_8_M1_s N_8_M0_d VSS PM_HAXP5_ASAP7_75T_R%8
cc_1 N_A_M0_g N_B_M1_g 0.00344695f $X=0.081 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_2 N_A_c_2_p N_B_M1_g 2.38942e-19 $X=0.144 $Y=0.036 $X2=0.135 $Y2=0.0675
cc_3 N_A_M3_g N_B_M2_g 0.00323392f $X=0.351 $Y=0.0675 $X2=0.297 $Y2=0.0675
cc_4 N_A_c_4_p N_B_M2_g 2.45429e-19 $X=0.299 $Y=0.072 $X2=0.297 $Y2=0.0675
cc_5 N_A_c_5_p N_B_c_42_n 8.12544e-19 $X=0.081 $Y=0.135 $X2=0.297 $Y2=0.135
cc_6 N_A_c_6_p N_B_c_42_n 0.00106649f $X=0.351 $Y=0.135 $X2=0.297 $Y2=0.135
cc_7 N_A_c_7_p N_B_c_42_n 3.32907e-19 $X=0.207 $Y=0.036 $X2=0.297 $Y2=0.135
cc_8 N_A_c_8_p N_B_c_42_n 0.00124812f $X=0.225 $Y=0.072 $X2=0.297 $Y2=0.135
cc_9 N_A_c_9_p B 2.57131e-19 $X=0.018 $Y=0.126 $X2=0.136 $Y2=0.135
cc_10 N_A_c_10_p B 2.3692e-19 $X=0.018 $Y=0.081 $X2=0.136 $Y2=0.135
cc_11 N_A_c_2_p B 0.00409303f $X=0.144 $Y=0.036 $X2=0.136 $Y2=0.135
cc_12 A B 4.29558e-19 $X=0.06 $Y=0.136 $X2=0.136 $Y2=0.135
cc_13 N_A_c_8_p B 3.32918e-19 $X=0.225 $Y=0.072 $X2=0.136 $Y2=0.135
cc_14 N_A_c_14_p B 8.13002e-19 $X=0.018 $Y=0.135 $X2=0.136 $Y2=0.135
cc_15 N_A_M3_g N_CON_M4_g 0.00323392f $X=0.351 $Y=0.0675 $X2=0.135 $Y2=0.0675
cc_16 N_A_c_6_p N_CON_c_72_n 9.46013e-19 $X=0.351 $Y=0.135 $X2=0.135 $Y2=0.135
cc_17 N_A_c_7_p N_CON_c_73_n 0.00142006f $X=0.207 $Y=0.036 $X2=0.297 $Y2=0.135
cc_18 N_A_c_18_p N_CON_c_73_n 0.00161143f $X=0.162 $Y=0.036 $X2=0.297 $Y2=0.135
cc_19 N_A_c_19_p N_CON_c_73_n 0.00130888f $X=0.18 $Y=0.036 $X2=0.297 $Y2=0.135
cc_20 N_A_c_20_p N_CON_c_73_n 7.82924e-19 $X=0.216 $Y=0.063 $X2=0.297 $Y2=0.135
cc_21 N_A_c_19_p N_CON_c_77_n 8.69266e-19 $X=0.18 $Y=0.036 $X2=0 $Y2=0
cc_22 N_A_c_8_p N_CON_c_77_n 3.12063e-19 $X=0.225 $Y=0.072 $X2=0 $Y2=0
cc_23 N_A_c_14_p N_CON_c_77_n 2.69986e-19 $X=0.018 $Y=0.135 $X2=0 $Y2=0
cc_24 N_A_c_8_p N_CON_c_80_n 7.71444e-19 $X=0.225 $Y=0.072 $X2=0 $Y2=0
cc_25 N_A_c_4_p N_CON_c_81_n 7.71444e-19 $X=0.299 $Y=0.072 $X2=0 $Y2=0
cc_26 N_A_M3_g N_CON_c_82_n 3.0688e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_27 N_A_c_27_p N_CON_c_82_n 8.07817e-19 $X=0.351 $Y=0.135 $X2=0 $Y2=0
cc_28 N_A_c_28_p N_CON_c_84_n 0.00118958f $X=0.351 $Y=0.128 $X2=0 $Y2=0
cc_29 VSS N_A_c_4_p 3.29233e-19 $X=0.299 $Y=0.072 $X2=0.135 $Y2=0.0675
cc_30 VSS N_A_c_20_p 6.7861e-19 $X=0.216 $Y=0.063 $X2=0.297 $Y2=0.135
cc_31 VSS N_A_c_4_p 0.00219077f $X=0.299 $Y=0.072 $X2=0.297 $Y2=0.135
cc_32 VSS N_A_c_32_p 0.00158538f $X=0.342 $Y=0.072 $X2=0 $Y2=0
cc_33 VSS N_A_M3_g 2.34993e-19 $X=0.351 $Y=0.0675 $X2=0 $Y2=0
cc_34 VSS N_A_c_7_p 0.00123555f $X=0.207 $Y=0.036 $X2=0 $Y2=0
cc_35 VSS N_A_c_4_p 0.00880208f $X=0.299 $Y=0.072 $X2=0 $Y2=0
cc_36 N_A_M3_g N_SN_c_110_n 2.38303e-19 $X=0.351 $Y=0.0675 $X2=0.136 $Y2=0.135
cc_37 N_A_c_32_p N_SN_c_111_n 6.03287e-19 $X=0.342 $Y=0.072 $X2=0 $Y2=0
cc_38 N_B_M2_g N_CON_M4_g 2.34385e-19 $X=0.297 $Y=0.0675 $X2=0.081 $Y2=0.0675
cc_39 N_B_c_42_n N_CON_c_73_n 0.00369057f $X=0.297 $Y=0.135 $X2=0.351 $Y2=0.135
cc_40 B N_CON_c_73_n 5.10449e-19 $X=0.136 $Y=0.135 $X2=0.351 $Y2=0.135
cc_41 B N_CON_c_88_n 0.00184579f $X=0.136 $Y=0.135 $X2=0.018 $Y2=0.126
cc_42 N_B_M1_g N_CON_c_89_n 2.35623e-19 $X=0.135 $Y=0.0675 $X2=0.207 $Y2=0.036
cc_43 B N_CON_c_89_n 0.00374777f $X=0.136 $Y=0.135 $X2=0.207 $Y2=0.036
cc_44 N_B_c_42_n N_CON_c_91_n 2.91977e-19 $X=0.297 $Y=0.135 $X2=0.027 $Y2=0.036
cc_45 B N_CON_c_92_n 0.00183916f $X=0.136 $Y=0.135 $X2=0.078 $Y2=0.036
cc_46 N_B_c_42_n N_CON_c_77_n 0.00250832f $X=0.297 $Y=0.135 $X2=0.106 $Y2=0.036
cc_47 B N_CON_c_77_n 0.00551748f $X=0.136 $Y=0.135 $X2=0.106 $Y2=0.036
cc_48 B N_CON_c_95_n 0.00183916f $X=0.136 $Y=0.135 $X2=0.06 $Y2=0.136
cc_49 N_B_c_42_n N_CON_c_96_n 0.00135939f $X=0.297 $Y=0.135 $X2=0.225 $Y2=0.072
cc_50 N_B_M2_g N_CON_c_81_n 4.09048e-19 $X=0.297 $Y=0.0675 $X2=0.299 $Y2=0.072
cc_51 B N_CON_c_98_n 0.00183916f $X=0.136 $Y=0.135 $X2=0.081 $Y2=0.135
cc_52 VSS N_B_c_42_n 6.8292e-19 $X=0.297 $Y=0.135 $X2=0.351 $Y2=0.135
cc_53 VSS N_B_M2_g 2.65491e-19 $X=0.297 $Y=0.0675 $X2=0.018 $Y2=0.126
cc_54 N_B_c_42_n N_SN_c_112_n 6.8292e-19 $X=0.297 $Y=0.135 $X2=0.351 $Y2=0.0675
cc_55 N_B_M2_g N_SN_c_110_n 2.65491e-19 $X=0.297 $Y=0.0675 $X2=0 $Y2=0
cc_56 B N_8_M1_s 2.02285e-19 $X=0.136 $Y=0.135 $X2=0.081 $Y2=0.0675
cc_57 VSS N_CON_c_73_n 0.00221794f $X=0.16 $Y=0.0675 $X2=0.351 $Y2=0.135
cc_58 N_CON_c_81_n N_SN_M7_s 3.29233e-19 $X=0.342 $Y=0.198 $X2=0.081 $Y2=0.216
cc_59 N_CON_c_95_n N_SN_c_112_n 5.55768e-19 $X=0.171 $Y=0.1695 $X2=0.351
+ $Y2=0.0675
cc_60 N_CON_c_102_p N_SN_c_112_n 2.38811e-19 $X=0.171 $Y=0.225 $X2=0.351
+ $Y2=0.0675
cc_61 N_CON_c_81_n N_SN_c_112_n 0.00284111f $X=0.342 $Y=0.198 $X2=0.351
+ $Y2=0.0675
cc_62 N_CON_c_104_p N_SN_c_118_n 0.00135952f $X=0.405 $Y=0.1695 $X2=0.351
+ $Y2=0.2025
cc_63 N_CON_M4_g N_SN_c_110_n 2.34993e-19 $X=0.405 $Y=0.0675 $X2=0 $Y2=0
cc_64 N_CON_c_106_p N_SN_c_110_n 5.49907e-19 $X=0.162 $Y=0.234 $X2=0 $Y2=0
cc_65 N_CON_c_81_n N_SN_c_110_n 0.0133208f $X=0.342 $Y=0.198 $X2=0 $Y2=0
cc_66 N_CON_c_84_n SN 0.0034418f $X=0.405 $Y=0.135 $X2=0.094 $Y2=0.036
cc_67 VSS N_CON_c_81_n 5.15356e-19 $X=0.342 $Y=0.198 $X2=0.081 $Y2=0.0675
cc_68 VSS N_SN_c_112_n 0.00169333f $X=0.27 $Y=0.036 $X2=0.351 $Y2=0.0675
cc_69 VSS N_SN_c_124_n 0.00395939f $X=0.378 $Y=0.036 $X2=0.06 $Y2=0.136
cc_70 VSS N_SN_c_125_n 6.5272e-19 $X=0.378 $Y=0.036 $X2=0 $Y2=0
cc_71 VSS N_SN_c_110_n 3.33359e-19 $X=0.414 $Y=0.234 $X2=0.081 $Y2=0.0675

* END of "./HAxp5_ASAP7_75t_R.pex.sp.HAXP5_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: TIEHIx1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:06:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "TIEHIx1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./TIEHIx1_ASAP7_75t_R.pex.sp.pex"
* File: TIEHIx1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:06:03 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_TIEHIX1_ASAP7_75T_R%H 2 5 7 10 14 19 24 25 26 VSS
c12 34 VSS 0.00256321f $X=0.126 $Y=0.234
c13 33 VSS 0.00278032f $X=0.135 $Y=0.234
c14 28 VSS 0.00175467f $X=0.108 $Y=0.234
c15 26 VSS 0.00114837f $X=0.135 $Y=0.146
c16 25 VSS 0.00182701f $X=0.135 $Y=0.128
c17 22 VSS 0.00397056f $X=0.135 $Y=0.225
c18 20 VSS 2.74234e-19 $X=0.1105 $Y=0.079
c19 19 VSS 5.05338e-19 $X=0.095 $Y=0.079
c20 14 VSS 3.32709e-19 $X=0.081 $Y=0.079
c21 12 VSS 0.00267656f $X=0.126 $Y=0.079
c22 10 VSS 0.00782082f $X=0.106 $Y=0.2025
c23 5 VSS 0.00449381f $X=0.081 $Y=0.079
r24 34 35 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r25 33 35 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.234 $X2=0.1305 $Y2=0.234
r26 28 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.234 $X2=0.126 $Y2=0.234
r27 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.128 $X2=0.135 $Y2=0.146
r28 24 26 3.22531 $w=1.8e-08 $l=4.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.1935 $X2=0.135 $Y2=0.146
r29 22 33 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.234
r30 22 24 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.225 $X2=0.135 $Y2=0.1935
r31 21 25 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.088 $X2=0.135 $Y2=0.128
r32 19 20 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.079 $X2=0.1105 $Y2=0.079
r33 14 19 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.079 $X2=0.095 $Y2=0.079
r34 12 21 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.126 $Y=0.079 $X2=0.135 $Y2=0.088
r35 12 20 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.079 $X2=0.1105 $Y2=0.079
r36 10 28 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.234 $X2=0.108
+ $Y2=0.234
r37 7 10 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.2025 $X2=0.106 $Y2=0.2025
r38 5 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.079 $X2=0.081
+ $Y2=0.079
r39 2 5 137.749 $w=2e-08 $l=3.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0405 $X2=0.081 $Y2=0.079
.ends

.subckt PM_TIEHIX1_ASAP7_75T_R%4 2 5 7 10 13 14 15 18 21 VSS
c12 30 VSS 7.11107e-19 $X=0.045 $Y=0.036
c13 29 VSS 0.00327678f $X=0.036 $Y=0.036
c14 27 VSS 0.00319097f $X=0.054 $Y=0.036
c15 21 VSS 8.592e-20 $X=0.074 $Y=0.137
c16 20 VSS 8.34396e-19 $X=0.067 $Y=0.137
c17 18 VSS 3.52763e-19 $X=0.081 $Y=0.137
c18 16 VSS 0.0019543f $X=0.036 $Y=0.137
c19 15 VSS 7.43234e-19 $X=0.027 $Y=0.088
c20 14 VSS 0.00125918f $X=0.027 $Y=0.07
c21 13 VSS 0.00182701f $X=0.027 $Y=0.128
c22 10 VSS 0.00470034f $X=0.056 $Y=0.0405
c23 7 VSS 4.65731e-19 $X=0.071 $Y=0.0405
c24 2 VSS 0.0898363f $X=0.081 $Y=0.137
r25 29 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.036 $X2=0.045 $Y2=0.036
r26 27 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.036 $X2=0.045 $Y2=0.036
r27 24 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.036 $X2=0.036 $Y2=0.036
r28 20 21 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.067
+ $Y=0.137 $X2=0.074 $Y2=0.137
r29 18 21 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.137 $X2=0.074 $Y2=0.137
r30 16 20 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.137 $X2=0.067 $Y2=0.137
r31 14 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.07 $X2=0.027 $Y2=0.088
r32 13 16 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.128 $X2=0.036 $Y2=0.137
r33 13 15 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.128 $X2=0.027 $Y2=0.088
r34 12 24 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.036
r35 12 14 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.045 $X2=0.027 $Y2=0.07
r36 10 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.036 $X2=0.054
+ $Y2=0.036
r37 7 10 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.0405 $X2=0.056 $Y2=0.0405
r38 2 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.137 $X2=0.081
+ $Y2=0.137
r39 2 5 240.554 $w=2e-08 $l=6.55e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.137 $X2=0.081 $Y2=0.2025
.ends


* END of "./TIEHIx1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt TIEHIx1_ASAP7_75t_R  VSS VDD H
* 
* H	H
M0 VSS N_H_M0_g N_4_M0_s VSS NMOS_RVT L=2e-08 W=2.7e-08 NFIN=1 $X=0.071 $Y=0.027
M1 N_H_M1_d N_4_M1_g VDD VDD PMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.162
*
* 
* .include "TIEHIx1_ASAP7_75t_R.pex.sp.TIEHIX1_ASAP7_75T_R.pxi"
* BEGIN of "./TIEHIx1_ASAP7_75t_R.pex.sp.TIEHIX1_ASAP7_75T_R.pxi"
* File: TIEHIx1_ASAP7_75t_R.pex.sp.TIEHIX1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:06:03 2017
* 
x_PM_TIEHIX1_ASAP7_75T_R%H N_H_M0_g N_H_c_1_p N_H_M1_d N_H_c_2_p N_H_c_3_p
+ N_H_c_10_p H N_H_c_4_p N_H_c_11_p VSS PM_TIEHIX1_ASAP7_75T_R%H
x_PM_TIEHIX1_ASAP7_75T_R%4 N_4_c_13_n N_4_M1_g N_4_M0_s N_4_c_17_n N_4_c_18_n
+ N_4_c_19_n N_4_c_20_n N_4_c_21_n N_4_c_24_n VSS PM_TIEHIX1_ASAP7_75T_R%4
cc_1 N_H_c_1_p N_4_c_13_n 0.00553621f $X=0.081 $Y=0.079 $X2=0.081 $Y2=0.137
cc_2 N_H_c_2_p N_4_c_13_n 5.73423e-19 $X=0.106 $Y=0.2025 $X2=0.081 $Y2=0.137
cc_3 N_H_c_3_p N_4_c_13_n 2.12306e-19 $X=0.081 $Y=0.079 $X2=0.081 $Y2=0.137
cc_4 N_H_c_4_p N_4_c_13_n 5.60768e-19 $X=0.135 $Y=0.128 $X2=0.081 $Y2=0.137
cc_5 N_H_c_1_p N_4_c_17_n 4.40669e-19 $X=0.081 $Y=0.079 $X2=0.056 $Y2=0.0405
cc_6 N_H_c_4_p N_4_c_18_n 7.07225e-19 $X=0.135 $Y=0.128 $X2=0.027 $Y2=0.128
cc_7 N_H_c_1_p N_4_c_19_n 5.65652e-19 $X=0.081 $Y=0.079 $X2=0.027 $Y2=0.07
cc_8 N_H_c_3_p N_4_c_20_n 8.26176e-19 $X=0.081 $Y=0.079 $X2=0.027 $Y2=0.088
cc_9 N_H_c_3_p N_4_c_21_n 2.65646e-19 $X=0.081 $Y=0.079 $X2=0.081 $Y2=0.137
cc_10 N_H_c_10_p N_4_c_21_n 2.65646e-19 $X=0.095 $Y=0.079 $X2=0.081 $Y2=0.137
cc_11 N_H_c_11_p N_4_c_21_n 8.2057e-19 $X=0.135 $Y=0.146 $X2=0.081 $Y2=0.137
cc_12 N_H_c_3_p N_4_c_24_n 2.65646e-19 $X=0.081 $Y=0.079 $X2=0.074 $Y2=0.137

* END of "./TIEHIx1_ASAP7_75t_R.pex.sp.TIEHIX1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

* File: TIELOx1_ASAP7_75t_R.pex.sp
* Created: Tue Sep  5 13:06:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* 
* 
* .include "TIELOx1_ASAP7_75t_R.pex.sp.pex"
* BEGIN of "./TIELOx1_ASAP7_75t_R.pex.sp.pex"
* File: TIELOx1_ASAP7_75t_R.pex.sp.pex
* Created: Tue Sep  5 13:06:25 2017
* Program "Calibre xRC"
* Version "v2017.1_34.33"
* Nominal Temperature: 25C
* Circuit Temperature: 27C
* 
.subckt PM_TIELOX1_ASAP7_75T_R%3 2 5 7 10 14 15 18 21 VSS
c12 30 VSS 7.11107e-19 $X=0.045 $Y=0.234
c13 29 VSS 0.00327678f $X=0.036 $Y=0.234
c14 27 VSS 0.00319097f $X=0.054 $Y=0.234
c15 21 VSS 8.592e-20 $X=0.074 $Y=0.133
c16 20 VSS 8.34396e-19 $X=0.067 $Y=0.133
c17 18 VSS 3.52763e-19 $X=0.081 $Y=0.133
c18 16 VSS 0.00196342f $X=0.036 $Y=0.133
c19 15 VSS 7.43234e-19 $X=0.027 $Y=0.2
c20 14 VSS 0.00182701f $X=0.027 $Y=0.182
c21 13 VSS 0.00125918f $X=0.027 $Y=0.225
c22 10 VSS 0.00470034f $X=0.056 $Y=0.2295
c23 7 VSS 4.65731e-19 $X=0.071 $Y=0.2295
c24 5 VSS 0.00393353f $X=0.081 $Y=0.133
c25 2 VSS 0.0354269f $X=0.081 $Y=0.0675
r26 29 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.234 $X2=0.045 $Y2=0.234
r27 27 30 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.054
+ $Y=0.234 $X2=0.045 $Y2=0.234
r28 24 29 0.611111 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.234 $X2=0.036 $Y2=0.234
r29 20 21 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.067
+ $Y=0.133 $X2=0.074 $Y2=0.133
r30 18 21 0.475309 $w=1.8e-08 $l=7e-09 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.133 $X2=0.074 $Y2=0.133
r31 16 20 2.10494 $w=1.8e-08 $l=3.1e-08 $layer=M1 $thickness=3.6e-08 $X=0.036
+ $Y=0.133 $X2=0.067 $Y2=0.133
r32 14 15 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.182 $X2=0.027 $Y2=0.2
r33 13 24 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.234
r34 13 15 1.69753 $w=1.8e-08 $l=2.5e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.225 $X2=0.027 $Y2=0.2
r35 12 16 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.027 $Y=0.142 $X2=0.036 $Y2=0.133
r36 12 14 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.027
+ $Y=0.142 $X2=0.027 $Y2=0.182
r37 10 27 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.054 $Y=0.234 $X2=0.054
+ $Y2=0.234
r38 7 10 22.2222 $w=2.7e-08 $l=1.5e-08 $layer=P_src_drn $thickness=1e-09
+ $X=0.071 $Y=0.2295 $X2=0.056 $Y2=0.2295
r39 5 18 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.133 $X2=0.081
+ $Y2=0.133
r40 2 5 240.554 $w=2e-08 $l=6.55e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.0675 $X2=0.081 $Y2=0.133
.ends

.subckt PM_TIELOX1_ASAP7_75T_R%L 2 5 7 14 19 22 24 26 29 VSS
c12 34 VSS 0.00256321f $X=0.126 $Y=0.036
c13 33 VSS 0.00278032f $X=0.135 $Y=0.036
c14 29 VSS 0.00733468f $X=0.108 $Y=0.036
c15 28 VSS 0.00175467f $X=0.108 $Y=0.036
c16 26 VSS 0.00114837f $X=0.135 $Y=0.142
c17 24 VSS 0.00397056f $X=0.137 $Y=0.0765
c18 22 VSS 0.00182701f $X=0.135 $Y=0.182
c19 20 VSS 2.74234e-19 $X=0.1105 $Y=0.191
c20 19 VSS 5.05338e-19 $X=0.095 $Y=0.191
c21 14 VSS 3.32709e-19 $X=0.081 $Y=0.191
c22 12 VSS 0.00267656f $X=0.126 $Y=0.191
c23 10 VSS 4.86139e-19 $X=0.106 $Y=0.0675
c24 2 VSS 0.0549696f $X=0.081 $Y=0.191
r25 34 35 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r26 33 35 0.305556 $w=1.8e-08 $l=4.5e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.036 $X2=0.1305 $Y2=0.036
r27 28 34 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.108
+ $Y=0.036 $X2=0.126 $Y2=0.036
r28 28 29 6.07099 $a=3.24e-16 $layer=V0LISD $count=1 $X=0.108 $Y=0.036 $X2=0.108
+ $Y2=0.036
r29 25 26 1.22222 $w=1.8e-08 $l=1.8e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.124 $X2=0.135 $Y2=0.142
r30 24 25 3.22531 $w=1.8e-08 $l=4.75e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.0765 $X2=0.135 $Y2=0.124
r31 22 26 2.71605 $w=1.8e-08 $l=4e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.182 $X2=0.135 $Y2=0.142
r32 21 33 0.0717796 $w=1.8e-08 $l=9e-09 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.036
r33 21 24 2.13889 $w=1.8e-08 $l=3.15e-08 $layer=M1 $thickness=3.6e-08 $X=0.135
+ $Y=0.045 $X2=0.135 $Y2=0.0765
r34 19 20 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.095
+ $Y=0.191 $X2=0.1105 $Y2=0.191
r35 14 19 0.950617 $w=1.8e-08 $l=1.4e-08 $layer=M1 $thickness=3.6e-08 $X=0.081
+ $Y=0.191 $X2=0.095 $Y2=0.191
r36 12 22 0.682891 $w=1.8e-08 $l=1.27279e-08 $layer=M1 $thickness=3.6e-08
+ $X=0.126 $Y=0.191 $X2=0.135 $Y2=0.182
r37 12 20 1.05247 $w=1.8e-08 $l=1.55e-08 $layer=M1 $thickness=3.6e-08 $X=0.126
+ $Y=0.191 $X2=0.1105 $Y2=0.191
r38 10 29 27.1875 $w=2.4e-08 $l=3.15e-08 $layer=LISD $thickness=2.8e-08 $X=0.108
+ $Y=0.0675 $X2=0.108 $Y2=0.036
r39 7 10 7.40741 $w=8.1e-08 $l=1.5e-08 $layer=N_src_drn $thickness=1e-09
+ $X=0.091 $Y=0.0675 $X2=0.106 $Y2=0.0675
r40 2 14 6.07099 $a=3.24e-16 $layer=V0LIG $count=1 $X=0.081 $Y=0.191 $X2=0.081
+ $Y2=0.191
r41 2 5 137.749 $w=2e-08 $l=3.85e-08 $layer=Gate_1 $thickness=5.6e-08 $X=0.081
+ $Y=0.191 $X2=0.081 $Y2=0.2295
.ends


* END of "./TIELOx1_ASAP7_75t_R.pex.sp.pex"
* 
.subckt TIELOx1_ASAP7_75t_R  VSS VDD L
* 
* L	L
M0 N_L_M0_d N_3_M0_g VSS VSS NMOS_RVT L=2e-08 W=8.1e-08 NFIN=3 $X=0.071 $Y=0.027
M1 VDD N_L_M1_g N_3_M1_s VDD PMOS_RVT L=2e-08 W=2.7e-08 NFIN=1 $X=0.071 $Y=0.216
*
* 
* .include "TIELOx1_ASAP7_75t_R.pex.sp.TIELOX1_ASAP7_75T_R.pxi"
* BEGIN of "./TIELOx1_ASAP7_75t_R.pex.sp.TIELOX1_ASAP7_75T_R.pxi"
* File: TIELOx1_ASAP7_75t_R.pex.sp.TIELOX1_ASAP7_75T_R.pxi
* Created: Tue Sep  5 13:06:25 2017
* 
x_PM_TIELOX1_ASAP7_75T_R%3 N_3_M0_g N_3_c_1_p N_3_M1_s N_3_c_2_p N_3_c_3_p
+ N_3_c_5_p N_3_c_6_p N_3_c_7_p VSS PM_TIELOX1_ASAP7_75T_R%3
x_PM_TIELOX1_ASAP7_75T_R%L N_L_c_13_n N_L_M1_g N_L_M0_d N_L_c_16_n N_L_c_20_n
+ N_L_c_21_n L N_L_c_23_n N_L_c_24_n VSS PM_TIELOX1_ASAP7_75T_R%L
cc_1 N_3_c_1_p N_L_c_13_n 0.00414874f $X=0.081 $Y=0.133 $X2=0.081 $Y2=0.191
cc_2 N_3_c_2_p N_L_c_13_n 4.40669e-19 $X=0.056 $Y=0.2295 $X2=0.081 $Y2=0.191
cc_3 N_3_c_3_p N_L_c_13_n 5.65652e-19 $X=0.027 $Y=0.182 $X2=0.081 $Y2=0.191
cc_4 N_3_c_1_p N_L_c_16_n 2.12306e-19 $X=0.081 $Y=0.133 $X2=0.081 $Y2=0.191
cc_5 N_3_c_5_p N_L_c_16_n 8.26176e-19 $X=0.027 $Y=0.2 $X2=0.081 $Y2=0.191
cc_6 N_3_c_6_p N_L_c_16_n 2.65646e-19 $X=0.081 $Y=0.133 $X2=0.081 $Y2=0.191
cc_7 N_3_c_7_p N_L_c_16_n 2.65646e-19 $X=0.074 $Y=0.133 $X2=0.081 $Y2=0.191
cc_8 N_3_c_6_p N_L_c_20_n 2.65646e-19 $X=0.081 $Y=0.133 $X2=0.095 $Y2=0.191
cc_9 N_3_c_3_p N_L_c_21_n 7.07225e-19 $X=0.027 $Y=0.182 $X2=0.135 $Y2=0.182
cc_10 N_3_c_1_p L 5.60768e-19 $X=0.081 $Y=0.133 $X2=0.137 $Y2=0.0765
cc_11 N_3_c_6_p N_L_c_23_n 8.2057e-19 $X=0.081 $Y=0.133 $X2=0.135 $Y2=0.142
cc_12 N_3_c_1_p N_L_c_24_n 5.73423e-19 $X=0.081 $Y=0.133 $X2=0.108 $Y2=0.036

* END of "./TIELOx1_ASAP7_75t_R.pex.sp.TIELOX1_ASAP7_75T_R.pxi"
* 
*
.ends
*
*

